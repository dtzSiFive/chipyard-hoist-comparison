// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module LSU_1(
  input         clock,
                reset,
                io_ptw_req_ready,
                io_ptw_resp_valid,
                io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
                io_ptw_resp_bits_pte_a,
                io_ptw_resp_bits_pte_g,
                io_ptw_resp_bits_pte_u,
                io_ptw_resp_bits_pte_x,
                io_ptw_resp_bits_pte_w,
                io_ptw_resp_bits_pte_r,
                io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
                io_ptw_status_sum,
                io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
                io_ptw_pmp_0_cfg_w,
                io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
                io_ptw_pmp_1_cfg_w,
                io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
                io_ptw_pmp_2_cfg_w,
                io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
                io_ptw_pmp_3_cfg_w,
                io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
                io_ptw_pmp_4_cfg_w,
                io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
                io_ptw_pmp_5_cfg_w,
                io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
                io_ptw_pmp_6_cfg_w,
                io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
                io_ptw_pmp_7_cfg_w,
                io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_core_exe_0_req_valid,
  input  [6:0]  io_core_exe_0_req_bits_uop_uopc,
  input  [31:0] io_core_exe_0_req_bits_uop_inst,
                io_core_exe_0_req_bits_uop_debug_inst,
  input         io_core_exe_0_req_bits_uop_is_rvc,
  input  [39:0] io_core_exe_0_req_bits_uop_debug_pc,
  input  [2:0]  io_core_exe_0_req_bits_uop_iq_type,
  input  [9:0]  io_core_exe_0_req_bits_uop_fu_code,
  input  [3:0]  io_core_exe_0_req_bits_uop_ctrl_br_type,
  input  [1:0]  io_core_exe_0_req_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_core_exe_0_req_bits_uop_ctrl_op2_sel,
                io_core_exe_0_req_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_core_exe_0_req_bits_uop_ctrl_op_fcn,
  input         io_core_exe_0_req_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_core_exe_0_req_bits_uop_ctrl_csr_cmd,
  input         io_core_exe_0_req_bits_uop_ctrl_is_load,
                io_core_exe_0_req_bits_uop_ctrl_is_sta,
                io_core_exe_0_req_bits_uop_ctrl_is_std,
  input  [1:0]  io_core_exe_0_req_bits_uop_iw_state,
  input         io_core_exe_0_req_bits_uop_iw_p1_poisoned,
                io_core_exe_0_req_bits_uop_iw_p2_poisoned,
                io_core_exe_0_req_bits_uop_is_br,
                io_core_exe_0_req_bits_uop_is_jalr,
                io_core_exe_0_req_bits_uop_is_jal,
                io_core_exe_0_req_bits_uop_is_sfb,
  input  [15:0] io_core_exe_0_req_bits_uop_br_mask,
  input  [3:0]  io_core_exe_0_req_bits_uop_br_tag,
  input  [4:0]  io_core_exe_0_req_bits_uop_ftq_idx,
  input         io_core_exe_0_req_bits_uop_edge_inst,
  input  [5:0]  io_core_exe_0_req_bits_uop_pc_lob,
  input         io_core_exe_0_req_bits_uop_taken,
  input  [19:0] io_core_exe_0_req_bits_uop_imm_packed,
  input  [11:0] io_core_exe_0_req_bits_uop_csr_addr,
  input  [6:0]  io_core_exe_0_req_bits_uop_rob_idx,
  input  [4:0]  io_core_exe_0_req_bits_uop_ldq_idx,
                io_core_exe_0_req_bits_uop_stq_idx,
  input  [1:0]  io_core_exe_0_req_bits_uop_rxq_idx,
  input  [6:0]  io_core_exe_0_req_bits_uop_pdst,
                io_core_exe_0_req_bits_uop_prs1,
                io_core_exe_0_req_bits_uop_prs2,
                io_core_exe_0_req_bits_uop_prs3,
  input  [4:0]  io_core_exe_0_req_bits_uop_ppred,
  input         io_core_exe_0_req_bits_uop_prs1_busy,
                io_core_exe_0_req_bits_uop_prs2_busy,
                io_core_exe_0_req_bits_uop_prs3_busy,
                io_core_exe_0_req_bits_uop_ppred_busy,
  input  [6:0]  io_core_exe_0_req_bits_uop_stale_pdst,
  input         io_core_exe_0_req_bits_uop_exception,
  input  [63:0] io_core_exe_0_req_bits_uop_exc_cause,
  input         io_core_exe_0_req_bits_uop_bypassable,
  input  [4:0]  io_core_exe_0_req_bits_uop_mem_cmd,
  input  [1:0]  io_core_exe_0_req_bits_uop_mem_size,
  input         io_core_exe_0_req_bits_uop_mem_signed,
                io_core_exe_0_req_bits_uop_is_fence,
                io_core_exe_0_req_bits_uop_is_fencei,
                io_core_exe_0_req_bits_uop_is_amo,
                io_core_exe_0_req_bits_uop_uses_ldq,
                io_core_exe_0_req_bits_uop_uses_stq,
                io_core_exe_0_req_bits_uop_is_sys_pc2epc,
                io_core_exe_0_req_bits_uop_is_unique,
                io_core_exe_0_req_bits_uop_flush_on_commit,
                io_core_exe_0_req_bits_uop_ldst_is_rs1,
  input  [5:0]  io_core_exe_0_req_bits_uop_ldst,
                io_core_exe_0_req_bits_uop_lrs1,
                io_core_exe_0_req_bits_uop_lrs2,
                io_core_exe_0_req_bits_uop_lrs3,
  input         io_core_exe_0_req_bits_uop_ldst_val,
  input  [1:0]  io_core_exe_0_req_bits_uop_dst_rtype,
                io_core_exe_0_req_bits_uop_lrs1_rtype,
                io_core_exe_0_req_bits_uop_lrs2_rtype,
  input         io_core_exe_0_req_bits_uop_frs3_en,
                io_core_exe_0_req_bits_uop_fp_val,
                io_core_exe_0_req_bits_uop_fp_single,
                io_core_exe_0_req_bits_uop_xcpt_pf_if,
                io_core_exe_0_req_bits_uop_xcpt_ae_if,
                io_core_exe_0_req_bits_uop_xcpt_ma_if,
                io_core_exe_0_req_bits_uop_bp_debug_if,
                io_core_exe_0_req_bits_uop_bp_xcpt_if,
  input  [1:0]  io_core_exe_0_req_bits_uop_debug_fsrc,
                io_core_exe_0_req_bits_uop_debug_tsrc,
  input  [63:0] io_core_exe_0_req_bits_data,
  input  [39:0] io_core_exe_0_req_bits_addr,
  input         io_core_exe_0_req_bits_mxcpt_valid,
                io_core_exe_0_req_bits_sfence_valid,
                io_core_exe_0_req_bits_sfence_bits_rs1,
                io_core_exe_0_req_bits_sfence_bits_rs2,
  input  [38:0] io_core_exe_0_req_bits_sfence_bits_addr,
  input         io_core_dis_uops_0_valid,
  input  [6:0]  io_core_dis_uops_0_bits_uopc,
  input  [31:0] io_core_dis_uops_0_bits_inst,
                io_core_dis_uops_0_bits_debug_inst,
  input         io_core_dis_uops_0_bits_is_rvc,
  input  [39:0] io_core_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_0_bits_iq_type,
  input  [9:0]  io_core_dis_uops_0_bits_fu_code,
  input  [3:0]  io_core_dis_uops_0_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_0_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_0_bits_ctrl_op2_sel,
                io_core_dis_uops_0_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_0_bits_ctrl_op_fcn,
  input         io_core_dis_uops_0_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_0_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_0_bits_ctrl_is_load,
                io_core_dis_uops_0_bits_ctrl_is_sta,
                io_core_dis_uops_0_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_0_bits_iw_state,
  input         io_core_dis_uops_0_bits_iw_p1_poisoned,
                io_core_dis_uops_0_bits_iw_p2_poisoned,
                io_core_dis_uops_0_bits_is_br,
                io_core_dis_uops_0_bits_is_jalr,
                io_core_dis_uops_0_bits_is_jal,
                io_core_dis_uops_0_bits_is_sfb,
  input  [15:0] io_core_dis_uops_0_bits_br_mask,
  input  [3:0]  io_core_dis_uops_0_bits_br_tag,
  input  [4:0]  io_core_dis_uops_0_bits_ftq_idx,
  input         io_core_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_0_bits_pc_lob,
  input         io_core_dis_uops_0_bits_taken,
  input  [19:0] io_core_dis_uops_0_bits_imm_packed,
  input  [11:0] io_core_dis_uops_0_bits_csr_addr,
  input  [6:0]  io_core_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_0_bits_ldq_idx,
                io_core_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_0_bits_pdst,
                io_core_dis_uops_0_bits_prs1,
                io_core_dis_uops_0_bits_prs2,
                io_core_dis_uops_0_bits_prs3,
  input         io_core_dis_uops_0_bits_prs1_busy,
                io_core_dis_uops_0_bits_prs2_busy,
                io_core_dis_uops_0_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_0_bits_stale_pdst,
  input         io_core_dis_uops_0_bits_exception,
  input  [63:0] io_core_dis_uops_0_bits_exc_cause,
  input         io_core_dis_uops_0_bits_bypassable,
  input  [4:0]  io_core_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_0_bits_mem_size,
  input         io_core_dis_uops_0_bits_mem_signed,
                io_core_dis_uops_0_bits_is_fence,
                io_core_dis_uops_0_bits_is_fencei,
                io_core_dis_uops_0_bits_is_amo,
                io_core_dis_uops_0_bits_uses_ldq,
                io_core_dis_uops_0_bits_uses_stq,
                io_core_dis_uops_0_bits_is_sys_pc2epc,
                io_core_dis_uops_0_bits_is_unique,
                io_core_dis_uops_0_bits_flush_on_commit,
                io_core_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_0_bits_ldst,
                io_core_dis_uops_0_bits_lrs1,
                io_core_dis_uops_0_bits_lrs2,
                io_core_dis_uops_0_bits_lrs3,
  input         io_core_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_0_bits_dst_rtype,
                io_core_dis_uops_0_bits_lrs1_rtype,
                io_core_dis_uops_0_bits_lrs2_rtype,
  input         io_core_dis_uops_0_bits_frs3_en,
                io_core_dis_uops_0_bits_fp_val,
                io_core_dis_uops_0_bits_fp_single,
                io_core_dis_uops_0_bits_xcpt_pf_if,
                io_core_dis_uops_0_bits_xcpt_ae_if,
                io_core_dis_uops_0_bits_xcpt_ma_if,
                io_core_dis_uops_0_bits_bp_debug_if,
                io_core_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_0_bits_debug_fsrc,
                io_core_dis_uops_0_bits_debug_tsrc,
  input         io_core_dis_uops_1_valid,
  input  [6:0]  io_core_dis_uops_1_bits_uopc,
  input  [31:0] io_core_dis_uops_1_bits_inst,
                io_core_dis_uops_1_bits_debug_inst,
  input         io_core_dis_uops_1_bits_is_rvc,
  input  [39:0] io_core_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_1_bits_iq_type,
  input  [9:0]  io_core_dis_uops_1_bits_fu_code,
  input  [3:0]  io_core_dis_uops_1_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_1_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_1_bits_ctrl_op2_sel,
                io_core_dis_uops_1_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_1_bits_ctrl_op_fcn,
  input         io_core_dis_uops_1_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_1_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_1_bits_ctrl_is_load,
                io_core_dis_uops_1_bits_ctrl_is_sta,
                io_core_dis_uops_1_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_1_bits_iw_state,
  input         io_core_dis_uops_1_bits_iw_p1_poisoned,
                io_core_dis_uops_1_bits_iw_p2_poisoned,
                io_core_dis_uops_1_bits_is_br,
                io_core_dis_uops_1_bits_is_jalr,
                io_core_dis_uops_1_bits_is_jal,
                io_core_dis_uops_1_bits_is_sfb,
  input  [15:0] io_core_dis_uops_1_bits_br_mask,
  input  [3:0]  io_core_dis_uops_1_bits_br_tag,
  input  [4:0]  io_core_dis_uops_1_bits_ftq_idx,
  input         io_core_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_1_bits_pc_lob,
  input         io_core_dis_uops_1_bits_taken,
  input  [19:0] io_core_dis_uops_1_bits_imm_packed,
  input  [11:0] io_core_dis_uops_1_bits_csr_addr,
  input  [6:0]  io_core_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_1_bits_ldq_idx,
                io_core_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_1_bits_pdst,
                io_core_dis_uops_1_bits_prs1,
                io_core_dis_uops_1_bits_prs2,
                io_core_dis_uops_1_bits_prs3,
  input         io_core_dis_uops_1_bits_prs1_busy,
                io_core_dis_uops_1_bits_prs2_busy,
                io_core_dis_uops_1_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_1_bits_stale_pdst,
  input         io_core_dis_uops_1_bits_exception,
  input  [63:0] io_core_dis_uops_1_bits_exc_cause,
  input         io_core_dis_uops_1_bits_bypassable,
  input  [4:0]  io_core_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_1_bits_mem_size,
  input         io_core_dis_uops_1_bits_mem_signed,
                io_core_dis_uops_1_bits_is_fence,
                io_core_dis_uops_1_bits_is_fencei,
                io_core_dis_uops_1_bits_is_amo,
                io_core_dis_uops_1_bits_uses_ldq,
                io_core_dis_uops_1_bits_uses_stq,
                io_core_dis_uops_1_bits_is_sys_pc2epc,
                io_core_dis_uops_1_bits_is_unique,
                io_core_dis_uops_1_bits_flush_on_commit,
                io_core_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_1_bits_ldst,
                io_core_dis_uops_1_bits_lrs1,
                io_core_dis_uops_1_bits_lrs2,
                io_core_dis_uops_1_bits_lrs3,
  input         io_core_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_1_bits_dst_rtype,
                io_core_dis_uops_1_bits_lrs1_rtype,
                io_core_dis_uops_1_bits_lrs2_rtype,
  input         io_core_dis_uops_1_bits_frs3_en,
                io_core_dis_uops_1_bits_fp_val,
                io_core_dis_uops_1_bits_fp_single,
                io_core_dis_uops_1_bits_xcpt_pf_if,
                io_core_dis_uops_1_bits_xcpt_ae_if,
                io_core_dis_uops_1_bits_xcpt_ma_if,
                io_core_dis_uops_1_bits_bp_debug_if,
                io_core_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_1_bits_debug_fsrc,
                io_core_dis_uops_1_bits_debug_tsrc,
  input         io_core_dis_uops_2_valid,
  input  [6:0]  io_core_dis_uops_2_bits_uopc,
  input  [31:0] io_core_dis_uops_2_bits_inst,
                io_core_dis_uops_2_bits_debug_inst,
  input         io_core_dis_uops_2_bits_is_rvc,
  input  [39:0] io_core_dis_uops_2_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_2_bits_iq_type,
  input  [9:0]  io_core_dis_uops_2_bits_fu_code,
  input  [3:0]  io_core_dis_uops_2_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_2_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_2_bits_ctrl_op2_sel,
                io_core_dis_uops_2_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_2_bits_ctrl_op_fcn,
  input         io_core_dis_uops_2_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_2_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_2_bits_ctrl_is_load,
                io_core_dis_uops_2_bits_ctrl_is_sta,
                io_core_dis_uops_2_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_2_bits_iw_state,
  input         io_core_dis_uops_2_bits_iw_p1_poisoned,
                io_core_dis_uops_2_bits_iw_p2_poisoned,
                io_core_dis_uops_2_bits_is_br,
                io_core_dis_uops_2_bits_is_jalr,
                io_core_dis_uops_2_bits_is_jal,
                io_core_dis_uops_2_bits_is_sfb,
  input  [15:0] io_core_dis_uops_2_bits_br_mask,
  input  [3:0]  io_core_dis_uops_2_bits_br_tag,
  input  [4:0]  io_core_dis_uops_2_bits_ftq_idx,
  input         io_core_dis_uops_2_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_2_bits_pc_lob,
  input         io_core_dis_uops_2_bits_taken,
  input  [19:0] io_core_dis_uops_2_bits_imm_packed,
  input  [11:0] io_core_dis_uops_2_bits_csr_addr,
  input  [6:0]  io_core_dis_uops_2_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_2_bits_ldq_idx,
                io_core_dis_uops_2_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_2_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_2_bits_pdst,
                io_core_dis_uops_2_bits_prs1,
                io_core_dis_uops_2_bits_prs2,
                io_core_dis_uops_2_bits_prs3,
  input         io_core_dis_uops_2_bits_prs1_busy,
                io_core_dis_uops_2_bits_prs2_busy,
                io_core_dis_uops_2_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_2_bits_stale_pdst,
  input         io_core_dis_uops_2_bits_exception,
  input  [63:0] io_core_dis_uops_2_bits_exc_cause,
  input         io_core_dis_uops_2_bits_bypassable,
  input  [4:0]  io_core_dis_uops_2_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_2_bits_mem_size,
  input         io_core_dis_uops_2_bits_mem_signed,
                io_core_dis_uops_2_bits_is_fence,
                io_core_dis_uops_2_bits_is_fencei,
                io_core_dis_uops_2_bits_is_amo,
                io_core_dis_uops_2_bits_uses_ldq,
                io_core_dis_uops_2_bits_uses_stq,
                io_core_dis_uops_2_bits_is_sys_pc2epc,
                io_core_dis_uops_2_bits_is_unique,
                io_core_dis_uops_2_bits_flush_on_commit,
                io_core_dis_uops_2_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_2_bits_ldst,
                io_core_dis_uops_2_bits_lrs1,
                io_core_dis_uops_2_bits_lrs2,
                io_core_dis_uops_2_bits_lrs3,
  input         io_core_dis_uops_2_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_2_bits_dst_rtype,
                io_core_dis_uops_2_bits_lrs1_rtype,
                io_core_dis_uops_2_bits_lrs2_rtype,
  input         io_core_dis_uops_2_bits_frs3_en,
                io_core_dis_uops_2_bits_fp_val,
                io_core_dis_uops_2_bits_fp_single,
                io_core_dis_uops_2_bits_xcpt_pf_if,
                io_core_dis_uops_2_bits_xcpt_ae_if,
                io_core_dis_uops_2_bits_xcpt_ma_if,
                io_core_dis_uops_2_bits_bp_debug_if,
                io_core_dis_uops_2_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_2_bits_debug_fsrc,
                io_core_dis_uops_2_bits_debug_tsrc,
  input         io_core_fp_stdata_valid,
  input  [15:0] io_core_fp_stdata_bits_uop_br_mask,
  input  [6:0]  io_core_fp_stdata_bits_uop_rob_idx,
  input  [4:0]  io_core_fp_stdata_bits_uop_stq_idx,
  input  [63:0] io_core_fp_stdata_bits_data,
  input         io_core_commit_valids_0,
                io_core_commit_valids_1,
                io_core_commit_valids_2,
                io_core_commit_uops_0_uses_ldq,
                io_core_commit_uops_0_uses_stq,
                io_core_commit_uops_1_uses_ldq,
                io_core_commit_uops_1_uses_stq,
                io_core_commit_uops_2_uses_ldq,
                io_core_commit_uops_2_uses_stq,
                io_core_commit_load_at_rob_head,
                io_core_fence_dmem,
  input  [15:0] io_core_brupdate_b1_resolve_mask,
                io_core_brupdate_b1_mispredict_mask,
  input  [4:0]  io_core_brupdate_b2_uop_ldq_idx,
                io_core_brupdate_b2_uop_stq_idx,
  input         io_core_brupdate_b2_mispredict,
  input  [6:0]  io_core_rob_head_idx,
  input         io_core_exception,
                io_dmem_req_ready,
                io_dmem_resp_0_valid,
  input  [4:0]  io_dmem_resp_0_bits_uop_ldq_idx,
                io_dmem_resp_0_bits_uop_stq_idx,
  input         io_dmem_resp_0_bits_uop_is_amo,
                io_dmem_resp_0_bits_uop_uses_ldq,
                io_dmem_resp_0_bits_uop_uses_stq,
  input  [63:0] io_dmem_resp_0_bits_data,
  input         io_dmem_resp_0_bits_is_hella,
                io_dmem_nack_0_valid,
  input  [4:0]  io_dmem_nack_0_bits_uop_ldq_idx,
                io_dmem_nack_0_bits_uop_stq_idx,
  input         io_dmem_nack_0_bits_uop_uses_ldq,
                io_dmem_nack_0_bits_uop_uses_stq,
                io_dmem_nack_0_bits_is_hella,
                io_dmem_release_valid,
  input  [31:0] io_dmem_release_bits_address,
  input         io_dmem_ordered,
                io_hellacache_req_valid,
  input  [39:0] io_hellacache_req_bits_addr,
  input         io_hellacache_s1_kill,
  output        io_ptw_req_valid,
                io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  output        io_core_exe_0_iresp_valid,
  output [6:0]  io_core_exe_0_iresp_bits_uop_rob_idx,
                io_core_exe_0_iresp_bits_uop_pdst,
  output        io_core_exe_0_iresp_bits_uop_is_amo,
                io_core_exe_0_iresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_iresp_bits_uop_dst_rtype,
  output [63:0] io_core_exe_0_iresp_bits_data,
  output        io_core_exe_0_fresp_valid,
  output [6:0]  io_core_exe_0_fresp_bits_uop_uopc,
  output [15:0] io_core_exe_0_fresp_bits_uop_br_mask,
  output [6:0]  io_core_exe_0_fresp_bits_uop_rob_idx,
  output [4:0]  io_core_exe_0_fresp_bits_uop_stq_idx,
  output [6:0]  io_core_exe_0_fresp_bits_uop_pdst,
  output [1:0]  io_core_exe_0_fresp_bits_uop_mem_size,
  output        io_core_exe_0_fresp_bits_uop_is_amo,
                io_core_exe_0_fresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_fresp_bits_uop_dst_rtype,
  output        io_core_exe_0_fresp_bits_uop_fp_val,
  output [64:0] io_core_exe_0_fresp_bits_data,
  output [4:0]  io_core_dis_ldq_idx_0,
                io_core_dis_ldq_idx_1,
                io_core_dis_ldq_idx_2,
                io_core_dis_stq_idx_0,
                io_core_dis_stq_idx_1,
                io_core_dis_stq_idx_2,
  output        io_core_ldq_full_0,
                io_core_ldq_full_1,
                io_core_ldq_full_2,
                io_core_stq_full_0,
                io_core_stq_full_1,
                io_core_stq_full_2,
                io_core_fp_stdata_ready,
                io_core_clr_bsy_0_valid,
  output [6:0]  io_core_clr_bsy_0_bits,
  output        io_core_clr_bsy_1_valid,
  output [6:0]  io_core_clr_bsy_1_bits,
  output        io_core_spec_ld_wakeup_0_valid,
  output [6:0]  io_core_spec_ld_wakeup_0_bits,
  output        io_core_ld_miss,
                io_core_fencei_rdy,
                io_core_lxcpt_valid,
  output [15:0] io_core_lxcpt_bits_uop_br_mask,
  output [6:0]  io_core_lxcpt_bits_uop_rob_idx,
  output [4:0]  io_core_lxcpt_bits_cause,
  output [39:0] io_core_lxcpt_bits_badvaddr,
  output        io_dmem_req_valid,
                io_dmem_req_bits_0_valid,
  output [6:0]  io_dmem_req_bits_0_bits_uop_uopc,
  output [31:0] io_dmem_req_bits_0_bits_uop_inst,
                io_dmem_req_bits_0_bits_uop_debug_inst,
  output        io_dmem_req_bits_0_bits_uop_is_rvc,
  output [39:0] io_dmem_req_bits_0_bits_uop_debug_pc,
  output [2:0]  io_dmem_req_bits_0_bits_uop_iq_type,
  output [9:0]  io_dmem_req_bits_0_bits_uop_fu_code,
  output [3:0]  io_dmem_req_bits_0_bits_uop_ctrl_br_type,
  output [1:0]  io_dmem_req_bits_0_bits_uop_ctrl_op1_sel,
  output [2:0]  io_dmem_req_bits_0_bits_uop_ctrl_op2_sel,
                io_dmem_req_bits_0_bits_uop_ctrl_imm_sel,
  output [3:0]  io_dmem_req_bits_0_bits_uop_ctrl_op_fcn,
  output        io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd,
  output        io_dmem_req_bits_0_bits_uop_ctrl_is_load,
                io_dmem_req_bits_0_bits_uop_ctrl_is_sta,
                io_dmem_req_bits_0_bits_uop_ctrl_is_std,
  output [1:0]  io_dmem_req_bits_0_bits_uop_iw_state,
  output        io_dmem_req_bits_0_bits_uop_iw_p1_poisoned,
                io_dmem_req_bits_0_bits_uop_iw_p2_poisoned,
                io_dmem_req_bits_0_bits_uop_is_br,
                io_dmem_req_bits_0_bits_uop_is_jalr,
                io_dmem_req_bits_0_bits_uop_is_jal,
                io_dmem_req_bits_0_bits_uop_is_sfb,
  output [15:0] io_dmem_req_bits_0_bits_uop_br_mask,
  output [3:0]  io_dmem_req_bits_0_bits_uop_br_tag,
  output [4:0]  io_dmem_req_bits_0_bits_uop_ftq_idx,
  output        io_dmem_req_bits_0_bits_uop_edge_inst,
  output [5:0]  io_dmem_req_bits_0_bits_uop_pc_lob,
  output        io_dmem_req_bits_0_bits_uop_taken,
  output [19:0] io_dmem_req_bits_0_bits_uop_imm_packed,
  output [11:0] io_dmem_req_bits_0_bits_uop_csr_addr,
  output [6:0]  io_dmem_req_bits_0_bits_uop_rob_idx,
  output [4:0]  io_dmem_req_bits_0_bits_uop_ldq_idx,
                io_dmem_req_bits_0_bits_uop_stq_idx,
  output [1:0]  io_dmem_req_bits_0_bits_uop_rxq_idx,
  output [6:0]  io_dmem_req_bits_0_bits_uop_pdst,
                io_dmem_req_bits_0_bits_uop_prs1,
                io_dmem_req_bits_0_bits_uop_prs2,
                io_dmem_req_bits_0_bits_uop_prs3,
  output [4:0]  io_dmem_req_bits_0_bits_uop_ppred,
  output        io_dmem_req_bits_0_bits_uop_prs1_busy,
                io_dmem_req_bits_0_bits_uop_prs2_busy,
                io_dmem_req_bits_0_bits_uop_prs3_busy,
                io_dmem_req_bits_0_bits_uop_ppred_busy,
  output [6:0]  io_dmem_req_bits_0_bits_uop_stale_pdst,
  output        io_dmem_req_bits_0_bits_uop_exception,
  output [63:0] io_dmem_req_bits_0_bits_uop_exc_cause,
  output        io_dmem_req_bits_0_bits_uop_bypassable,
  output [4:0]  io_dmem_req_bits_0_bits_uop_mem_cmd,
  output [1:0]  io_dmem_req_bits_0_bits_uop_mem_size,
  output        io_dmem_req_bits_0_bits_uop_mem_signed,
                io_dmem_req_bits_0_bits_uop_is_fence,
                io_dmem_req_bits_0_bits_uop_is_fencei,
                io_dmem_req_bits_0_bits_uop_is_amo,
                io_dmem_req_bits_0_bits_uop_uses_ldq,
                io_dmem_req_bits_0_bits_uop_uses_stq,
                io_dmem_req_bits_0_bits_uop_is_sys_pc2epc,
                io_dmem_req_bits_0_bits_uop_is_unique,
                io_dmem_req_bits_0_bits_uop_flush_on_commit,
                io_dmem_req_bits_0_bits_uop_ldst_is_rs1,
  output [5:0]  io_dmem_req_bits_0_bits_uop_ldst,
                io_dmem_req_bits_0_bits_uop_lrs1,
                io_dmem_req_bits_0_bits_uop_lrs2,
                io_dmem_req_bits_0_bits_uop_lrs3,
  output        io_dmem_req_bits_0_bits_uop_ldst_val,
  output [1:0]  io_dmem_req_bits_0_bits_uop_dst_rtype,
                io_dmem_req_bits_0_bits_uop_lrs1_rtype,
                io_dmem_req_bits_0_bits_uop_lrs2_rtype,
  output        io_dmem_req_bits_0_bits_uop_frs3_en,
                io_dmem_req_bits_0_bits_uop_fp_val,
                io_dmem_req_bits_0_bits_uop_fp_single,
                io_dmem_req_bits_0_bits_uop_xcpt_pf_if,
                io_dmem_req_bits_0_bits_uop_xcpt_ae_if,
                io_dmem_req_bits_0_bits_uop_xcpt_ma_if,
                io_dmem_req_bits_0_bits_uop_bp_debug_if,
                io_dmem_req_bits_0_bits_uop_bp_xcpt_if,
  output [1:0]  io_dmem_req_bits_0_bits_uop_debug_fsrc,
                io_dmem_req_bits_0_bits_uop_debug_tsrc,
  output [39:0] io_dmem_req_bits_0_bits_addr,
  output [63:0] io_dmem_req_bits_0_bits_data,
  output        io_dmem_req_bits_0_bits_is_hella,
                io_dmem_s1_kill_0,
  output [15:0] io_dmem_brupdate_b1_resolve_mask,
                io_dmem_brupdate_b1_mispredict_mask,
  output        io_dmem_exception,
                io_dmem_release_ready,
                io_dmem_force_order,
                io_hellacache_req_ready,
                io_hellacache_s2_nack,
                io_hellacache_resp_valid,
  output [63:0] io_hellacache_resp_bits_data,
  output        io_hellacache_s2_xcpt_ae_ld
);

  wire              _GEN;	// lsu.scala:1527:34, :1533:38, :1550:43, :1553:38, :1560:40, :1576:42
  wire              store_needs_order;	// lsu.scala:1495:3, :1496:64
  wire              nacking_loads_23;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_22;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_21;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_20;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_19;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_18;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_17;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_16;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_15;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_14;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_13;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_12;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_11;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_10;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_9;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_8;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_7;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_6;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_5;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_4;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_3;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_2;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_1;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_0;	// lsu.scala:1284:5, :1287:7
  wire              block_load_wakeup;	// lsu.scala:1199:80, :1210:43, :1211:25
  wire              _GEN_0;	// lsu.scala:820:26
  wire              _GEN_1;	// lsu.scala:803:26
  reg               mem_xcpt_valids_0;	// lsu.scala:667:32
  wire              _will_fire_store_commit_0_T_2;	// lsu.scala:538:31
  wire [4:0]        _forwarding_age_logic_0_io_forwarding_idx;	// lsu.scala:1178:57
  wire              _dtlb_io_miss_rdy;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_miss;	// lsu.scala:249:20
  wire [31:0]       _dtlb_io_resp_0_paddr;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_pf_ld;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_pf_st;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ae_ld;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ae_st;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ma_ld;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ma_st;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_cacheable;	// lsu.scala:249:20
  reg               ldq_0_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_0_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_0_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_0_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_0_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_0_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_0_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_0_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_0_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_0_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_0_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_0_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_0_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_0_bits_executed;	// lsu.scala:210:16
  reg               ldq_0_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_0_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_0_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_0_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_0_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_1_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_1_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_1_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_1_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_1_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_1_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_1_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_1_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_1_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_1_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_1_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_1_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_1_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_1_bits_executed;	// lsu.scala:210:16
  reg               ldq_1_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_1_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_1_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_1_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_1_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_2_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_2_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_2_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_2_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_2_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_2_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_2_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_2_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_2_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_2_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_2_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_2_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_2_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_2_bits_executed;	// lsu.scala:210:16
  reg               ldq_2_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_2_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_2_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_2_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_2_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_3_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_3_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_3_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_3_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_3_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_3_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_3_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_3_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_3_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_3_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_3_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_3_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_3_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_3_bits_executed;	// lsu.scala:210:16
  reg               ldq_3_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_3_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_3_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_3_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_3_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_4_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_4_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_4_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_4_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_4_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_4_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_4_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_4_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_4_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_4_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_4_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_4_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_4_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_4_bits_executed;	// lsu.scala:210:16
  reg               ldq_4_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_4_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_4_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_4_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_4_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_5_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_5_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_5_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_5_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_5_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_5_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_5_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_5_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_5_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_5_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_5_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_5_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_5_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_5_bits_executed;	// lsu.scala:210:16
  reg               ldq_5_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_5_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_5_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_5_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_5_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_6_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_6_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_6_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_6_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_6_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_6_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_6_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_6_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_6_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_6_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_6_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_6_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_6_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_6_bits_executed;	// lsu.scala:210:16
  reg               ldq_6_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_6_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_6_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_6_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_6_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_7_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_7_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_7_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_7_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_7_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_7_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_7_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_7_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_7_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_7_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_7_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_7_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_7_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_7_bits_executed;	// lsu.scala:210:16
  reg               ldq_7_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_7_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_7_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_7_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_7_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_8_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_8_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_8_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_8_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_8_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_8_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_8_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_8_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_8_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_8_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_8_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_8_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_8_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_8_bits_executed;	// lsu.scala:210:16
  reg               ldq_8_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_8_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_8_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_8_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_8_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_9_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_9_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_9_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_9_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_9_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_9_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_9_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_9_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_9_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_9_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_9_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_9_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_9_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_9_bits_executed;	// lsu.scala:210:16
  reg               ldq_9_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_9_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_9_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_9_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_9_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_10_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_10_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_10_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_10_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_10_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_10_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_10_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_10_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_10_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_10_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_10_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_10_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_10_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_10_bits_executed;	// lsu.scala:210:16
  reg               ldq_10_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_10_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_10_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_10_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_10_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_11_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_11_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_11_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_11_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_11_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_11_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_11_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_11_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_11_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_11_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_11_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_11_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_11_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_11_bits_executed;	// lsu.scala:210:16
  reg               ldq_11_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_11_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_11_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_11_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_11_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_12_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_12_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_12_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_12_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_12_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_12_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_12_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_12_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_12_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_12_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_12_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_12_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_12_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_12_bits_executed;	// lsu.scala:210:16
  reg               ldq_12_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_12_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_12_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_12_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_12_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_13_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_13_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_13_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_13_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_13_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_13_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_13_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_13_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_13_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_13_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_13_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_13_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_13_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_13_bits_executed;	// lsu.scala:210:16
  reg               ldq_13_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_13_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_13_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_13_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_13_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_14_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_14_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_14_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_14_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_14_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_14_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_14_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_14_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_14_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_14_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_14_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_14_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_14_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_14_bits_executed;	// lsu.scala:210:16
  reg               ldq_14_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_14_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_14_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_14_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_14_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_15_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_15_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_15_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_15_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_15_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_15_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_15_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_15_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_15_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_15_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_15_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_15_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_15_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_15_bits_executed;	// lsu.scala:210:16
  reg               ldq_15_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_15_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_15_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_15_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_15_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_16_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_16_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_16_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_16_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_16_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_16_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_16_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_16_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_16_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_16_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_16_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_16_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_16_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_16_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_16_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_16_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_16_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_16_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_16_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_16_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_16_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_16_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_16_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_16_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_16_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_16_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_16_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_16_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_16_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_16_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_16_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_16_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_16_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_16_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_16_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_16_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_16_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_16_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_16_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_16_bits_executed;	// lsu.scala:210:16
  reg               ldq_16_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_16_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_16_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_16_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_16_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_16_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_16_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_17_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_17_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_17_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_17_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_17_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_17_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_17_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_17_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_17_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_17_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_17_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_17_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_17_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_17_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_17_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_17_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_17_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_17_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_17_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_17_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_17_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_17_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_17_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_17_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_17_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_17_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_17_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_17_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_17_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_17_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_17_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_17_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_17_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_17_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_17_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_17_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_17_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_17_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_17_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_17_bits_executed;	// lsu.scala:210:16
  reg               ldq_17_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_17_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_17_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_17_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_17_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_17_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_17_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_18_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_18_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_18_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_18_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_18_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_18_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_18_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_18_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_18_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_18_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_18_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_18_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_18_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_18_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_18_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_18_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_18_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_18_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_18_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_18_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_18_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_18_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_18_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_18_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_18_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_18_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_18_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_18_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_18_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_18_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_18_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_18_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_18_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_18_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_18_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_18_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_18_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_18_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_18_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_18_bits_executed;	// lsu.scala:210:16
  reg               ldq_18_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_18_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_18_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_18_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_18_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_18_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_18_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_19_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_19_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_19_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_19_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_19_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_19_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_19_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_19_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_19_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_19_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_19_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_19_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_19_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_19_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_19_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_19_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_19_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_19_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_19_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_19_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_19_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_19_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_19_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_19_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_19_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_19_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_19_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_19_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_19_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_19_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_19_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_19_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_19_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_19_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_19_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_19_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_19_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_19_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_19_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_19_bits_executed;	// lsu.scala:210:16
  reg               ldq_19_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_19_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_19_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_19_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_19_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_19_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_19_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_20_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_20_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_20_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_20_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_20_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_20_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_20_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_20_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_20_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_20_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_20_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_20_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_20_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_20_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_20_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_20_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_20_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_20_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_20_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_20_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_20_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_20_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_20_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_20_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_20_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_20_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_20_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_20_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_20_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_20_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_20_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_20_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_20_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_20_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_20_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_20_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_20_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_20_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_20_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_20_bits_executed;	// lsu.scala:210:16
  reg               ldq_20_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_20_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_20_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_20_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_20_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_20_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_20_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_21_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_21_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_21_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_21_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_21_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_21_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_21_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_21_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_21_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_21_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_21_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_21_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_21_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_21_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_21_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_21_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_21_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_21_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_21_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_21_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_21_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_21_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_21_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_21_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_21_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_21_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_21_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_21_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_21_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_21_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_21_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_21_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_21_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_21_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_21_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_21_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_21_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_21_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_21_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_21_bits_executed;	// lsu.scala:210:16
  reg               ldq_21_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_21_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_21_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_21_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_21_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_21_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_21_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_22_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_22_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_22_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_22_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_22_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_22_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_22_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_22_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_22_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_22_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_22_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_22_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_22_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_22_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_22_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_22_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_22_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_22_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_22_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_22_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_22_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_22_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_22_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_22_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_22_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_22_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_22_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_22_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_22_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_22_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_22_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_22_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_22_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_22_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_22_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_22_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_22_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_22_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_22_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_22_bits_executed;	// lsu.scala:210:16
  reg               ldq_22_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_22_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_22_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_22_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_22_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_22_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_22_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_23_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_23_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_23_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_23_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_23_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_23_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_23_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_23_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_23_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_23_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_23_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_23_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [15:0]       ldq_23_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_23_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_23_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_23_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_23_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_23_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [6:0]        ldq_23_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_23_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [4:0]        ldq_23_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_23_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_23_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_23_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_23_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_23_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_23_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_23_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_23_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_23_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_23_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_23_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_23_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_23_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_23_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_23_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_23_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_23_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_23_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_23_bits_executed;	// lsu.scala:210:16
  reg               ldq_23_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_23_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_23_bits_observed;	// lsu.scala:210:16
  reg  [23:0]       ldq_23_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [4:0]        ldq_23_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_23_bits_forward_std_val;	// lsu.scala:210:16
  reg  [4:0]        ldq_23_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               stq_0_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_0_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_0_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_0_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_0_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_0_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_0_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_0_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_0_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_0_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_0_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_0_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_0_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_0_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_0_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_0_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_0_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_0_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_0_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_0_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_0_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_0_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_0_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_0_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_0_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_0_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_0_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_0_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_0_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_0_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_0_bits_data_bits;	// lsu.scala:211:16
  reg               stq_0_bits_committed;	// lsu.scala:211:16
  reg               stq_0_bits_succeeded;	// lsu.scala:211:16
  reg               stq_1_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_1_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_1_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_1_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_1_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_1_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_1_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_1_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_1_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_1_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_1_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_1_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_1_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_1_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_1_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_1_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_1_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_1_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_1_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_1_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_1_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_1_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_1_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_1_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_1_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_1_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_1_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_1_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_1_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_1_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_1_bits_data_bits;	// lsu.scala:211:16
  reg               stq_1_bits_committed;	// lsu.scala:211:16
  reg               stq_1_bits_succeeded;	// lsu.scala:211:16
  reg               stq_2_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_2_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_2_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_2_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_2_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_2_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_2_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_2_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_2_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_2_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_2_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_2_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_2_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_2_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_2_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_2_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_2_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_2_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_2_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_2_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_2_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_2_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_2_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_2_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_2_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_2_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_2_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_2_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_2_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_2_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_2_bits_data_bits;	// lsu.scala:211:16
  reg               stq_2_bits_committed;	// lsu.scala:211:16
  reg               stq_2_bits_succeeded;	// lsu.scala:211:16
  reg               stq_3_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_3_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_3_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_3_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_3_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_3_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_3_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_3_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_3_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_3_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_3_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_3_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_3_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_3_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_3_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_3_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_3_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_3_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_3_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_3_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_3_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_3_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_3_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_3_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_3_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_3_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_3_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_3_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_3_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_3_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_3_bits_data_bits;	// lsu.scala:211:16
  reg               stq_3_bits_committed;	// lsu.scala:211:16
  reg               stq_3_bits_succeeded;	// lsu.scala:211:16
  reg               stq_4_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_4_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_4_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_4_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_4_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_4_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_4_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_4_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_4_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_4_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_4_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_4_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_4_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_4_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_4_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_4_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_4_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_4_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_4_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_4_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_4_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_4_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_4_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_4_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_4_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_4_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_4_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_4_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_4_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_4_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_4_bits_data_bits;	// lsu.scala:211:16
  reg               stq_4_bits_committed;	// lsu.scala:211:16
  reg               stq_4_bits_succeeded;	// lsu.scala:211:16
  reg               stq_5_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_5_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_5_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_5_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_5_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_5_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_5_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_5_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_5_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_5_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_5_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_5_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_5_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_5_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_5_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_5_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_5_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_5_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_5_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_5_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_5_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_5_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_5_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_5_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_5_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_5_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_5_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_5_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_5_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_5_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_5_bits_data_bits;	// lsu.scala:211:16
  reg               stq_5_bits_committed;	// lsu.scala:211:16
  reg               stq_5_bits_succeeded;	// lsu.scala:211:16
  reg               stq_6_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_6_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_6_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_6_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_6_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_6_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_6_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_6_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_6_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_6_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_6_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_6_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_6_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_6_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_6_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_6_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_6_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_6_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_6_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_6_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_6_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_6_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_6_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_6_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_6_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_6_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_6_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_6_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_6_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_6_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_6_bits_data_bits;	// lsu.scala:211:16
  reg               stq_6_bits_committed;	// lsu.scala:211:16
  reg               stq_6_bits_succeeded;	// lsu.scala:211:16
  reg               stq_7_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_7_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_7_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_7_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_7_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_7_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_7_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_7_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_7_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_7_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_7_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_7_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_7_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_7_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_7_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_7_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_7_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_7_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_7_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_7_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_7_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_7_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_7_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_7_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_7_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_7_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_7_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_7_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_7_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_7_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_7_bits_data_bits;	// lsu.scala:211:16
  reg               stq_7_bits_committed;	// lsu.scala:211:16
  reg               stq_7_bits_succeeded;	// lsu.scala:211:16
  reg               stq_8_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_8_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_8_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_8_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_8_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_8_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_8_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_8_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_8_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_8_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_8_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_8_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_8_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_8_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_8_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_8_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_8_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_8_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_8_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_8_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_8_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_8_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_8_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_8_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_8_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_8_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_8_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_8_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_8_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_8_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_8_bits_data_bits;	// lsu.scala:211:16
  reg               stq_8_bits_committed;	// lsu.scala:211:16
  reg               stq_8_bits_succeeded;	// lsu.scala:211:16
  reg               stq_9_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_9_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_9_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_9_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_9_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_9_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_9_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_9_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_9_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_9_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_9_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_9_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_9_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_9_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_9_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_9_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_9_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_9_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_9_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_9_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_9_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_9_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_9_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_9_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_9_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_9_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_9_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_9_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_9_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_9_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_9_bits_data_bits;	// lsu.scala:211:16
  reg               stq_9_bits_committed;	// lsu.scala:211:16
  reg               stq_9_bits_succeeded;	// lsu.scala:211:16
  reg               stq_10_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_10_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_10_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_10_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_10_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_10_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_10_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_10_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_10_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_10_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_10_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_10_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_10_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_10_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_10_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_10_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_10_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_10_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_10_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_10_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_10_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_10_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_10_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_10_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_10_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_10_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_10_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_10_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_10_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_10_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_10_bits_data_bits;	// lsu.scala:211:16
  reg               stq_10_bits_committed;	// lsu.scala:211:16
  reg               stq_10_bits_succeeded;	// lsu.scala:211:16
  reg               stq_11_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_11_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_11_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_11_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_11_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_11_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_11_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_11_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_11_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_11_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_11_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_11_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_11_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_11_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_11_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_11_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_11_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_11_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_11_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_11_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_11_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_11_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_11_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_11_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_11_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_11_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_11_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_11_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_11_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_11_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_11_bits_data_bits;	// lsu.scala:211:16
  reg               stq_11_bits_committed;	// lsu.scala:211:16
  reg               stq_11_bits_succeeded;	// lsu.scala:211:16
  reg               stq_12_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_12_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_12_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_12_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_12_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_12_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_12_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_12_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_12_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_12_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_12_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_12_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_12_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_12_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_12_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_12_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_12_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_12_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_12_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_12_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_12_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_12_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_12_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_12_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_12_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_12_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_12_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_12_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_12_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_12_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_12_bits_data_bits;	// lsu.scala:211:16
  reg               stq_12_bits_committed;	// lsu.scala:211:16
  reg               stq_12_bits_succeeded;	// lsu.scala:211:16
  reg               stq_13_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_13_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_13_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_13_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_13_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_13_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_13_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_13_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_13_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_13_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_13_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_13_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_13_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_13_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_13_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_13_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_13_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_13_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_13_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_13_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_13_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_13_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_13_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_13_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_13_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_13_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_13_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_13_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_13_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_13_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_13_bits_data_bits;	// lsu.scala:211:16
  reg               stq_13_bits_committed;	// lsu.scala:211:16
  reg               stq_13_bits_succeeded;	// lsu.scala:211:16
  reg               stq_14_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_14_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_14_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_14_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_14_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_14_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_14_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_14_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_14_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_14_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_14_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_14_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_14_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_14_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_14_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_14_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_14_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_14_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_14_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_14_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_14_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_14_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_14_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_14_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_14_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_14_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_14_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_14_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_14_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_14_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_14_bits_data_bits;	// lsu.scala:211:16
  reg               stq_14_bits_committed;	// lsu.scala:211:16
  reg               stq_14_bits_succeeded;	// lsu.scala:211:16
  reg               stq_15_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_15_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_15_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_15_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_15_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_15_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_15_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_15_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_15_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_15_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_15_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_15_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_15_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_15_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_15_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_15_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_15_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_15_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_15_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_15_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_15_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_15_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_15_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_15_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_15_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_15_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_15_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_15_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_15_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_15_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_15_bits_data_bits;	// lsu.scala:211:16
  reg               stq_15_bits_committed;	// lsu.scala:211:16
  reg               stq_15_bits_succeeded;	// lsu.scala:211:16
  reg               stq_16_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_16_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_16_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_16_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_16_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_16_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_16_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_16_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_16_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_16_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_16_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_16_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_16_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_16_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_16_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_16_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_16_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_16_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_16_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_16_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_16_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_16_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_16_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_16_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_16_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_16_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_16_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_16_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_16_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_16_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_16_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_16_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_16_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_16_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_16_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_16_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_16_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_16_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_16_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_16_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_16_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_16_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_16_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_16_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_16_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_16_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_16_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_16_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_16_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_16_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_16_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_16_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_16_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_16_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_16_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_16_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_16_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_16_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_16_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_16_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_16_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_16_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_16_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_16_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_16_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_16_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_16_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_16_bits_data_bits;	// lsu.scala:211:16
  reg               stq_16_bits_committed;	// lsu.scala:211:16
  reg               stq_16_bits_succeeded;	// lsu.scala:211:16
  reg               stq_17_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_17_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_17_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_17_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_17_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_17_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_17_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_17_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_17_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_17_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_17_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_17_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_17_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_17_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_17_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_17_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_17_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_17_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_17_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_17_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_17_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_17_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_17_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_17_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_17_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_17_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_17_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_17_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_17_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_17_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_17_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_17_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_17_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_17_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_17_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_17_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_17_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_17_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_17_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_17_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_17_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_17_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_17_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_17_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_17_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_17_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_17_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_17_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_17_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_17_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_17_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_17_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_17_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_17_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_17_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_17_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_17_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_17_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_17_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_17_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_17_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_17_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_17_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_17_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_17_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_17_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_17_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_17_bits_data_bits;	// lsu.scala:211:16
  reg               stq_17_bits_committed;	// lsu.scala:211:16
  reg               stq_17_bits_succeeded;	// lsu.scala:211:16
  reg               stq_18_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_18_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_18_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_18_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_18_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_18_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_18_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_18_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_18_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_18_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_18_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_18_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_18_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_18_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_18_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_18_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_18_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_18_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_18_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_18_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_18_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_18_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_18_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_18_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_18_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_18_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_18_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_18_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_18_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_18_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_18_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_18_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_18_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_18_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_18_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_18_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_18_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_18_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_18_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_18_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_18_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_18_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_18_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_18_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_18_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_18_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_18_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_18_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_18_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_18_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_18_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_18_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_18_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_18_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_18_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_18_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_18_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_18_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_18_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_18_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_18_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_18_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_18_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_18_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_18_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_18_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_18_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_18_bits_data_bits;	// lsu.scala:211:16
  reg               stq_18_bits_committed;	// lsu.scala:211:16
  reg               stq_18_bits_succeeded;	// lsu.scala:211:16
  reg               stq_19_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_19_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_19_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_19_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_19_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_19_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_19_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_19_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_19_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_19_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_19_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_19_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_19_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_19_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_19_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_19_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_19_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_19_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_19_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_19_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_19_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_19_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_19_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_19_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_19_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_19_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_19_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_19_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_19_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_19_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_19_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_19_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_19_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_19_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_19_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_19_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_19_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_19_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_19_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_19_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_19_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_19_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_19_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_19_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_19_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_19_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_19_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_19_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_19_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_19_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_19_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_19_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_19_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_19_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_19_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_19_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_19_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_19_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_19_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_19_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_19_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_19_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_19_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_19_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_19_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_19_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_19_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_19_bits_data_bits;	// lsu.scala:211:16
  reg               stq_19_bits_committed;	// lsu.scala:211:16
  reg               stq_19_bits_succeeded;	// lsu.scala:211:16
  reg               stq_20_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_20_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_20_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_20_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_20_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_20_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_20_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_20_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_20_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_20_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_20_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_20_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_20_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_20_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_20_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_20_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_20_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_20_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_20_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_20_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_20_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_20_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_20_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_20_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_20_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_20_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_20_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_20_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_20_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_20_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_20_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_20_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_20_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_20_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_20_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_20_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_20_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_20_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_20_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_20_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_20_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_20_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_20_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_20_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_20_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_20_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_20_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_20_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_20_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_20_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_20_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_20_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_20_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_20_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_20_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_20_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_20_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_20_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_20_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_20_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_20_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_20_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_20_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_20_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_20_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_20_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_20_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_20_bits_data_bits;	// lsu.scala:211:16
  reg               stq_20_bits_committed;	// lsu.scala:211:16
  reg               stq_20_bits_succeeded;	// lsu.scala:211:16
  reg               stq_21_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_21_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_21_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_21_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_21_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_21_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_21_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_21_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_21_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_21_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_21_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_21_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_21_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_21_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_21_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_21_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_21_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_21_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_21_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_21_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_21_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_21_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_21_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_21_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_21_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_21_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_21_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_21_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_21_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_21_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_21_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_21_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_21_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_21_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_21_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_21_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_21_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_21_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_21_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_21_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_21_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_21_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_21_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_21_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_21_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_21_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_21_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_21_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_21_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_21_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_21_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_21_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_21_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_21_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_21_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_21_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_21_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_21_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_21_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_21_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_21_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_21_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_21_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_21_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_21_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_21_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_21_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_21_bits_data_bits;	// lsu.scala:211:16
  reg               stq_21_bits_committed;	// lsu.scala:211:16
  reg               stq_21_bits_succeeded;	// lsu.scala:211:16
  reg               stq_22_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_22_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_22_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_22_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_22_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_22_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_22_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_22_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_22_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_22_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_22_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_22_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_22_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_22_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_22_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_22_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_22_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_22_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_22_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_22_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_22_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_22_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_22_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_22_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_22_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_22_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_22_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_22_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_22_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_22_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_22_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_22_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_22_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_22_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_22_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_22_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_22_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_22_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_22_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_22_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_22_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_22_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_22_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_22_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_22_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_22_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_22_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_22_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_22_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_22_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_22_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_22_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_22_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_22_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_22_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_22_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_22_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_22_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_22_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_22_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_22_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_22_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_22_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_22_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_22_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_22_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_22_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_22_bits_data_bits;	// lsu.scala:211:16
  reg               stq_22_bits_committed;	// lsu.scala:211:16
  reg               stq_22_bits_succeeded;	// lsu.scala:211:16
  reg               stq_23_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_23_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_23_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_23_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_23_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_23_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_23_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_23_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_23_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_23_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_23_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_23_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_23_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_23_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_23_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_23_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_23_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_23_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [15:0]       stq_23_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_23_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_23_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_23_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_23_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_23_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_23_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_23_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [6:0]        stq_23_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_23_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [4:0]        stq_23_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_23_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_23_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_23_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_23_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_23_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_23_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_23_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_23_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_23_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_23_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_23_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_23_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_23_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_23_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_23_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_23_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_23_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_23_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_23_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_23_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_23_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_23_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_23_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_23_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_23_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_23_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_23_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_23_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_23_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_23_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_23_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_23_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_23_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_23_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_23_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_23_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_23_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_23_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_23_bits_data_bits;	// lsu.scala:211:16
  reg               stq_23_bits_committed;	// lsu.scala:211:16
  reg               stq_23_bits_succeeded;	// lsu.scala:211:16
  reg  [4:0]        ldq_head;	// lsu.scala:215:29
  reg  [4:0]        ldq_tail;	// lsu.scala:216:29
  reg  [4:0]        stq_head;	// lsu.scala:217:29
  reg  [4:0]        stq_tail;	// lsu.scala:218:29
  reg  [4:0]        stq_commit_head;	// lsu.scala:219:29
  reg  [4:0]        stq_execute_head;	// lsu.scala:220:29
  wire [31:0]       _GEN_2 =
    {{stq_0_valid},
     {stq_0_valid},
     {stq_0_valid},
     {stq_0_valid},
     {stq_0_valid},
     {stq_0_valid},
     {stq_0_valid},
     {stq_0_valid},
     {stq_23_valid},
     {stq_22_valid},
     {stq_21_valid},
     {stq_20_valid},
     {stq_19_valid},
     {stq_18_valid},
     {stq_17_valid},
     {stq_16_valid},
     {stq_15_valid},
     {stq_14_valid},
     {stq_13_valid},
     {stq_12_valid},
     {stq_11_valid},
     {stq_10_valid},
     {stq_9_valid},
     {stq_8_valid},
     {stq_7_valid},
     {stq_6_valid},
     {stq_5_valid},
     {stq_4_valid},
     {stq_3_valid},
     {stq_2_valid},
     {stq_1_valid},
     {stq_0_valid}};	// lsu.scala:211:16, :224:42
  wire              _GEN_3 = _GEN_2[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [31:0][6:0]  _GEN_4 =
    {{stq_0_bits_uop_uopc},
     {stq_0_bits_uop_uopc},
     {stq_0_bits_uop_uopc},
     {stq_0_bits_uop_uopc},
     {stq_0_bits_uop_uopc},
     {stq_0_bits_uop_uopc},
     {stq_0_bits_uop_uopc},
     {stq_0_bits_uop_uopc},
     {stq_23_bits_uop_uopc},
     {stq_22_bits_uop_uopc},
     {stq_21_bits_uop_uopc},
     {stq_20_bits_uop_uopc},
     {stq_19_bits_uop_uopc},
     {stq_18_bits_uop_uopc},
     {stq_17_bits_uop_uopc},
     {stq_16_bits_uop_uopc},
     {stq_15_bits_uop_uopc},
     {stq_14_bits_uop_uopc},
     {stq_13_bits_uop_uopc},
     {stq_12_bits_uop_uopc},
     {stq_11_bits_uop_uopc},
     {stq_10_bits_uop_uopc},
     {stq_9_bits_uop_uopc},
     {stq_8_bits_uop_uopc},
     {stq_7_bits_uop_uopc},
     {stq_6_bits_uop_uopc},
     {stq_5_bits_uop_uopc},
     {stq_4_bits_uop_uopc},
     {stq_3_bits_uop_uopc},
     {stq_2_bits_uop_uopc},
     {stq_1_bits_uop_uopc},
     {stq_0_bits_uop_uopc}};	// lsu.scala:211:16, :224:42
  wire [31:0][31:0] _GEN_5 =
    {{stq_0_bits_uop_inst},
     {stq_0_bits_uop_inst},
     {stq_0_bits_uop_inst},
     {stq_0_bits_uop_inst},
     {stq_0_bits_uop_inst},
     {stq_0_bits_uop_inst},
     {stq_0_bits_uop_inst},
     {stq_0_bits_uop_inst},
     {stq_23_bits_uop_inst},
     {stq_22_bits_uop_inst},
     {stq_21_bits_uop_inst},
     {stq_20_bits_uop_inst},
     {stq_19_bits_uop_inst},
     {stq_18_bits_uop_inst},
     {stq_17_bits_uop_inst},
     {stq_16_bits_uop_inst},
     {stq_15_bits_uop_inst},
     {stq_14_bits_uop_inst},
     {stq_13_bits_uop_inst},
     {stq_12_bits_uop_inst},
     {stq_11_bits_uop_inst},
     {stq_10_bits_uop_inst},
     {stq_9_bits_uop_inst},
     {stq_8_bits_uop_inst},
     {stq_7_bits_uop_inst},
     {stq_6_bits_uop_inst},
     {stq_5_bits_uop_inst},
     {stq_4_bits_uop_inst},
     {stq_3_bits_uop_inst},
     {stq_2_bits_uop_inst},
     {stq_1_bits_uop_inst},
     {stq_0_bits_uop_inst}};	// lsu.scala:211:16, :224:42
  wire [31:0][31:0] _GEN_6 =
    {{stq_0_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst},
     {stq_23_bits_uop_debug_inst},
     {stq_22_bits_uop_debug_inst},
     {stq_21_bits_uop_debug_inst},
     {stq_20_bits_uop_debug_inst},
     {stq_19_bits_uop_debug_inst},
     {stq_18_bits_uop_debug_inst},
     {stq_17_bits_uop_debug_inst},
     {stq_16_bits_uop_debug_inst},
     {stq_15_bits_uop_debug_inst},
     {stq_14_bits_uop_debug_inst},
     {stq_13_bits_uop_debug_inst},
     {stq_12_bits_uop_debug_inst},
     {stq_11_bits_uop_debug_inst},
     {stq_10_bits_uop_debug_inst},
     {stq_9_bits_uop_debug_inst},
     {stq_8_bits_uop_debug_inst},
     {stq_7_bits_uop_debug_inst},
     {stq_6_bits_uop_debug_inst},
     {stq_5_bits_uop_debug_inst},
     {stq_4_bits_uop_debug_inst},
     {stq_3_bits_uop_debug_inst},
     {stq_2_bits_uop_debug_inst},
     {stq_1_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_7 =
    {{stq_0_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc},
     {stq_23_bits_uop_is_rvc},
     {stq_22_bits_uop_is_rvc},
     {stq_21_bits_uop_is_rvc},
     {stq_20_bits_uop_is_rvc},
     {stq_19_bits_uop_is_rvc},
     {stq_18_bits_uop_is_rvc},
     {stq_17_bits_uop_is_rvc},
     {stq_16_bits_uop_is_rvc},
     {stq_15_bits_uop_is_rvc},
     {stq_14_bits_uop_is_rvc},
     {stq_13_bits_uop_is_rvc},
     {stq_12_bits_uop_is_rvc},
     {stq_11_bits_uop_is_rvc},
     {stq_10_bits_uop_is_rvc},
     {stq_9_bits_uop_is_rvc},
     {stq_8_bits_uop_is_rvc},
     {stq_7_bits_uop_is_rvc},
     {stq_6_bits_uop_is_rvc},
     {stq_5_bits_uop_is_rvc},
     {stq_4_bits_uop_is_rvc},
     {stq_3_bits_uop_is_rvc},
     {stq_2_bits_uop_is_rvc},
     {stq_1_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc}};	// lsu.scala:211:16, :224:42
  wire [31:0][39:0] _GEN_8 =
    {{stq_0_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc},
     {stq_23_bits_uop_debug_pc},
     {stq_22_bits_uop_debug_pc},
     {stq_21_bits_uop_debug_pc},
     {stq_20_bits_uop_debug_pc},
     {stq_19_bits_uop_debug_pc},
     {stq_18_bits_uop_debug_pc},
     {stq_17_bits_uop_debug_pc},
     {stq_16_bits_uop_debug_pc},
     {stq_15_bits_uop_debug_pc},
     {stq_14_bits_uop_debug_pc},
     {stq_13_bits_uop_debug_pc},
     {stq_12_bits_uop_debug_pc},
     {stq_11_bits_uop_debug_pc},
     {stq_10_bits_uop_debug_pc},
     {stq_9_bits_uop_debug_pc},
     {stq_8_bits_uop_debug_pc},
     {stq_7_bits_uop_debug_pc},
     {stq_6_bits_uop_debug_pc},
     {stq_5_bits_uop_debug_pc},
     {stq_4_bits_uop_debug_pc},
     {stq_3_bits_uop_debug_pc},
     {stq_2_bits_uop_debug_pc},
     {stq_1_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc}};	// lsu.scala:211:16, :224:42
  wire [31:0][2:0]  _GEN_9 =
    {{stq_0_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type},
     {stq_23_bits_uop_iq_type},
     {stq_22_bits_uop_iq_type},
     {stq_21_bits_uop_iq_type},
     {stq_20_bits_uop_iq_type},
     {stq_19_bits_uop_iq_type},
     {stq_18_bits_uop_iq_type},
     {stq_17_bits_uop_iq_type},
     {stq_16_bits_uop_iq_type},
     {stq_15_bits_uop_iq_type},
     {stq_14_bits_uop_iq_type},
     {stq_13_bits_uop_iq_type},
     {stq_12_bits_uop_iq_type},
     {stq_11_bits_uop_iq_type},
     {stq_10_bits_uop_iq_type},
     {stq_9_bits_uop_iq_type},
     {stq_8_bits_uop_iq_type},
     {stq_7_bits_uop_iq_type},
     {stq_6_bits_uop_iq_type},
     {stq_5_bits_uop_iq_type},
     {stq_4_bits_uop_iq_type},
     {stq_3_bits_uop_iq_type},
     {stq_2_bits_uop_iq_type},
     {stq_1_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type}};	// lsu.scala:211:16, :224:42
  wire [31:0][9:0]  _GEN_10 =
    {{stq_0_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code},
     {stq_23_bits_uop_fu_code},
     {stq_22_bits_uop_fu_code},
     {stq_21_bits_uop_fu_code},
     {stq_20_bits_uop_fu_code},
     {stq_19_bits_uop_fu_code},
     {stq_18_bits_uop_fu_code},
     {stq_17_bits_uop_fu_code},
     {stq_16_bits_uop_fu_code},
     {stq_15_bits_uop_fu_code},
     {stq_14_bits_uop_fu_code},
     {stq_13_bits_uop_fu_code},
     {stq_12_bits_uop_fu_code},
     {stq_11_bits_uop_fu_code},
     {stq_10_bits_uop_fu_code},
     {stq_9_bits_uop_fu_code},
     {stq_8_bits_uop_fu_code},
     {stq_7_bits_uop_fu_code},
     {stq_6_bits_uop_fu_code},
     {stq_5_bits_uop_fu_code},
     {stq_4_bits_uop_fu_code},
     {stq_3_bits_uop_fu_code},
     {stq_2_bits_uop_fu_code},
     {stq_1_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code}};	// lsu.scala:211:16, :224:42
  wire [31:0][3:0]  _GEN_11 =
    {{stq_0_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type},
     {stq_23_bits_uop_ctrl_br_type},
     {stq_22_bits_uop_ctrl_br_type},
     {stq_21_bits_uop_ctrl_br_type},
     {stq_20_bits_uop_ctrl_br_type},
     {stq_19_bits_uop_ctrl_br_type},
     {stq_18_bits_uop_ctrl_br_type},
     {stq_17_bits_uop_ctrl_br_type},
     {stq_16_bits_uop_ctrl_br_type},
     {stq_15_bits_uop_ctrl_br_type},
     {stq_14_bits_uop_ctrl_br_type},
     {stq_13_bits_uop_ctrl_br_type},
     {stq_12_bits_uop_ctrl_br_type},
     {stq_11_bits_uop_ctrl_br_type},
     {stq_10_bits_uop_ctrl_br_type},
     {stq_9_bits_uop_ctrl_br_type},
     {stq_8_bits_uop_ctrl_br_type},
     {stq_7_bits_uop_ctrl_br_type},
     {stq_6_bits_uop_ctrl_br_type},
     {stq_5_bits_uop_ctrl_br_type},
     {stq_4_bits_uop_ctrl_br_type},
     {stq_3_bits_uop_ctrl_br_type},
     {stq_2_bits_uop_ctrl_br_type},
     {stq_1_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_12 =
    {{stq_0_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel},
     {stq_23_bits_uop_ctrl_op1_sel},
     {stq_22_bits_uop_ctrl_op1_sel},
     {stq_21_bits_uop_ctrl_op1_sel},
     {stq_20_bits_uop_ctrl_op1_sel},
     {stq_19_bits_uop_ctrl_op1_sel},
     {stq_18_bits_uop_ctrl_op1_sel},
     {stq_17_bits_uop_ctrl_op1_sel},
     {stq_16_bits_uop_ctrl_op1_sel},
     {stq_15_bits_uop_ctrl_op1_sel},
     {stq_14_bits_uop_ctrl_op1_sel},
     {stq_13_bits_uop_ctrl_op1_sel},
     {stq_12_bits_uop_ctrl_op1_sel},
     {stq_11_bits_uop_ctrl_op1_sel},
     {stq_10_bits_uop_ctrl_op1_sel},
     {stq_9_bits_uop_ctrl_op1_sel},
     {stq_8_bits_uop_ctrl_op1_sel},
     {stq_7_bits_uop_ctrl_op1_sel},
     {stq_6_bits_uop_ctrl_op1_sel},
     {stq_5_bits_uop_ctrl_op1_sel},
     {stq_4_bits_uop_ctrl_op1_sel},
     {stq_3_bits_uop_ctrl_op1_sel},
     {stq_2_bits_uop_ctrl_op1_sel},
     {stq_1_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel}};	// lsu.scala:211:16, :224:42
  wire [31:0][2:0]  _GEN_13 =
    {{stq_0_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel},
     {stq_23_bits_uop_ctrl_op2_sel},
     {stq_22_bits_uop_ctrl_op2_sel},
     {stq_21_bits_uop_ctrl_op2_sel},
     {stq_20_bits_uop_ctrl_op2_sel},
     {stq_19_bits_uop_ctrl_op2_sel},
     {stq_18_bits_uop_ctrl_op2_sel},
     {stq_17_bits_uop_ctrl_op2_sel},
     {stq_16_bits_uop_ctrl_op2_sel},
     {stq_15_bits_uop_ctrl_op2_sel},
     {stq_14_bits_uop_ctrl_op2_sel},
     {stq_13_bits_uop_ctrl_op2_sel},
     {stq_12_bits_uop_ctrl_op2_sel},
     {stq_11_bits_uop_ctrl_op2_sel},
     {stq_10_bits_uop_ctrl_op2_sel},
     {stq_9_bits_uop_ctrl_op2_sel},
     {stq_8_bits_uop_ctrl_op2_sel},
     {stq_7_bits_uop_ctrl_op2_sel},
     {stq_6_bits_uop_ctrl_op2_sel},
     {stq_5_bits_uop_ctrl_op2_sel},
     {stq_4_bits_uop_ctrl_op2_sel},
     {stq_3_bits_uop_ctrl_op2_sel},
     {stq_2_bits_uop_ctrl_op2_sel},
     {stq_1_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel}};	// lsu.scala:211:16, :224:42
  wire [31:0][2:0]  _GEN_14 =
    {{stq_0_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel},
     {stq_23_bits_uop_ctrl_imm_sel},
     {stq_22_bits_uop_ctrl_imm_sel},
     {stq_21_bits_uop_ctrl_imm_sel},
     {stq_20_bits_uop_ctrl_imm_sel},
     {stq_19_bits_uop_ctrl_imm_sel},
     {stq_18_bits_uop_ctrl_imm_sel},
     {stq_17_bits_uop_ctrl_imm_sel},
     {stq_16_bits_uop_ctrl_imm_sel},
     {stq_15_bits_uop_ctrl_imm_sel},
     {stq_14_bits_uop_ctrl_imm_sel},
     {stq_13_bits_uop_ctrl_imm_sel},
     {stq_12_bits_uop_ctrl_imm_sel},
     {stq_11_bits_uop_ctrl_imm_sel},
     {stq_10_bits_uop_ctrl_imm_sel},
     {stq_9_bits_uop_ctrl_imm_sel},
     {stq_8_bits_uop_ctrl_imm_sel},
     {stq_7_bits_uop_ctrl_imm_sel},
     {stq_6_bits_uop_ctrl_imm_sel},
     {stq_5_bits_uop_ctrl_imm_sel},
     {stq_4_bits_uop_ctrl_imm_sel},
     {stq_3_bits_uop_ctrl_imm_sel},
     {stq_2_bits_uop_ctrl_imm_sel},
     {stq_1_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel}};	// lsu.scala:211:16, :224:42
  wire [31:0][3:0]  _GEN_15 =
    {{stq_0_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn},
     {stq_23_bits_uop_ctrl_op_fcn},
     {stq_22_bits_uop_ctrl_op_fcn},
     {stq_21_bits_uop_ctrl_op_fcn},
     {stq_20_bits_uop_ctrl_op_fcn},
     {stq_19_bits_uop_ctrl_op_fcn},
     {stq_18_bits_uop_ctrl_op_fcn},
     {stq_17_bits_uop_ctrl_op_fcn},
     {stq_16_bits_uop_ctrl_op_fcn},
     {stq_15_bits_uop_ctrl_op_fcn},
     {stq_14_bits_uop_ctrl_op_fcn},
     {stq_13_bits_uop_ctrl_op_fcn},
     {stq_12_bits_uop_ctrl_op_fcn},
     {stq_11_bits_uop_ctrl_op_fcn},
     {stq_10_bits_uop_ctrl_op_fcn},
     {stq_9_bits_uop_ctrl_op_fcn},
     {stq_8_bits_uop_ctrl_op_fcn},
     {stq_7_bits_uop_ctrl_op_fcn},
     {stq_6_bits_uop_ctrl_op_fcn},
     {stq_5_bits_uop_ctrl_op_fcn},
     {stq_4_bits_uop_ctrl_op_fcn},
     {stq_3_bits_uop_ctrl_op_fcn},
     {stq_2_bits_uop_ctrl_op_fcn},
     {stq_1_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_16 =
    {{stq_0_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw},
     {stq_23_bits_uop_ctrl_fcn_dw},
     {stq_22_bits_uop_ctrl_fcn_dw},
     {stq_21_bits_uop_ctrl_fcn_dw},
     {stq_20_bits_uop_ctrl_fcn_dw},
     {stq_19_bits_uop_ctrl_fcn_dw},
     {stq_18_bits_uop_ctrl_fcn_dw},
     {stq_17_bits_uop_ctrl_fcn_dw},
     {stq_16_bits_uop_ctrl_fcn_dw},
     {stq_15_bits_uop_ctrl_fcn_dw},
     {stq_14_bits_uop_ctrl_fcn_dw},
     {stq_13_bits_uop_ctrl_fcn_dw},
     {stq_12_bits_uop_ctrl_fcn_dw},
     {stq_11_bits_uop_ctrl_fcn_dw},
     {stq_10_bits_uop_ctrl_fcn_dw},
     {stq_9_bits_uop_ctrl_fcn_dw},
     {stq_8_bits_uop_ctrl_fcn_dw},
     {stq_7_bits_uop_ctrl_fcn_dw},
     {stq_6_bits_uop_ctrl_fcn_dw},
     {stq_5_bits_uop_ctrl_fcn_dw},
     {stq_4_bits_uop_ctrl_fcn_dw},
     {stq_3_bits_uop_ctrl_fcn_dw},
     {stq_2_bits_uop_ctrl_fcn_dw},
     {stq_1_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw}};	// lsu.scala:211:16, :224:42
  wire [31:0][2:0]  _GEN_17 =
    {{stq_0_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd},
     {stq_23_bits_uop_ctrl_csr_cmd},
     {stq_22_bits_uop_ctrl_csr_cmd},
     {stq_21_bits_uop_ctrl_csr_cmd},
     {stq_20_bits_uop_ctrl_csr_cmd},
     {stq_19_bits_uop_ctrl_csr_cmd},
     {stq_18_bits_uop_ctrl_csr_cmd},
     {stq_17_bits_uop_ctrl_csr_cmd},
     {stq_16_bits_uop_ctrl_csr_cmd},
     {stq_15_bits_uop_ctrl_csr_cmd},
     {stq_14_bits_uop_ctrl_csr_cmd},
     {stq_13_bits_uop_ctrl_csr_cmd},
     {stq_12_bits_uop_ctrl_csr_cmd},
     {stq_11_bits_uop_ctrl_csr_cmd},
     {stq_10_bits_uop_ctrl_csr_cmd},
     {stq_9_bits_uop_ctrl_csr_cmd},
     {stq_8_bits_uop_ctrl_csr_cmd},
     {stq_7_bits_uop_ctrl_csr_cmd},
     {stq_6_bits_uop_ctrl_csr_cmd},
     {stq_5_bits_uop_ctrl_csr_cmd},
     {stq_4_bits_uop_ctrl_csr_cmd},
     {stq_3_bits_uop_ctrl_csr_cmd},
     {stq_2_bits_uop_ctrl_csr_cmd},
     {stq_1_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_18 =
    {{stq_0_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load},
     {stq_23_bits_uop_ctrl_is_load},
     {stq_22_bits_uop_ctrl_is_load},
     {stq_21_bits_uop_ctrl_is_load},
     {stq_20_bits_uop_ctrl_is_load},
     {stq_19_bits_uop_ctrl_is_load},
     {stq_18_bits_uop_ctrl_is_load},
     {stq_17_bits_uop_ctrl_is_load},
     {stq_16_bits_uop_ctrl_is_load},
     {stq_15_bits_uop_ctrl_is_load},
     {stq_14_bits_uop_ctrl_is_load},
     {stq_13_bits_uop_ctrl_is_load},
     {stq_12_bits_uop_ctrl_is_load},
     {stq_11_bits_uop_ctrl_is_load},
     {stq_10_bits_uop_ctrl_is_load},
     {stq_9_bits_uop_ctrl_is_load},
     {stq_8_bits_uop_ctrl_is_load},
     {stq_7_bits_uop_ctrl_is_load},
     {stq_6_bits_uop_ctrl_is_load},
     {stq_5_bits_uop_ctrl_is_load},
     {stq_4_bits_uop_ctrl_is_load},
     {stq_3_bits_uop_ctrl_is_load},
     {stq_2_bits_uop_ctrl_is_load},
     {stq_1_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_19 =
    {{stq_0_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta},
     {stq_23_bits_uop_ctrl_is_sta},
     {stq_22_bits_uop_ctrl_is_sta},
     {stq_21_bits_uop_ctrl_is_sta},
     {stq_20_bits_uop_ctrl_is_sta},
     {stq_19_bits_uop_ctrl_is_sta},
     {stq_18_bits_uop_ctrl_is_sta},
     {stq_17_bits_uop_ctrl_is_sta},
     {stq_16_bits_uop_ctrl_is_sta},
     {stq_15_bits_uop_ctrl_is_sta},
     {stq_14_bits_uop_ctrl_is_sta},
     {stq_13_bits_uop_ctrl_is_sta},
     {stq_12_bits_uop_ctrl_is_sta},
     {stq_11_bits_uop_ctrl_is_sta},
     {stq_10_bits_uop_ctrl_is_sta},
     {stq_9_bits_uop_ctrl_is_sta},
     {stq_8_bits_uop_ctrl_is_sta},
     {stq_7_bits_uop_ctrl_is_sta},
     {stq_6_bits_uop_ctrl_is_sta},
     {stq_5_bits_uop_ctrl_is_sta},
     {stq_4_bits_uop_ctrl_is_sta},
     {stq_3_bits_uop_ctrl_is_sta},
     {stq_2_bits_uop_ctrl_is_sta},
     {stq_1_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_20 =
    {{stq_0_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std},
     {stq_23_bits_uop_ctrl_is_std},
     {stq_22_bits_uop_ctrl_is_std},
     {stq_21_bits_uop_ctrl_is_std},
     {stq_20_bits_uop_ctrl_is_std},
     {stq_19_bits_uop_ctrl_is_std},
     {stq_18_bits_uop_ctrl_is_std},
     {stq_17_bits_uop_ctrl_is_std},
     {stq_16_bits_uop_ctrl_is_std},
     {stq_15_bits_uop_ctrl_is_std},
     {stq_14_bits_uop_ctrl_is_std},
     {stq_13_bits_uop_ctrl_is_std},
     {stq_12_bits_uop_ctrl_is_std},
     {stq_11_bits_uop_ctrl_is_std},
     {stq_10_bits_uop_ctrl_is_std},
     {stq_9_bits_uop_ctrl_is_std},
     {stq_8_bits_uop_ctrl_is_std},
     {stq_7_bits_uop_ctrl_is_std},
     {stq_6_bits_uop_ctrl_is_std},
     {stq_5_bits_uop_ctrl_is_std},
     {stq_4_bits_uop_ctrl_is_std},
     {stq_3_bits_uop_ctrl_is_std},
     {stq_2_bits_uop_ctrl_is_std},
     {stq_1_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_21 =
    {{stq_0_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state},
     {stq_23_bits_uop_iw_state},
     {stq_22_bits_uop_iw_state},
     {stq_21_bits_uop_iw_state},
     {stq_20_bits_uop_iw_state},
     {stq_19_bits_uop_iw_state},
     {stq_18_bits_uop_iw_state},
     {stq_17_bits_uop_iw_state},
     {stq_16_bits_uop_iw_state},
     {stq_15_bits_uop_iw_state},
     {stq_14_bits_uop_iw_state},
     {stq_13_bits_uop_iw_state},
     {stq_12_bits_uop_iw_state},
     {stq_11_bits_uop_iw_state},
     {stq_10_bits_uop_iw_state},
     {stq_9_bits_uop_iw_state},
     {stq_8_bits_uop_iw_state},
     {stq_7_bits_uop_iw_state},
     {stq_6_bits_uop_iw_state},
     {stq_5_bits_uop_iw_state},
     {stq_4_bits_uop_iw_state},
     {stq_3_bits_uop_iw_state},
     {stq_2_bits_uop_iw_state},
     {stq_1_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_22 =
    {{stq_0_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned},
     {stq_23_bits_uop_iw_p1_poisoned},
     {stq_22_bits_uop_iw_p1_poisoned},
     {stq_21_bits_uop_iw_p1_poisoned},
     {stq_20_bits_uop_iw_p1_poisoned},
     {stq_19_bits_uop_iw_p1_poisoned},
     {stq_18_bits_uop_iw_p1_poisoned},
     {stq_17_bits_uop_iw_p1_poisoned},
     {stq_16_bits_uop_iw_p1_poisoned},
     {stq_15_bits_uop_iw_p1_poisoned},
     {stq_14_bits_uop_iw_p1_poisoned},
     {stq_13_bits_uop_iw_p1_poisoned},
     {stq_12_bits_uop_iw_p1_poisoned},
     {stq_11_bits_uop_iw_p1_poisoned},
     {stq_10_bits_uop_iw_p1_poisoned},
     {stq_9_bits_uop_iw_p1_poisoned},
     {stq_8_bits_uop_iw_p1_poisoned},
     {stq_7_bits_uop_iw_p1_poisoned},
     {stq_6_bits_uop_iw_p1_poisoned},
     {stq_5_bits_uop_iw_p1_poisoned},
     {stq_4_bits_uop_iw_p1_poisoned},
     {stq_3_bits_uop_iw_p1_poisoned},
     {stq_2_bits_uop_iw_p1_poisoned},
     {stq_1_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_23 =
    {{stq_0_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned},
     {stq_23_bits_uop_iw_p2_poisoned},
     {stq_22_bits_uop_iw_p2_poisoned},
     {stq_21_bits_uop_iw_p2_poisoned},
     {stq_20_bits_uop_iw_p2_poisoned},
     {stq_19_bits_uop_iw_p2_poisoned},
     {stq_18_bits_uop_iw_p2_poisoned},
     {stq_17_bits_uop_iw_p2_poisoned},
     {stq_16_bits_uop_iw_p2_poisoned},
     {stq_15_bits_uop_iw_p2_poisoned},
     {stq_14_bits_uop_iw_p2_poisoned},
     {stq_13_bits_uop_iw_p2_poisoned},
     {stq_12_bits_uop_iw_p2_poisoned},
     {stq_11_bits_uop_iw_p2_poisoned},
     {stq_10_bits_uop_iw_p2_poisoned},
     {stq_9_bits_uop_iw_p2_poisoned},
     {stq_8_bits_uop_iw_p2_poisoned},
     {stq_7_bits_uop_iw_p2_poisoned},
     {stq_6_bits_uop_iw_p2_poisoned},
     {stq_5_bits_uop_iw_p2_poisoned},
     {stq_4_bits_uop_iw_p2_poisoned},
     {stq_3_bits_uop_iw_p2_poisoned},
     {stq_2_bits_uop_iw_p2_poisoned},
     {stq_1_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_24 =
    {{stq_0_bits_uop_is_br},
     {stq_0_bits_uop_is_br},
     {stq_0_bits_uop_is_br},
     {stq_0_bits_uop_is_br},
     {stq_0_bits_uop_is_br},
     {stq_0_bits_uop_is_br},
     {stq_0_bits_uop_is_br},
     {stq_0_bits_uop_is_br},
     {stq_23_bits_uop_is_br},
     {stq_22_bits_uop_is_br},
     {stq_21_bits_uop_is_br},
     {stq_20_bits_uop_is_br},
     {stq_19_bits_uop_is_br},
     {stq_18_bits_uop_is_br},
     {stq_17_bits_uop_is_br},
     {stq_16_bits_uop_is_br},
     {stq_15_bits_uop_is_br},
     {stq_14_bits_uop_is_br},
     {stq_13_bits_uop_is_br},
     {stq_12_bits_uop_is_br},
     {stq_11_bits_uop_is_br},
     {stq_10_bits_uop_is_br},
     {stq_9_bits_uop_is_br},
     {stq_8_bits_uop_is_br},
     {stq_7_bits_uop_is_br},
     {stq_6_bits_uop_is_br},
     {stq_5_bits_uop_is_br},
     {stq_4_bits_uop_is_br},
     {stq_3_bits_uop_is_br},
     {stq_2_bits_uop_is_br},
     {stq_1_bits_uop_is_br},
     {stq_0_bits_uop_is_br}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_25 =
    {{stq_0_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr},
     {stq_23_bits_uop_is_jalr},
     {stq_22_bits_uop_is_jalr},
     {stq_21_bits_uop_is_jalr},
     {stq_20_bits_uop_is_jalr},
     {stq_19_bits_uop_is_jalr},
     {stq_18_bits_uop_is_jalr},
     {stq_17_bits_uop_is_jalr},
     {stq_16_bits_uop_is_jalr},
     {stq_15_bits_uop_is_jalr},
     {stq_14_bits_uop_is_jalr},
     {stq_13_bits_uop_is_jalr},
     {stq_12_bits_uop_is_jalr},
     {stq_11_bits_uop_is_jalr},
     {stq_10_bits_uop_is_jalr},
     {stq_9_bits_uop_is_jalr},
     {stq_8_bits_uop_is_jalr},
     {stq_7_bits_uop_is_jalr},
     {stq_6_bits_uop_is_jalr},
     {stq_5_bits_uop_is_jalr},
     {stq_4_bits_uop_is_jalr},
     {stq_3_bits_uop_is_jalr},
     {stq_2_bits_uop_is_jalr},
     {stq_1_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_26 =
    {{stq_0_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal},
     {stq_23_bits_uop_is_jal},
     {stq_22_bits_uop_is_jal},
     {stq_21_bits_uop_is_jal},
     {stq_20_bits_uop_is_jal},
     {stq_19_bits_uop_is_jal},
     {stq_18_bits_uop_is_jal},
     {stq_17_bits_uop_is_jal},
     {stq_16_bits_uop_is_jal},
     {stq_15_bits_uop_is_jal},
     {stq_14_bits_uop_is_jal},
     {stq_13_bits_uop_is_jal},
     {stq_12_bits_uop_is_jal},
     {stq_11_bits_uop_is_jal},
     {stq_10_bits_uop_is_jal},
     {stq_9_bits_uop_is_jal},
     {stq_8_bits_uop_is_jal},
     {stq_7_bits_uop_is_jal},
     {stq_6_bits_uop_is_jal},
     {stq_5_bits_uop_is_jal},
     {stq_4_bits_uop_is_jal},
     {stq_3_bits_uop_is_jal},
     {stq_2_bits_uop_is_jal},
     {stq_1_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_27 =
    {{stq_0_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb},
     {stq_23_bits_uop_is_sfb},
     {stq_22_bits_uop_is_sfb},
     {stq_21_bits_uop_is_sfb},
     {stq_20_bits_uop_is_sfb},
     {stq_19_bits_uop_is_sfb},
     {stq_18_bits_uop_is_sfb},
     {stq_17_bits_uop_is_sfb},
     {stq_16_bits_uop_is_sfb},
     {stq_15_bits_uop_is_sfb},
     {stq_14_bits_uop_is_sfb},
     {stq_13_bits_uop_is_sfb},
     {stq_12_bits_uop_is_sfb},
     {stq_11_bits_uop_is_sfb},
     {stq_10_bits_uop_is_sfb},
     {stq_9_bits_uop_is_sfb},
     {stq_8_bits_uop_is_sfb},
     {stq_7_bits_uop_is_sfb},
     {stq_6_bits_uop_is_sfb},
     {stq_5_bits_uop_is_sfb},
     {stq_4_bits_uop_is_sfb},
     {stq_3_bits_uop_is_sfb},
     {stq_2_bits_uop_is_sfb},
     {stq_1_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb}};	// lsu.scala:211:16, :224:42
  wire [31:0][15:0] _GEN_28 =
    {{stq_0_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask},
     {stq_23_bits_uop_br_mask},
     {stq_22_bits_uop_br_mask},
     {stq_21_bits_uop_br_mask},
     {stq_20_bits_uop_br_mask},
     {stq_19_bits_uop_br_mask},
     {stq_18_bits_uop_br_mask},
     {stq_17_bits_uop_br_mask},
     {stq_16_bits_uop_br_mask},
     {stq_15_bits_uop_br_mask},
     {stq_14_bits_uop_br_mask},
     {stq_13_bits_uop_br_mask},
     {stq_12_bits_uop_br_mask},
     {stq_11_bits_uop_br_mask},
     {stq_10_bits_uop_br_mask},
     {stq_9_bits_uop_br_mask},
     {stq_8_bits_uop_br_mask},
     {stq_7_bits_uop_br_mask},
     {stq_6_bits_uop_br_mask},
     {stq_5_bits_uop_br_mask},
     {stq_4_bits_uop_br_mask},
     {stq_3_bits_uop_br_mask},
     {stq_2_bits_uop_br_mask},
     {stq_1_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask}};	// lsu.scala:211:16, :224:42
  wire [31:0][3:0]  _GEN_29 =
    {{stq_0_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag},
     {stq_23_bits_uop_br_tag},
     {stq_22_bits_uop_br_tag},
     {stq_21_bits_uop_br_tag},
     {stq_20_bits_uop_br_tag},
     {stq_19_bits_uop_br_tag},
     {stq_18_bits_uop_br_tag},
     {stq_17_bits_uop_br_tag},
     {stq_16_bits_uop_br_tag},
     {stq_15_bits_uop_br_tag},
     {stq_14_bits_uop_br_tag},
     {stq_13_bits_uop_br_tag},
     {stq_12_bits_uop_br_tag},
     {stq_11_bits_uop_br_tag},
     {stq_10_bits_uop_br_tag},
     {stq_9_bits_uop_br_tag},
     {stq_8_bits_uop_br_tag},
     {stq_7_bits_uop_br_tag},
     {stq_6_bits_uop_br_tag},
     {stq_5_bits_uop_br_tag},
     {stq_4_bits_uop_br_tag},
     {stq_3_bits_uop_br_tag},
     {stq_2_bits_uop_br_tag},
     {stq_1_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag}};	// lsu.scala:211:16, :224:42
  wire [31:0][4:0]  _GEN_30 =
    {{stq_0_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx},
     {stq_23_bits_uop_ftq_idx},
     {stq_22_bits_uop_ftq_idx},
     {stq_21_bits_uop_ftq_idx},
     {stq_20_bits_uop_ftq_idx},
     {stq_19_bits_uop_ftq_idx},
     {stq_18_bits_uop_ftq_idx},
     {stq_17_bits_uop_ftq_idx},
     {stq_16_bits_uop_ftq_idx},
     {stq_15_bits_uop_ftq_idx},
     {stq_14_bits_uop_ftq_idx},
     {stq_13_bits_uop_ftq_idx},
     {stq_12_bits_uop_ftq_idx},
     {stq_11_bits_uop_ftq_idx},
     {stq_10_bits_uop_ftq_idx},
     {stq_9_bits_uop_ftq_idx},
     {stq_8_bits_uop_ftq_idx},
     {stq_7_bits_uop_ftq_idx},
     {stq_6_bits_uop_ftq_idx},
     {stq_5_bits_uop_ftq_idx},
     {stq_4_bits_uop_ftq_idx},
     {stq_3_bits_uop_ftq_idx},
     {stq_2_bits_uop_ftq_idx},
     {stq_1_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_31 =
    {{stq_0_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst},
     {stq_23_bits_uop_edge_inst},
     {stq_22_bits_uop_edge_inst},
     {stq_21_bits_uop_edge_inst},
     {stq_20_bits_uop_edge_inst},
     {stq_19_bits_uop_edge_inst},
     {stq_18_bits_uop_edge_inst},
     {stq_17_bits_uop_edge_inst},
     {stq_16_bits_uop_edge_inst},
     {stq_15_bits_uop_edge_inst},
     {stq_14_bits_uop_edge_inst},
     {stq_13_bits_uop_edge_inst},
     {stq_12_bits_uop_edge_inst},
     {stq_11_bits_uop_edge_inst},
     {stq_10_bits_uop_edge_inst},
     {stq_9_bits_uop_edge_inst},
     {stq_8_bits_uop_edge_inst},
     {stq_7_bits_uop_edge_inst},
     {stq_6_bits_uop_edge_inst},
     {stq_5_bits_uop_edge_inst},
     {stq_4_bits_uop_edge_inst},
     {stq_3_bits_uop_edge_inst},
     {stq_2_bits_uop_edge_inst},
     {stq_1_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst}};	// lsu.scala:211:16, :224:42
  wire [31:0][5:0]  _GEN_32 =
    {{stq_0_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob},
     {stq_23_bits_uop_pc_lob},
     {stq_22_bits_uop_pc_lob},
     {stq_21_bits_uop_pc_lob},
     {stq_20_bits_uop_pc_lob},
     {stq_19_bits_uop_pc_lob},
     {stq_18_bits_uop_pc_lob},
     {stq_17_bits_uop_pc_lob},
     {stq_16_bits_uop_pc_lob},
     {stq_15_bits_uop_pc_lob},
     {stq_14_bits_uop_pc_lob},
     {stq_13_bits_uop_pc_lob},
     {stq_12_bits_uop_pc_lob},
     {stq_11_bits_uop_pc_lob},
     {stq_10_bits_uop_pc_lob},
     {stq_9_bits_uop_pc_lob},
     {stq_8_bits_uop_pc_lob},
     {stq_7_bits_uop_pc_lob},
     {stq_6_bits_uop_pc_lob},
     {stq_5_bits_uop_pc_lob},
     {stq_4_bits_uop_pc_lob},
     {stq_3_bits_uop_pc_lob},
     {stq_2_bits_uop_pc_lob},
     {stq_1_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_33 =
    {{stq_0_bits_uop_taken},
     {stq_0_bits_uop_taken},
     {stq_0_bits_uop_taken},
     {stq_0_bits_uop_taken},
     {stq_0_bits_uop_taken},
     {stq_0_bits_uop_taken},
     {stq_0_bits_uop_taken},
     {stq_0_bits_uop_taken},
     {stq_23_bits_uop_taken},
     {stq_22_bits_uop_taken},
     {stq_21_bits_uop_taken},
     {stq_20_bits_uop_taken},
     {stq_19_bits_uop_taken},
     {stq_18_bits_uop_taken},
     {stq_17_bits_uop_taken},
     {stq_16_bits_uop_taken},
     {stq_15_bits_uop_taken},
     {stq_14_bits_uop_taken},
     {stq_13_bits_uop_taken},
     {stq_12_bits_uop_taken},
     {stq_11_bits_uop_taken},
     {stq_10_bits_uop_taken},
     {stq_9_bits_uop_taken},
     {stq_8_bits_uop_taken},
     {stq_7_bits_uop_taken},
     {stq_6_bits_uop_taken},
     {stq_5_bits_uop_taken},
     {stq_4_bits_uop_taken},
     {stq_3_bits_uop_taken},
     {stq_2_bits_uop_taken},
     {stq_1_bits_uop_taken},
     {stq_0_bits_uop_taken}};	// lsu.scala:211:16, :224:42
  wire [31:0][19:0] _GEN_34 =
    {{stq_0_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed},
     {stq_23_bits_uop_imm_packed},
     {stq_22_bits_uop_imm_packed},
     {stq_21_bits_uop_imm_packed},
     {stq_20_bits_uop_imm_packed},
     {stq_19_bits_uop_imm_packed},
     {stq_18_bits_uop_imm_packed},
     {stq_17_bits_uop_imm_packed},
     {stq_16_bits_uop_imm_packed},
     {stq_15_bits_uop_imm_packed},
     {stq_14_bits_uop_imm_packed},
     {stq_13_bits_uop_imm_packed},
     {stq_12_bits_uop_imm_packed},
     {stq_11_bits_uop_imm_packed},
     {stq_10_bits_uop_imm_packed},
     {stq_9_bits_uop_imm_packed},
     {stq_8_bits_uop_imm_packed},
     {stq_7_bits_uop_imm_packed},
     {stq_6_bits_uop_imm_packed},
     {stq_5_bits_uop_imm_packed},
     {stq_4_bits_uop_imm_packed},
     {stq_3_bits_uop_imm_packed},
     {stq_2_bits_uop_imm_packed},
     {stq_1_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed}};	// lsu.scala:211:16, :224:42
  wire [31:0][11:0] _GEN_35 =
    {{stq_0_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr},
     {stq_23_bits_uop_csr_addr},
     {stq_22_bits_uop_csr_addr},
     {stq_21_bits_uop_csr_addr},
     {stq_20_bits_uop_csr_addr},
     {stq_19_bits_uop_csr_addr},
     {stq_18_bits_uop_csr_addr},
     {stq_17_bits_uop_csr_addr},
     {stq_16_bits_uop_csr_addr},
     {stq_15_bits_uop_csr_addr},
     {stq_14_bits_uop_csr_addr},
     {stq_13_bits_uop_csr_addr},
     {stq_12_bits_uop_csr_addr},
     {stq_11_bits_uop_csr_addr},
     {stq_10_bits_uop_csr_addr},
     {stq_9_bits_uop_csr_addr},
     {stq_8_bits_uop_csr_addr},
     {stq_7_bits_uop_csr_addr},
     {stq_6_bits_uop_csr_addr},
     {stq_5_bits_uop_csr_addr},
     {stq_4_bits_uop_csr_addr},
     {stq_3_bits_uop_csr_addr},
     {stq_2_bits_uop_csr_addr},
     {stq_1_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr}};	// lsu.scala:211:16, :224:42
  wire [31:0][6:0]  _GEN_36 =
    {{stq_0_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx},
     {stq_23_bits_uop_rob_idx},
     {stq_22_bits_uop_rob_idx},
     {stq_21_bits_uop_rob_idx},
     {stq_20_bits_uop_rob_idx},
     {stq_19_bits_uop_rob_idx},
     {stq_18_bits_uop_rob_idx},
     {stq_17_bits_uop_rob_idx},
     {stq_16_bits_uop_rob_idx},
     {stq_15_bits_uop_rob_idx},
     {stq_14_bits_uop_rob_idx},
     {stq_13_bits_uop_rob_idx},
     {stq_12_bits_uop_rob_idx},
     {stq_11_bits_uop_rob_idx},
     {stq_10_bits_uop_rob_idx},
     {stq_9_bits_uop_rob_idx},
     {stq_8_bits_uop_rob_idx},
     {stq_7_bits_uop_rob_idx},
     {stq_6_bits_uop_rob_idx},
     {stq_5_bits_uop_rob_idx},
     {stq_4_bits_uop_rob_idx},
     {stq_3_bits_uop_rob_idx},
     {stq_2_bits_uop_rob_idx},
     {stq_1_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx}};	// lsu.scala:211:16, :224:42
  wire [31:0][4:0]  _GEN_37 =
    {{stq_0_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx},
     {stq_23_bits_uop_ldq_idx},
     {stq_22_bits_uop_ldq_idx},
     {stq_21_bits_uop_ldq_idx},
     {stq_20_bits_uop_ldq_idx},
     {stq_19_bits_uop_ldq_idx},
     {stq_18_bits_uop_ldq_idx},
     {stq_17_bits_uop_ldq_idx},
     {stq_16_bits_uop_ldq_idx},
     {stq_15_bits_uop_ldq_idx},
     {stq_14_bits_uop_ldq_idx},
     {stq_13_bits_uop_ldq_idx},
     {stq_12_bits_uop_ldq_idx},
     {stq_11_bits_uop_ldq_idx},
     {stq_10_bits_uop_ldq_idx},
     {stq_9_bits_uop_ldq_idx},
     {stq_8_bits_uop_ldq_idx},
     {stq_7_bits_uop_ldq_idx},
     {stq_6_bits_uop_ldq_idx},
     {stq_5_bits_uop_ldq_idx},
     {stq_4_bits_uop_ldq_idx},
     {stq_3_bits_uop_ldq_idx},
     {stq_2_bits_uop_ldq_idx},
     {stq_1_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx}};	// lsu.scala:211:16, :224:42
  wire [31:0][4:0]  _GEN_38 =
    {{stq_0_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx},
     {stq_23_bits_uop_stq_idx},
     {stq_22_bits_uop_stq_idx},
     {stq_21_bits_uop_stq_idx},
     {stq_20_bits_uop_stq_idx},
     {stq_19_bits_uop_stq_idx},
     {stq_18_bits_uop_stq_idx},
     {stq_17_bits_uop_stq_idx},
     {stq_16_bits_uop_stq_idx},
     {stq_15_bits_uop_stq_idx},
     {stq_14_bits_uop_stq_idx},
     {stq_13_bits_uop_stq_idx},
     {stq_12_bits_uop_stq_idx},
     {stq_11_bits_uop_stq_idx},
     {stq_10_bits_uop_stq_idx},
     {stq_9_bits_uop_stq_idx},
     {stq_8_bits_uop_stq_idx},
     {stq_7_bits_uop_stq_idx},
     {stq_6_bits_uop_stq_idx},
     {stq_5_bits_uop_stq_idx},
     {stq_4_bits_uop_stq_idx},
     {stq_3_bits_uop_stq_idx},
     {stq_2_bits_uop_stq_idx},
     {stq_1_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_39 =
    {{stq_0_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx},
     {stq_23_bits_uop_rxq_idx},
     {stq_22_bits_uop_rxq_idx},
     {stq_21_bits_uop_rxq_idx},
     {stq_20_bits_uop_rxq_idx},
     {stq_19_bits_uop_rxq_idx},
     {stq_18_bits_uop_rxq_idx},
     {stq_17_bits_uop_rxq_idx},
     {stq_16_bits_uop_rxq_idx},
     {stq_15_bits_uop_rxq_idx},
     {stq_14_bits_uop_rxq_idx},
     {stq_13_bits_uop_rxq_idx},
     {stq_12_bits_uop_rxq_idx},
     {stq_11_bits_uop_rxq_idx},
     {stq_10_bits_uop_rxq_idx},
     {stq_9_bits_uop_rxq_idx},
     {stq_8_bits_uop_rxq_idx},
     {stq_7_bits_uop_rxq_idx},
     {stq_6_bits_uop_rxq_idx},
     {stq_5_bits_uop_rxq_idx},
     {stq_4_bits_uop_rxq_idx},
     {stq_3_bits_uop_rxq_idx},
     {stq_2_bits_uop_rxq_idx},
     {stq_1_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx}};	// lsu.scala:211:16, :224:42
  wire [31:0][6:0]  _GEN_40 =
    {{stq_0_bits_uop_pdst},
     {stq_0_bits_uop_pdst},
     {stq_0_bits_uop_pdst},
     {stq_0_bits_uop_pdst},
     {stq_0_bits_uop_pdst},
     {stq_0_bits_uop_pdst},
     {stq_0_bits_uop_pdst},
     {stq_0_bits_uop_pdst},
     {stq_23_bits_uop_pdst},
     {stq_22_bits_uop_pdst},
     {stq_21_bits_uop_pdst},
     {stq_20_bits_uop_pdst},
     {stq_19_bits_uop_pdst},
     {stq_18_bits_uop_pdst},
     {stq_17_bits_uop_pdst},
     {stq_16_bits_uop_pdst},
     {stq_15_bits_uop_pdst},
     {stq_14_bits_uop_pdst},
     {stq_13_bits_uop_pdst},
     {stq_12_bits_uop_pdst},
     {stq_11_bits_uop_pdst},
     {stq_10_bits_uop_pdst},
     {stq_9_bits_uop_pdst},
     {stq_8_bits_uop_pdst},
     {stq_7_bits_uop_pdst},
     {stq_6_bits_uop_pdst},
     {stq_5_bits_uop_pdst},
     {stq_4_bits_uop_pdst},
     {stq_3_bits_uop_pdst},
     {stq_2_bits_uop_pdst},
     {stq_1_bits_uop_pdst},
     {stq_0_bits_uop_pdst}};	// lsu.scala:211:16, :224:42
  wire [31:0][6:0]  _GEN_41 =
    {{stq_0_bits_uop_prs1},
     {stq_0_bits_uop_prs1},
     {stq_0_bits_uop_prs1},
     {stq_0_bits_uop_prs1},
     {stq_0_bits_uop_prs1},
     {stq_0_bits_uop_prs1},
     {stq_0_bits_uop_prs1},
     {stq_0_bits_uop_prs1},
     {stq_23_bits_uop_prs1},
     {stq_22_bits_uop_prs1},
     {stq_21_bits_uop_prs1},
     {stq_20_bits_uop_prs1},
     {stq_19_bits_uop_prs1},
     {stq_18_bits_uop_prs1},
     {stq_17_bits_uop_prs1},
     {stq_16_bits_uop_prs1},
     {stq_15_bits_uop_prs1},
     {stq_14_bits_uop_prs1},
     {stq_13_bits_uop_prs1},
     {stq_12_bits_uop_prs1},
     {stq_11_bits_uop_prs1},
     {stq_10_bits_uop_prs1},
     {stq_9_bits_uop_prs1},
     {stq_8_bits_uop_prs1},
     {stq_7_bits_uop_prs1},
     {stq_6_bits_uop_prs1},
     {stq_5_bits_uop_prs1},
     {stq_4_bits_uop_prs1},
     {stq_3_bits_uop_prs1},
     {stq_2_bits_uop_prs1},
     {stq_1_bits_uop_prs1},
     {stq_0_bits_uop_prs1}};	// lsu.scala:211:16, :224:42
  wire [31:0][6:0]  _GEN_42 =
    {{stq_0_bits_uop_prs2},
     {stq_0_bits_uop_prs2},
     {stq_0_bits_uop_prs2},
     {stq_0_bits_uop_prs2},
     {stq_0_bits_uop_prs2},
     {stq_0_bits_uop_prs2},
     {stq_0_bits_uop_prs2},
     {stq_0_bits_uop_prs2},
     {stq_23_bits_uop_prs2},
     {stq_22_bits_uop_prs2},
     {stq_21_bits_uop_prs2},
     {stq_20_bits_uop_prs2},
     {stq_19_bits_uop_prs2},
     {stq_18_bits_uop_prs2},
     {stq_17_bits_uop_prs2},
     {stq_16_bits_uop_prs2},
     {stq_15_bits_uop_prs2},
     {stq_14_bits_uop_prs2},
     {stq_13_bits_uop_prs2},
     {stq_12_bits_uop_prs2},
     {stq_11_bits_uop_prs2},
     {stq_10_bits_uop_prs2},
     {stq_9_bits_uop_prs2},
     {stq_8_bits_uop_prs2},
     {stq_7_bits_uop_prs2},
     {stq_6_bits_uop_prs2},
     {stq_5_bits_uop_prs2},
     {stq_4_bits_uop_prs2},
     {stq_3_bits_uop_prs2},
     {stq_2_bits_uop_prs2},
     {stq_1_bits_uop_prs2},
     {stq_0_bits_uop_prs2}};	// lsu.scala:211:16, :224:42
  wire [31:0][6:0]  _GEN_43 =
    {{stq_0_bits_uop_prs3},
     {stq_0_bits_uop_prs3},
     {stq_0_bits_uop_prs3},
     {stq_0_bits_uop_prs3},
     {stq_0_bits_uop_prs3},
     {stq_0_bits_uop_prs3},
     {stq_0_bits_uop_prs3},
     {stq_0_bits_uop_prs3},
     {stq_23_bits_uop_prs3},
     {stq_22_bits_uop_prs3},
     {stq_21_bits_uop_prs3},
     {stq_20_bits_uop_prs3},
     {stq_19_bits_uop_prs3},
     {stq_18_bits_uop_prs3},
     {stq_17_bits_uop_prs3},
     {stq_16_bits_uop_prs3},
     {stq_15_bits_uop_prs3},
     {stq_14_bits_uop_prs3},
     {stq_13_bits_uop_prs3},
     {stq_12_bits_uop_prs3},
     {stq_11_bits_uop_prs3},
     {stq_10_bits_uop_prs3},
     {stq_9_bits_uop_prs3},
     {stq_8_bits_uop_prs3},
     {stq_7_bits_uop_prs3},
     {stq_6_bits_uop_prs3},
     {stq_5_bits_uop_prs3},
     {stq_4_bits_uop_prs3},
     {stq_3_bits_uop_prs3},
     {stq_2_bits_uop_prs3},
     {stq_1_bits_uop_prs3},
     {stq_0_bits_uop_prs3}};	// lsu.scala:211:16, :224:42
  wire [31:0][4:0]  _GEN_44 =
    {{stq_0_bits_uop_ppred},
     {stq_0_bits_uop_ppred},
     {stq_0_bits_uop_ppred},
     {stq_0_bits_uop_ppred},
     {stq_0_bits_uop_ppred},
     {stq_0_bits_uop_ppred},
     {stq_0_bits_uop_ppred},
     {stq_0_bits_uop_ppred},
     {stq_23_bits_uop_ppred},
     {stq_22_bits_uop_ppred},
     {stq_21_bits_uop_ppred},
     {stq_20_bits_uop_ppred},
     {stq_19_bits_uop_ppred},
     {stq_18_bits_uop_ppred},
     {stq_17_bits_uop_ppred},
     {stq_16_bits_uop_ppred},
     {stq_15_bits_uop_ppred},
     {stq_14_bits_uop_ppred},
     {stq_13_bits_uop_ppred},
     {stq_12_bits_uop_ppred},
     {stq_11_bits_uop_ppred},
     {stq_10_bits_uop_ppred},
     {stq_9_bits_uop_ppred},
     {stq_8_bits_uop_ppred},
     {stq_7_bits_uop_ppred},
     {stq_6_bits_uop_ppred},
     {stq_5_bits_uop_ppred},
     {stq_4_bits_uop_ppred},
     {stq_3_bits_uop_ppred},
     {stq_2_bits_uop_ppred},
     {stq_1_bits_uop_ppred},
     {stq_0_bits_uop_ppred}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_45 =
    {{stq_0_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy},
     {stq_23_bits_uop_prs1_busy},
     {stq_22_bits_uop_prs1_busy},
     {stq_21_bits_uop_prs1_busy},
     {stq_20_bits_uop_prs1_busy},
     {stq_19_bits_uop_prs1_busy},
     {stq_18_bits_uop_prs1_busy},
     {stq_17_bits_uop_prs1_busy},
     {stq_16_bits_uop_prs1_busy},
     {stq_15_bits_uop_prs1_busy},
     {stq_14_bits_uop_prs1_busy},
     {stq_13_bits_uop_prs1_busy},
     {stq_12_bits_uop_prs1_busy},
     {stq_11_bits_uop_prs1_busy},
     {stq_10_bits_uop_prs1_busy},
     {stq_9_bits_uop_prs1_busy},
     {stq_8_bits_uop_prs1_busy},
     {stq_7_bits_uop_prs1_busy},
     {stq_6_bits_uop_prs1_busy},
     {stq_5_bits_uop_prs1_busy},
     {stq_4_bits_uop_prs1_busy},
     {stq_3_bits_uop_prs1_busy},
     {stq_2_bits_uop_prs1_busy},
     {stq_1_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_46 =
    {{stq_0_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy},
     {stq_23_bits_uop_prs2_busy},
     {stq_22_bits_uop_prs2_busy},
     {stq_21_bits_uop_prs2_busy},
     {stq_20_bits_uop_prs2_busy},
     {stq_19_bits_uop_prs2_busy},
     {stq_18_bits_uop_prs2_busy},
     {stq_17_bits_uop_prs2_busy},
     {stq_16_bits_uop_prs2_busy},
     {stq_15_bits_uop_prs2_busy},
     {stq_14_bits_uop_prs2_busy},
     {stq_13_bits_uop_prs2_busy},
     {stq_12_bits_uop_prs2_busy},
     {stq_11_bits_uop_prs2_busy},
     {stq_10_bits_uop_prs2_busy},
     {stq_9_bits_uop_prs2_busy},
     {stq_8_bits_uop_prs2_busy},
     {stq_7_bits_uop_prs2_busy},
     {stq_6_bits_uop_prs2_busy},
     {stq_5_bits_uop_prs2_busy},
     {stq_4_bits_uop_prs2_busy},
     {stq_3_bits_uop_prs2_busy},
     {stq_2_bits_uop_prs2_busy},
     {stq_1_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_47 =
    {{stq_0_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy},
     {stq_23_bits_uop_prs3_busy},
     {stq_22_bits_uop_prs3_busy},
     {stq_21_bits_uop_prs3_busy},
     {stq_20_bits_uop_prs3_busy},
     {stq_19_bits_uop_prs3_busy},
     {stq_18_bits_uop_prs3_busy},
     {stq_17_bits_uop_prs3_busy},
     {stq_16_bits_uop_prs3_busy},
     {stq_15_bits_uop_prs3_busy},
     {stq_14_bits_uop_prs3_busy},
     {stq_13_bits_uop_prs3_busy},
     {stq_12_bits_uop_prs3_busy},
     {stq_11_bits_uop_prs3_busy},
     {stq_10_bits_uop_prs3_busy},
     {stq_9_bits_uop_prs3_busy},
     {stq_8_bits_uop_prs3_busy},
     {stq_7_bits_uop_prs3_busy},
     {stq_6_bits_uop_prs3_busy},
     {stq_5_bits_uop_prs3_busy},
     {stq_4_bits_uop_prs3_busy},
     {stq_3_bits_uop_prs3_busy},
     {stq_2_bits_uop_prs3_busy},
     {stq_1_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_48 =
    {{stq_0_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy},
     {stq_23_bits_uop_ppred_busy},
     {stq_22_bits_uop_ppred_busy},
     {stq_21_bits_uop_ppred_busy},
     {stq_20_bits_uop_ppred_busy},
     {stq_19_bits_uop_ppred_busy},
     {stq_18_bits_uop_ppred_busy},
     {stq_17_bits_uop_ppred_busy},
     {stq_16_bits_uop_ppred_busy},
     {stq_15_bits_uop_ppred_busy},
     {stq_14_bits_uop_ppred_busy},
     {stq_13_bits_uop_ppred_busy},
     {stq_12_bits_uop_ppred_busy},
     {stq_11_bits_uop_ppred_busy},
     {stq_10_bits_uop_ppred_busy},
     {stq_9_bits_uop_ppred_busy},
     {stq_8_bits_uop_ppred_busy},
     {stq_7_bits_uop_ppred_busy},
     {stq_6_bits_uop_ppred_busy},
     {stq_5_bits_uop_ppred_busy},
     {stq_4_bits_uop_ppred_busy},
     {stq_3_bits_uop_ppred_busy},
     {stq_2_bits_uop_ppred_busy},
     {stq_1_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy}};	// lsu.scala:211:16, :224:42
  wire [31:0][6:0]  _GEN_49 =
    {{stq_0_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst},
     {stq_23_bits_uop_stale_pdst},
     {stq_22_bits_uop_stale_pdst},
     {stq_21_bits_uop_stale_pdst},
     {stq_20_bits_uop_stale_pdst},
     {stq_19_bits_uop_stale_pdst},
     {stq_18_bits_uop_stale_pdst},
     {stq_17_bits_uop_stale_pdst},
     {stq_16_bits_uop_stale_pdst},
     {stq_15_bits_uop_stale_pdst},
     {stq_14_bits_uop_stale_pdst},
     {stq_13_bits_uop_stale_pdst},
     {stq_12_bits_uop_stale_pdst},
     {stq_11_bits_uop_stale_pdst},
     {stq_10_bits_uop_stale_pdst},
     {stq_9_bits_uop_stale_pdst},
     {stq_8_bits_uop_stale_pdst},
     {stq_7_bits_uop_stale_pdst},
     {stq_6_bits_uop_stale_pdst},
     {stq_5_bits_uop_stale_pdst},
     {stq_4_bits_uop_stale_pdst},
     {stq_3_bits_uop_stale_pdst},
     {stq_2_bits_uop_stale_pdst},
     {stq_1_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_50 =
    {{stq_0_bits_uop_exception},
     {stq_0_bits_uop_exception},
     {stq_0_bits_uop_exception},
     {stq_0_bits_uop_exception},
     {stq_0_bits_uop_exception},
     {stq_0_bits_uop_exception},
     {stq_0_bits_uop_exception},
     {stq_0_bits_uop_exception},
     {stq_23_bits_uop_exception},
     {stq_22_bits_uop_exception},
     {stq_21_bits_uop_exception},
     {stq_20_bits_uop_exception},
     {stq_19_bits_uop_exception},
     {stq_18_bits_uop_exception},
     {stq_17_bits_uop_exception},
     {stq_16_bits_uop_exception},
     {stq_15_bits_uop_exception},
     {stq_14_bits_uop_exception},
     {stq_13_bits_uop_exception},
     {stq_12_bits_uop_exception},
     {stq_11_bits_uop_exception},
     {stq_10_bits_uop_exception},
     {stq_9_bits_uop_exception},
     {stq_8_bits_uop_exception},
     {stq_7_bits_uop_exception},
     {stq_6_bits_uop_exception},
     {stq_5_bits_uop_exception},
     {stq_4_bits_uop_exception},
     {stq_3_bits_uop_exception},
     {stq_2_bits_uop_exception},
     {stq_1_bits_uop_exception},
     {stq_0_bits_uop_exception}};	// lsu.scala:211:16, :224:42
  wire              _GEN_51 = _GEN_50[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [31:0][63:0] _GEN_52 =
    {{stq_0_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause},
     {stq_23_bits_uop_exc_cause},
     {stq_22_bits_uop_exc_cause},
     {stq_21_bits_uop_exc_cause},
     {stq_20_bits_uop_exc_cause},
     {stq_19_bits_uop_exc_cause},
     {stq_18_bits_uop_exc_cause},
     {stq_17_bits_uop_exc_cause},
     {stq_16_bits_uop_exc_cause},
     {stq_15_bits_uop_exc_cause},
     {stq_14_bits_uop_exc_cause},
     {stq_13_bits_uop_exc_cause},
     {stq_12_bits_uop_exc_cause},
     {stq_11_bits_uop_exc_cause},
     {stq_10_bits_uop_exc_cause},
     {stq_9_bits_uop_exc_cause},
     {stq_8_bits_uop_exc_cause},
     {stq_7_bits_uop_exc_cause},
     {stq_6_bits_uop_exc_cause},
     {stq_5_bits_uop_exc_cause},
     {stq_4_bits_uop_exc_cause},
     {stq_3_bits_uop_exc_cause},
     {stq_2_bits_uop_exc_cause},
     {stq_1_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_53 =
    {{stq_0_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable},
     {stq_23_bits_uop_bypassable},
     {stq_22_bits_uop_bypassable},
     {stq_21_bits_uop_bypassable},
     {stq_20_bits_uop_bypassable},
     {stq_19_bits_uop_bypassable},
     {stq_18_bits_uop_bypassable},
     {stq_17_bits_uop_bypassable},
     {stq_16_bits_uop_bypassable},
     {stq_15_bits_uop_bypassable},
     {stq_14_bits_uop_bypassable},
     {stq_13_bits_uop_bypassable},
     {stq_12_bits_uop_bypassable},
     {stq_11_bits_uop_bypassable},
     {stq_10_bits_uop_bypassable},
     {stq_9_bits_uop_bypassable},
     {stq_8_bits_uop_bypassable},
     {stq_7_bits_uop_bypassable},
     {stq_6_bits_uop_bypassable},
     {stq_5_bits_uop_bypassable},
     {stq_4_bits_uop_bypassable},
     {stq_3_bits_uop_bypassable},
     {stq_2_bits_uop_bypassable},
     {stq_1_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable}};	// lsu.scala:211:16, :224:42
  wire [31:0][4:0]  _GEN_54 =
    {{stq_0_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd},
     {stq_23_bits_uop_mem_cmd},
     {stq_22_bits_uop_mem_cmd},
     {stq_21_bits_uop_mem_cmd},
     {stq_20_bits_uop_mem_cmd},
     {stq_19_bits_uop_mem_cmd},
     {stq_18_bits_uop_mem_cmd},
     {stq_17_bits_uop_mem_cmd},
     {stq_16_bits_uop_mem_cmd},
     {stq_15_bits_uop_mem_cmd},
     {stq_14_bits_uop_mem_cmd},
     {stq_13_bits_uop_mem_cmd},
     {stq_12_bits_uop_mem_cmd},
     {stq_11_bits_uop_mem_cmd},
     {stq_10_bits_uop_mem_cmd},
     {stq_9_bits_uop_mem_cmd},
     {stq_8_bits_uop_mem_cmd},
     {stq_7_bits_uop_mem_cmd},
     {stq_6_bits_uop_mem_cmd},
     {stq_5_bits_uop_mem_cmd},
     {stq_4_bits_uop_mem_cmd},
     {stq_3_bits_uop_mem_cmd},
     {stq_2_bits_uop_mem_cmd},
     {stq_1_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_55 =
    {{stq_0_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size},
     {stq_23_bits_uop_mem_size},
     {stq_22_bits_uop_mem_size},
     {stq_21_bits_uop_mem_size},
     {stq_20_bits_uop_mem_size},
     {stq_19_bits_uop_mem_size},
     {stq_18_bits_uop_mem_size},
     {stq_17_bits_uop_mem_size},
     {stq_16_bits_uop_mem_size},
     {stq_15_bits_uop_mem_size},
     {stq_14_bits_uop_mem_size},
     {stq_13_bits_uop_mem_size},
     {stq_12_bits_uop_mem_size},
     {stq_11_bits_uop_mem_size},
     {stq_10_bits_uop_mem_size},
     {stq_9_bits_uop_mem_size},
     {stq_8_bits_uop_mem_size},
     {stq_7_bits_uop_mem_size},
     {stq_6_bits_uop_mem_size},
     {stq_5_bits_uop_mem_size},
     {stq_4_bits_uop_mem_size},
     {stq_3_bits_uop_mem_size},
     {stq_2_bits_uop_mem_size},
     {stq_1_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size}};	// lsu.scala:211:16, :224:42
  wire [1:0]        _GEN_56 = _GEN_55[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [31:0]       _GEN_57 =
    {{stq_0_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed},
     {stq_23_bits_uop_mem_signed},
     {stq_22_bits_uop_mem_signed},
     {stq_21_bits_uop_mem_signed},
     {stq_20_bits_uop_mem_signed},
     {stq_19_bits_uop_mem_signed},
     {stq_18_bits_uop_mem_signed},
     {stq_17_bits_uop_mem_signed},
     {stq_16_bits_uop_mem_signed},
     {stq_15_bits_uop_mem_signed},
     {stq_14_bits_uop_mem_signed},
     {stq_13_bits_uop_mem_signed},
     {stq_12_bits_uop_mem_signed},
     {stq_11_bits_uop_mem_signed},
     {stq_10_bits_uop_mem_signed},
     {stq_9_bits_uop_mem_signed},
     {stq_8_bits_uop_mem_signed},
     {stq_7_bits_uop_mem_signed},
     {stq_6_bits_uop_mem_signed},
     {stq_5_bits_uop_mem_signed},
     {stq_4_bits_uop_mem_signed},
     {stq_3_bits_uop_mem_signed},
     {stq_2_bits_uop_mem_signed},
     {stq_1_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_58 =
    {{stq_0_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence},
     {stq_23_bits_uop_is_fence},
     {stq_22_bits_uop_is_fence},
     {stq_21_bits_uop_is_fence},
     {stq_20_bits_uop_is_fence},
     {stq_19_bits_uop_is_fence},
     {stq_18_bits_uop_is_fence},
     {stq_17_bits_uop_is_fence},
     {stq_16_bits_uop_is_fence},
     {stq_15_bits_uop_is_fence},
     {stq_14_bits_uop_is_fence},
     {stq_13_bits_uop_is_fence},
     {stq_12_bits_uop_is_fence},
     {stq_11_bits_uop_is_fence},
     {stq_10_bits_uop_is_fence},
     {stq_9_bits_uop_is_fence},
     {stq_8_bits_uop_is_fence},
     {stq_7_bits_uop_is_fence},
     {stq_6_bits_uop_is_fence},
     {stq_5_bits_uop_is_fence},
     {stq_4_bits_uop_is_fence},
     {stq_3_bits_uop_is_fence},
     {stq_2_bits_uop_is_fence},
     {stq_1_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence}};	// lsu.scala:211:16, :224:42
  wire              _GEN_59 = _GEN_58[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [31:0]       _GEN_60 =
    {{stq_0_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei},
     {stq_23_bits_uop_is_fencei},
     {stq_22_bits_uop_is_fencei},
     {stq_21_bits_uop_is_fencei},
     {stq_20_bits_uop_is_fencei},
     {stq_19_bits_uop_is_fencei},
     {stq_18_bits_uop_is_fencei},
     {stq_17_bits_uop_is_fencei},
     {stq_16_bits_uop_is_fencei},
     {stq_15_bits_uop_is_fencei},
     {stq_14_bits_uop_is_fencei},
     {stq_13_bits_uop_is_fencei},
     {stq_12_bits_uop_is_fencei},
     {stq_11_bits_uop_is_fencei},
     {stq_10_bits_uop_is_fencei},
     {stq_9_bits_uop_is_fencei},
     {stq_8_bits_uop_is_fencei},
     {stq_7_bits_uop_is_fencei},
     {stq_6_bits_uop_is_fencei},
     {stq_5_bits_uop_is_fencei},
     {stq_4_bits_uop_is_fencei},
     {stq_3_bits_uop_is_fencei},
     {stq_2_bits_uop_is_fencei},
     {stq_1_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_61 =
    {{stq_0_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo},
     {stq_23_bits_uop_is_amo},
     {stq_22_bits_uop_is_amo},
     {stq_21_bits_uop_is_amo},
     {stq_20_bits_uop_is_amo},
     {stq_19_bits_uop_is_amo},
     {stq_18_bits_uop_is_amo},
     {stq_17_bits_uop_is_amo},
     {stq_16_bits_uop_is_amo},
     {stq_15_bits_uop_is_amo},
     {stq_14_bits_uop_is_amo},
     {stq_13_bits_uop_is_amo},
     {stq_12_bits_uop_is_amo},
     {stq_11_bits_uop_is_amo},
     {stq_10_bits_uop_is_amo},
     {stq_9_bits_uop_is_amo},
     {stq_8_bits_uop_is_amo},
     {stq_7_bits_uop_is_amo},
     {stq_6_bits_uop_is_amo},
     {stq_5_bits_uop_is_amo},
     {stq_4_bits_uop_is_amo},
     {stq_3_bits_uop_is_amo},
     {stq_2_bits_uop_is_amo},
     {stq_1_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo}};	// lsu.scala:211:16, :224:42
  wire              _GEN_62 = _GEN_61[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [31:0]       _GEN_63 =
    {{stq_0_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq},
     {stq_23_bits_uop_uses_ldq},
     {stq_22_bits_uop_uses_ldq},
     {stq_21_bits_uop_uses_ldq},
     {stq_20_bits_uop_uses_ldq},
     {stq_19_bits_uop_uses_ldq},
     {stq_18_bits_uop_uses_ldq},
     {stq_17_bits_uop_uses_ldq},
     {stq_16_bits_uop_uses_ldq},
     {stq_15_bits_uop_uses_ldq},
     {stq_14_bits_uop_uses_ldq},
     {stq_13_bits_uop_uses_ldq},
     {stq_12_bits_uop_uses_ldq},
     {stq_11_bits_uop_uses_ldq},
     {stq_10_bits_uop_uses_ldq},
     {stq_9_bits_uop_uses_ldq},
     {stq_8_bits_uop_uses_ldq},
     {stq_7_bits_uop_uses_ldq},
     {stq_6_bits_uop_uses_ldq},
     {stq_5_bits_uop_uses_ldq},
     {stq_4_bits_uop_uses_ldq},
     {stq_3_bits_uop_uses_ldq},
     {stq_2_bits_uop_uses_ldq},
     {stq_1_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_64 =
    {{stq_0_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq},
     {stq_23_bits_uop_uses_stq},
     {stq_22_bits_uop_uses_stq},
     {stq_21_bits_uop_uses_stq},
     {stq_20_bits_uop_uses_stq},
     {stq_19_bits_uop_uses_stq},
     {stq_18_bits_uop_uses_stq},
     {stq_17_bits_uop_uses_stq},
     {stq_16_bits_uop_uses_stq},
     {stq_15_bits_uop_uses_stq},
     {stq_14_bits_uop_uses_stq},
     {stq_13_bits_uop_uses_stq},
     {stq_12_bits_uop_uses_stq},
     {stq_11_bits_uop_uses_stq},
     {stq_10_bits_uop_uses_stq},
     {stq_9_bits_uop_uses_stq},
     {stq_8_bits_uop_uses_stq},
     {stq_7_bits_uop_uses_stq},
     {stq_6_bits_uop_uses_stq},
     {stq_5_bits_uop_uses_stq},
     {stq_4_bits_uop_uses_stq},
     {stq_3_bits_uop_uses_stq},
     {stq_2_bits_uop_uses_stq},
     {stq_1_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_65 =
    {{stq_0_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc},
     {stq_23_bits_uop_is_sys_pc2epc},
     {stq_22_bits_uop_is_sys_pc2epc},
     {stq_21_bits_uop_is_sys_pc2epc},
     {stq_20_bits_uop_is_sys_pc2epc},
     {stq_19_bits_uop_is_sys_pc2epc},
     {stq_18_bits_uop_is_sys_pc2epc},
     {stq_17_bits_uop_is_sys_pc2epc},
     {stq_16_bits_uop_is_sys_pc2epc},
     {stq_15_bits_uop_is_sys_pc2epc},
     {stq_14_bits_uop_is_sys_pc2epc},
     {stq_13_bits_uop_is_sys_pc2epc},
     {stq_12_bits_uop_is_sys_pc2epc},
     {stq_11_bits_uop_is_sys_pc2epc},
     {stq_10_bits_uop_is_sys_pc2epc},
     {stq_9_bits_uop_is_sys_pc2epc},
     {stq_8_bits_uop_is_sys_pc2epc},
     {stq_7_bits_uop_is_sys_pc2epc},
     {stq_6_bits_uop_is_sys_pc2epc},
     {stq_5_bits_uop_is_sys_pc2epc},
     {stq_4_bits_uop_is_sys_pc2epc},
     {stq_3_bits_uop_is_sys_pc2epc},
     {stq_2_bits_uop_is_sys_pc2epc},
     {stq_1_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_66 =
    {{stq_0_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique},
     {stq_23_bits_uop_is_unique},
     {stq_22_bits_uop_is_unique},
     {stq_21_bits_uop_is_unique},
     {stq_20_bits_uop_is_unique},
     {stq_19_bits_uop_is_unique},
     {stq_18_bits_uop_is_unique},
     {stq_17_bits_uop_is_unique},
     {stq_16_bits_uop_is_unique},
     {stq_15_bits_uop_is_unique},
     {stq_14_bits_uop_is_unique},
     {stq_13_bits_uop_is_unique},
     {stq_12_bits_uop_is_unique},
     {stq_11_bits_uop_is_unique},
     {stq_10_bits_uop_is_unique},
     {stq_9_bits_uop_is_unique},
     {stq_8_bits_uop_is_unique},
     {stq_7_bits_uop_is_unique},
     {stq_6_bits_uop_is_unique},
     {stq_5_bits_uop_is_unique},
     {stq_4_bits_uop_is_unique},
     {stq_3_bits_uop_is_unique},
     {stq_2_bits_uop_is_unique},
     {stq_1_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_67 =
    {{stq_0_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit},
     {stq_23_bits_uop_flush_on_commit},
     {stq_22_bits_uop_flush_on_commit},
     {stq_21_bits_uop_flush_on_commit},
     {stq_20_bits_uop_flush_on_commit},
     {stq_19_bits_uop_flush_on_commit},
     {stq_18_bits_uop_flush_on_commit},
     {stq_17_bits_uop_flush_on_commit},
     {stq_16_bits_uop_flush_on_commit},
     {stq_15_bits_uop_flush_on_commit},
     {stq_14_bits_uop_flush_on_commit},
     {stq_13_bits_uop_flush_on_commit},
     {stq_12_bits_uop_flush_on_commit},
     {stq_11_bits_uop_flush_on_commit},
     {stq_10_bits_uop_flush_on_commit},
     {stq_9_bits_uop_flush_on_commit},
     {stq_8_bits_uop_flush_on_commit},
     {stq_7_bits_uop_flush_on_commit},
     {stq_6_bits_uop_flush_on_commit},
     {stq_5_bits_uop_flush_on_commit},
     {stq_4_bits_uop_flush_on_commit},
     {stq_3_bits_uop_flush_on_commit},
     {stq_2_bits_uop_flush_on_commit},
     {stq_1_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_68 =
    {{stq_0_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1},
     {stq_23_bits_uop_ldst_is_rs1},
     {stq_22_bits_uop_ldst_is_rs1},
     {stq_21_bits_uop_ldst_is_rs1},
     {stq_20_bits_uop_ldst_is_rs1},
     {stq_19_bits_uop_ldst_is_rs1},
     {stq_18_bits_uop_ldst_is_rs1},
     {stq_17_bits_uop_ldst_is_rs1},
     {stq_16_bits_uop_ldst_is_rs1},
     {stq_15_bits_uop_ldst_is_rs1},
     {stq_14_bits_uop_ldst_is_rs1},
     {stq_13_bits_uop_ldst_is_rs1},
     {stq_12_bits_uop_ldst_is_rs1},
     {stq_11_bits_uop_ldst_is_rs1},
     {stq_10_bits_uop_ldst_is_rs1},
     {stq_9_bits_uop_ldst_is_rs1},
     {stq_8_bits_uop_ldst_is_rs1},
     {stq_7_bits_uop_ldst_is_rs1},
     {stq_6_bits_uop_ldst_is_rs1},
     {stq_5_bits_uop_ldst_is_rs1},
     {stq_4_bits_uop_ldst_is_rs1},
     {stq_3_bits_uop_ldst_is_rs1},
     {stq_2_bits_uop_ldst_is_rs1},
     {stq_1_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1}};	// lsu.scala:211:16, :224:42
  wire [31:0][5:0]  _GEN_69 =
    {{stq_0_bits_uop_ldst},
     {stq_0_bits_uop_ldst},
     {stq_0_bits_uop_ldst},
     {stq_0_bits_uop_ldst},
     {stq_0_bits_uop_ldst},
     {stq_0_bits_uop_ldst},
     {stq_0_bits_uop_ldst},
     {stq_0_bits_uop_ldst},
     {stq_23_bits_uop_ldst},
     {stq_22_bits_uop_ldst},
     {stq_21_bits_uop_ldst},
     {stq_20_bits_uop_ldst},
     {stq_19_bits_uop_ldst},
     {stq_18_bits_uop_ldst},
     {stq_17_bits_uop_ldst},
     {stq_16_bits_uop_ldst},
     {stq_15_bits_uop_ldst},
     {stq_14_bits_uop_ldst},
     {stq_13_bits_uop_ldst},
     {stq_12_bits_uop_ldst},
     {stq_11_bits_uop_ldst},
     {stq_10_bits_uop_ldst},
     {stq_9_bits_uop_ldst},
     {stq_8_bits_uop_ldst},
     {stq_7_bits_uop_ldst},
     {stq_6_bits_uop_ldst},
     {stq_5_bits_uop_ldst},
     {stq_4_bits_uop_ldst},
     {stq_3_bits_uop_ldst},
     {stq_2_bits_uop_ldst},
     {stq_1_bits_uop_ldst},
     {stq_0_bits_uop_ldst}};	// lsu.scala:211:16, :224:42
  wire [31:0][5:0]  _GEN_70 =
    {{stq_0_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1},
     {stq_23_bits_uop_lrs1},
     {stq_22_bits_uop_lrs1},
     {stq_21_bits_uop_lrs1},
     {stq_20_bits_uop_lrs1},
     {stq_19_bits_uop_lrs1},
     {stq_18_bits_uop_lrs1},
     {stq_17_bits_uop_lrs1},
     {stq_16_bits_uop_lrs1},
     {stq_15_bits_uop_lrs1},
     {stq_14_bits_uop_lrs1},
     {stq_13_bits_uop_lrs1},
     {stq_12_bits_uop_lrs1},
     {stq_11_bits_uop_lrs1},
     {stq_10_bits_uop_lrs1},
     {stq_9_bits_uop_lrs1},
     {stq_8_bits_uop_lrs1},
     {stq_7_bits_uop_lrs1},
     {stq_6_bits_uop_lrs1},
     {stq_5_bits_uop_lrs1},
     {stq_4_bits_uop_lrs1},
     {stq_3_bits_uop_lrs1},
     {stq_2_bits_uop_lrs1},
     {stq_1_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1}};	// lsu.scala:211:16, :224:42
  wire [31:0][5:0]  _GEN_71 =
    {{stq_0_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2},
     {stq_23_bits_uop_lrs2},
     {stq_22_bits_uop_lrs2},
     {stq_21_bits_uop_lrs2},
     {stq_20_bits_uop_lrs2},
     {stq_19_bits_uop_lrs2},
     {stq_18_bits_uop_lrs2},
     {stq_17_bits_uop_lrs2},
     {stq_16_bits_uop_lrs2},
     {stq_15_bits_uop_lrs2},
     {stq_14_bits_uop_lrs2},
     {stq_13_bits_uop_lrs2},
     {stq_12_bits_uop_lrs2},
     {stq_11_bits_uop_lrs2},
     {stq_10_bits_uop_lrs2},
     {stq_9_bits_uop_lrs2},
     {stq_8_bits_uop_lrs2},
     {stq_7_bits_uop_lrs2},
     {stq_6_bits_uop_lrs2},
     {stq_5_bits_uop_lrs2},
     {stq_4_bits_uop_lrs2},
     {stq_3_bits_uop_lrs2},
     {stq_2_bits_uop_lrs2},
     {stq_1_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2}};	// lsu.scala:211:16, :224:42
  wire [31:0][5:0]  _GEN_72 =
    {{stq_0_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3},
     {stq_23_bits_uop_lrs3},
     {stq_22_bits_uop_lrs3},
     {stq_21_bits_uop_lrs3},
     {stq_20_bits_uop_lrs3},
     {stq_19_bits_uop_lrs3},
     {stq_18_bits_uop_lrs3},
     {stq_17_bits_uop_lrs3},
     {stq_16_bits_uop_lrs3},
     {stq_15_bits_uop_lrs3},
     {stq_14_bits_uop_lrs3},
     {stq_13_bits_uop_lrs3},
     {stq_12_bits_uop_lrs3},
     {stq_11_bits_uop_lrs3},
     {stq_10_bits_uop_lrs3},
     {stq_9_bits_uop_lrs3},
     {stq_8_bits_uop_lrs3},
     {stq_7_bits_uop_lrs3},
     {stq_6_bits_uop_lrs3},
     {stq_5_bits_uop_lrs3},
     {stq_4_bits_uop_lrs3},
     {stq_3_bits_uop_lrs3},
     {stq_2_bits_uop_lrs3},
     {stq_1_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_73 =
    {{stq_0_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val},
     {stq_23_bits_uop_ldst_val},
     {stq_22_bits_uop_ldst_val},
     {stq_21_bits_uop_ldst_val},
     {stq_20_bits_uop_ldst_val},
     {stq_19_bits_uop_ldst_val},
     {stq_18_bits_uop_ldst_val},
     {stq_17_bits_uop_ldst_val},
     {stq_16_bits_uop_ldst_val},
     {stq_15_bits_uop_ldst_val},
     {stq_14_bits_uop_ldst_val},
     {stq_13_bits_uop_ldst_val},
     {stq_12_bits_uop_ldst_val},
     {stq_11_bits_uop_ldst_val},
     {stq_10_bits_uop_ldst_val},
     {stq_9_bits_uop_ldst_val},
     {stq_8_bits_uop_ldst_val},
     {stq_7_bits_uop_ldst_val},
     {stq_6_bits_uop_ldst_val},
     {stq_5_bits_uop_ldst_val},
     {stq_4_bits_uop_ldst_val},
     {stq_3_bits_uop_ldst_val},
     {stq_2_bits_uop_ldst_val},
     {stq_1_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_74 =
    {{stq_0_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype},
     {stq_23_bits_uop_dst_rtype},
     {stq_22_bits_uop_dst_rtype},
     {stq_21_bits_uop_dst_rtype},
     {stq_20_bits_uop_dst_rtype},
     {stq_19_bits_uop_dst_rtype},
     {stq_18_bits_uop_dst_rtype},
     {stq_17_bits_uop_dst_rtype},
     {stq_16_bits_uop_dst_rtype},
     {stq_15_bits_uop_dst_rtype},
     {stq_14_bits_uop_dst_rtype},
     {stq_13_bits_uop_dst_rtype},
     {stq_12_bits_uop_dst_rtype},
     {stq_11_bits_uop_dst_rtype},
     {stq_10_bits_uop_dst_rtype},
     {stq_9_bits_uop_dst_rtype},
     {stq_8_bits_uop_dst_rtype},
     {stq_7_bits_uop_dst_rtype},
     {stq_6_bits_uop_dst_rtype},
     {stq_5_bits_uop_dst_rtype},
     {stq_4_bits_uop_dst_rtype},
     {stq_3_bits_uop_dst_rtype},
     {stq_2_bits_uop_dst_rtype},
     {stq_1_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_75 =
    {{stq_0_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype},
     {stq_23_bits_uop_lrs1_rtype},
     {stq_22_bits_uop_lrs1_rtype},
     {stq_21_bits_uop_lrs1_rtype},
     {stq_20_bits_uop_lrs1_rtype},
     {stq_19_bits_uop_lrs1_rtype},
     {stq_18_bits_uop_lrs1_rtype},
     {stq_17_bits_uop_lrs1_rtype},
     {stq_16_bits_uop_lrs1_rtype},
     {stq_15_bits_uop_lrs1_rtype},
     {stq_14_bits_uop_lrs1_rtype},
     {stq_13_bits_uop_lrs1_rtype},
     {stq_12_bits_uop_lrs1_rtype},
     {stq_11_bits_uop_lrs1_rtype},
     {stq_10_bits_uop_lrs1_rtype},
     {stq_9_bits_uop_lrs1_rtype},
     {stq_8_bits_uop_lrs1_rtype},
     {stq_7_bits_uop_lrs1_rtype},
     {stq_6_bits_uop_lrs1_rtype},
     {stq_5_bits_uop_lrs1_rtype},
     {stq_4_bits_uop_lrs1_rtype},
     {stq_3_bits_uop_lrs1_rtype},
     {stq_2_bits_uop_lrs1_rtype},
     {stq_1_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_76 =
    {{stq_0_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype},
     {stq_23_bits_uop_lrs2_rtype},
     {stq_22_bits_uop_lrs2_rtype},
     {stq_21_bits_uop_lrs2_rtype},
     {stq_20_bits_uop_lrs2_rtype},
     {stq_19_bits_uop_lrs2_rtype},
     {stq_18_bits_uop_lrs2_rtype},
     {stq_17_bits_uop_lrs2_rtype},
     {stq_16_bits_uop_lrs2_rtype},
     {stq_15_bits_uop_lrs2_rtype},
     {stq_14_bits_uop_lrs2_rtype},
     {stq_13_bits_uop_lrs2_rtype},
     {stq_12_bits_uop_lrs2_rtype},
     {stq_11_bits_uop_lrs2_rtype},
     {stq_10_bits_uop_lrs2_rtype},
     {stq_9_bits_uop_lrs2_rtype},
     {stq_8_bits_uop_lrs2_rtype},
     {stq_7_bits_uop_lrs2_rtype},
     {stq_6_bits_uop_lrs2_rtype},
     {stq_5_bits_uop_lrs2_rtype},
     {stq_4_bits_uop_lrs2_rtype},
     {stq_3_bits_uop_lrs2_rtype},
     {stq_2_bits_uop_lrs2_rtype},
     {stq_1_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_77 =
    {{stq_0_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en},
     {stq_23_bits_uop_frs3_en},
     {stq_22_bits_uop_frs3_en},
     {stq_21_bits_uop_frs3_en},
     {stq_20_bits_uop_frs3_en},
     {stq_19_bits_uop_frs3_en},
     {stq_18_bits_uop_frs3_en},
     {stq_17_bits_uop_frs3_en},
     {stq_16_bits_uop_frs3_en},
     {stq_15_bits_uop_frs3_en},
     {stq_14_bits_uop_frs3_en},
     {stq_13_bits_uop_frs3_en},
     {stq_12_bits_uop_frs3_en},
     {stq_11_bits_uop_frs3_en},
     {stq_10_bits_uop_frs3_en},
     {stq_9_bits_uop_frs3_en},
     {stq_8_bits_uop_frs3_en},
     {stq_7_bits_uop_frs3_en},
     {stq_6_bits_uop_frs3_en},
     {stq_5_bits_uop_frs3_en},
     {stq_4_bits_uop_frs3_en},
     {stq_3_bits_uop_frs3_en},
     {stq_2_bits_uop_frs3_en},
     {stq_1_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_78 =
    {{stq_0_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val},
     {stq_23_bits_uop_fp_val},
     {stq_22_bits_uop_fp_val},
     {stq_21_bits_uop_fp_val},
     {stq_20_bits_uop_fp_val},
     {stq_19_bits_uop_fp_val},
     {stq_18_bits_uop_fp_val},
     {stq_17_bits_uop_fp_val},
     {stq_16_bits_uop_fp_val},
     {stq_15_bits_uop_fp_val},
     {stq_14_bits_uop_fp_val},
     {stq_13_bits_uop_fp_val},
     {stq_12_bits_uop_fp_val},
     {stq_11_bits_uop_fp_val},
     {stq_10_bits_uop_fp_val},
     {stq_9_bits_uop_fp_val},
     {stq_8_bits_uop_fp_val},
     {stq_7_bits_uop_fp_val},
     {stq_6_bits_uop_fp_val},
     {stq_5_bits_uop_fp_val},
     {stq_4_bits_uop_fp_val},
     {stq_3_bits_uop_fp_val},
     {stq_2_bits_uop_fp_val},
     {stq_1_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_79 =
    {{stq_0_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single},
     {stq_23_bits_uop_fp_single},
     {stq_22_bits_uop_fp_single},
     {stq_21_bits_uop_fp_single},
     {stq_20_bits_uop_fp_single},
     {stq_19_bits_uop_fp_single},
     {stq_18_bits_uop_fp_single},
     {stq_17_bits_uop_fp_single},
     {stq_16_bits_uop_fp_single},
     {stq_15_bits_uop_fp_single},
     {stq_14_bits_uop_fp_single},
     {stq_13_bits_uop_fp_single},
     {stq_12_bits_uop_fp_single},
     {stq_11_bits_uop_fp_single},
     {stq_10_bits_uop_fp_single},
     {stq_9_bits_uop_fp_single},
     {stq_8_bits_uop_fp_single},
     {stq_7_bits_uop_fp_single},
     {stq_6_bits_uop_fp_single},
     {stq_5_bits_uop_fp_single},
     {stq_4_bits_uop_fp_single},
     {stq_3_bits_uop_fp_single},
     {stq_2_bits_uop_fp_single},
     {stq_1_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_80 =
    {{stq_0_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if},
     {stq_23_bits_uop_xcpt_pf_if},
     {stq_22_bits_uop_xcpt_pf_if},
     {stq_21_bits_uop_xcpt_pf_if},
     {stq_20_bits_uop_xcpt_pf_if},
     {stq_19_bits_uop_xcpt_pf_if},
     {stq_18_bits_uop_xcpt_pf_if},
     {stq_17_bits_uop_xcpt_pf_if},
     {stq_16_bits_uop_xcpt_pf_if},
     {stq_15_bits_uop_xcpt_pf_if},
     {stq_14_bits_uop_xcpt_pf_if},
     {stq_13_bits_uop_xcpt_pf_if},
     {stq_12_bits_uop_xcpt_pf_if},
     {stq_11_bits_uop_xcpt_pf_if},
     {stq_10_bits_uop_xcpt_pf_if},
     {stq_9_bits_uop_xcpt_pf_if},
     {stq_8_bits_uop_xcpt_pf_if},
     {stq_7_bits_uop_xcpt_pf_if},
     {stq_6_bits_uop_xcpt_pf_if},
     {stq_5_bits_uop_xcpt_pf_if},
     {stq_4_bits_uop_xcpt_pf_if},
     {stq_3_bits_uop_xcpt_pf_if},
     {stq_2_bits_uop_xcpt_pf_if},
     {stq_1_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_81 =
    {{stq_0_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if},
     {stq_23_bits_uop_xcpt_ae_if},
     {stq_22_bits_uop_xcpt_ae_if},
     {stq_21_bits_uop_xcpt_ae_if},
     {stq_20_bits_uop_xcpt_ae_if},
     {stq_19_bits_uop_xcpt_ae_if},
     {stq_18_bits_uop_xcpt_ae_if},
     {stq_17_bits_uop_xcpt_ae_if},
     {stq_16_bits_uop_xcpt_ae_if},
     {stq_15_bits_uop_xcpt_ae_if},
     {stq_14_bits_uop_xcpt_ae_if},
     {stq_13_bits_uop_xcpt_ae_if},
     {stq_12_bits_uop_xcpt_ae_if},
     {stq_11_bits_uop_xcpt_ae_if},
     {stq_10_bits_uop_xcpt_ae_if},
     {stq_9_bits_uop_xcpt_ae_if},
     {stq_8_bits_uop_xcpt_ae_if},
     {stq_7_bits_uop_xcpt_ae_if},
     {stq_6_bits_uop_xcpt_ae_if},
     {stq_5_bits_uop_xcpt_ae_if},
     {stq_4_bits_uop_xcpt_ae_if},
     {stq_3_bits_uop_xcpt_ae_if},
     {stq_2_bits_uop_xcpt_ae_if},
     {stq_1_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_82 =
    {{stq_0_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if},
     {stq_23_bits_uop_xcpt_ma_if},
     {stq_22_bits_uop_xcpt_ma_if},
     {stq_21_bits_uop_xcpt_ma_if},
     {stq_20_bits_uop_xcpt_ma_if},
     {stq_19_bits_uop_xcpt_ma_if},
     {stq_18_bits_uop_xcpt_ma_if},
     {stq_17_bits_uop_xcpt_ma_if},
     {stq_16_bits_uop_xcpt_ma_if},
     {stq_15_bits_uop_xcpt_ma_if},
     {stq_14_bits_uop_xcpt_ma_if},
     {stq_13_bits_uop_xcpt_ma_if},
     {stq_12_bits_uop_xcpt_ma_if},
     {stq_11_bits_uop_xcpt_ma_if},
     {stq_10_bits_uop_xcpt_ma_if},
     {stq_9_bits_uop_xcpt_ma_if},
     {stq_8_bits_uop_xcpt_ma_if},
     {stq_7_bits_uop_xcpt_ma_if},
     {stq_6_bits_uop_xcpt_ma_if},
     {stq_5_bits_uop_xcpt_ma_if},
     {stq_4_bits_uop_xcpt_ma_if},
     {stq_3_bits_uop_xcpt_ma_if},
     {stq_2_bits_uop_xcpt_ma_if},
     {stq_1_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_83 =
    {{stq_0_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if},
     {stq_23_bits_uop_bp_debug_if},
     {stq_22_bits_uop_bp_debug_if},
     {stq_21_bits_uop_bp_debug_if},
     {stq_20_bits_uop_bp_debug_if},
     {stq_19_bits_uop_bp_debug_if},
     {stq_18_bits_uop_bp_debug_if},
     {stq_17_bits_uop_bp_debug_if},
     {stq_16_bits_uop_bp_debug_if},
     {stq_15_bits_uop_bp_debug_if},
     {stq_14_bits_uop_bp_debug_if},
     {stq_13_bits_uop_bp_debug_if},
     {stq_12_bits_uop_bp_debug_if},
     {stq_11_bits_uop_bp_debug_if},
     {stq_10_bits_uop_bp_debug_if},
     {stq_9_bits_uop_bp_debug_if},
     {stq_8_bits_uop_bp_debug_if},
     {stq_7_bits_uop_bp_debug_if},
     {stq_6_bits_uop_bp_debug_if},
     {stq_5_bits_uop_bp_debug_if},
     {stq_4_bits_uop_bp_debug_if},
     {stq_3_bits_uop_bp_debug_if},
     {stq_2_bits_uop_bp_debug_if},
     {stq_1_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_84 =
    {{stq_0_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if},
     {stq_23_bits_uop_bp_xcpt_if},
     {stq_22_bits_uop_bp_xcpt_if},
     {stq_21_bits_uop_bp_xcpt_if},
     {stq_20_bits_uop_bp_xcpt_if},
     {stq_19_bits_uop_bp_xcpt_if},
     {stq_18_bits_uop_bp_xcpt_if},
     {stq_17_bits_uop_bp_xcpt_if},
     {stq_16_bits_uop_bp_xcpt_if},
     {stq_15_bits_uop_bp_xcpt_if},
     {stq_14_bits_uop_bp_xcpt_if},
     {stq_13_bits_uop_bp_xcpt_if},
     {stq_12_bits_uop_bp_xcpt_if},
     {stq_11_bits_uop_bp_xcpt_if},
     {stq_10_bits_uop_bp_xcpt_if},
     {stq_9_bits_uop_bp_xcpt_if},
     {stq_8_bits_uop_bp_xcpt_if},
     {stq_7_bits_uop_bp_xcpt_if},
     {stq_6_bits_uop_bp_xcpt_if},
     {stq_5_bits_uop_bp_xcpt_if},
     {stq_4_bits_uop_bp_xcpt_if},
     {stq_3_bits_uop_bp_xcpt_if},
     {stq_2_bits_uop_bp_xcpt_if},
     {stq_1_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_85 =
    {{stq_0_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc},
     {stq_23_bits_uop_debug_fsrc},
     {stq_22_bits_uop_debug_fsrc},
     {stq_21_bits_uop_debug_fsrc},
     {stq_20_bits_uop_debug_fsrc},
     {stq_19_bits_uop_debug_fsrc},
     {stq_18_bits_uop_debug_fsrc},
     {stq_17_bits_uop_debug_fsrc},
     {stq_16_bits_uop_debug_fsrc},
     {stq_15_bits_uop_debug_fsrc},
     {stq_14_bits_uop_debug_fsrc},
     {stq_13_bits_uop_debug_fsrc},
     {stq_12_bits_uop_debug_fsrc},
     {stq_11_bits_uop_debug_fsrc},
     {stq_10_bits_uop_debug_fsrc},
     {stq_9_bits_uop_debug_fsrc},
     {stq_8_bits_uop_debug_fsrc},
     {stq_7_bits_uop_debug_fsrc},
     {stq_6_bits_uop_debug_fsrc},
     {stq_5_bits_uop_debug_fsrc},
     {stq_4_bits_uop_debug_fsrc},
     {stq_3_bits_uop_debug_fsrc},
     {stq_2_bits_uop_debug_fsrc},
     {stq_1_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc}};	// lsu.scala:211:16, :224:42
  wire [31:0][1:0]  _GEN_86 =
    {{stq_0_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc},
     {stq_23_bits_uop_debug_tsrc},
     {stq_22_bits_uop_debug_tsrc},
     {stq_21_bits_uop_debug_tsrc},
     {stq_20_bits_uop_debug_tsrc},
     {stq_19_bits_uop_debug_tsrc},
     {stq_18_bits_uop_debug_tsrc},
     {stq_17_bits_uop_debug_tsrc},
     {stq_16_bits_uop_debug_tsrc},
     {stq_15_bits_uop_debug_tsrc},
     {stq_14_bits_uop_debug_tsrc},
     {stq_13_bits_uop_debug_tsrc},
     {stq_12_bits_uop_debug_tsrc},
     {stq_11_bits_uop_debug_tsrc},
     {stq_10_bits_uop_debug_tsrc},
     {stq_9_bits_uop_debug_tsrc},
     {stq_8_bits_uop_debug_tsrc},
     {stq_7_bits_uop_debug_tsrc},
     {stq_6_bits_uop_debug_tsrc},
     {stq_5_bits_uop_debug_tsrc},
     {stq_4_bits_uop_debug_tsrc},
     {stq_3_bits_uop_debug_tsrc},
     {stq_2_bits_uop_debug_tsrc},
     {stq_1_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_87 =
    {{stq_0_bits_addr_valid},
     {stq_0_bits_addr_valid},
     {stq_0_bits_addr_valid},
     {stq_0_bits_addr_valid},
     {stq_0_bits_addr_valid},
     {stq_0_bits_addr_valid},
     {stq_0_bits_addr_valid},
     {stq_0_bits_addr_valid},
     {stq_23_bits_addr_valid},
     {stq_22_bits_addr_valid},
     {stq_21_bits_addr_valid},
     {stq_20_bits_addr_valid},
     {stq_19_bits_addr_valid},
     {stq_18_bits_addr_valid},
     {stq_17_bits_addr_valid},
     {stq_16_bits_addr_valid},
     {stq_15_bits_addr_valid},
     {stq_14_bits_addr_valid},
     {stq_13_bits_addr_valid},
     {stq_12_bits_addr_valid},
     {stq_11_bits_addr_valid},
     {stq_10_bits_addr_valid},
     {stq_9_bits_addr_valid},
     {stq_8_bits_addr_valid},
     {stq_7_bits_addr_valid},
     {stq_6_bits_addr_valid},
     {stq_5_bits_addr_valid},
     {stq_4_bits_addr_valid},
     {stq_3_bits_addr_valid},
     {stq_2_bits_addr_valid},
     {stq_1_bits_addr_valid},
     {stq_0_bits_addr_valid}};	// lsu.scala:211:16, :224:42
  wire [31:0][39:0] _GEN_88 =
    {{stq_0_bits_addr_bits},
     {stq_0_bits_addr_bits},
     {stq_0_bits_addr_bits},
     {stq_0_bits_addr_bits},
     {stq_0_bits_addr_bits},
     {stq_0_bits_addr_bits},
     {stq_0_bits_addr_bits},
     {stq_0_bits_addr_bits},
     {stq_23_bits_addr_bits},
     {stq_22_bits_addr_bits},
     {stq_21_bits_addr_bits},
     {stq_20_bits_addr_bits},
     {stq_19_bits_addr_bits},
     {stq_18_bits_addr_bits},
     {stq_17_bits_addr_bits},
     {stq_16_bits_addr_bits},
     {stq_15_bits_addr_bits},
     {stq_14_bits_addr_bits},
     {stq_13_bits_addr_bits},
     {stq_12_bits_addr_bits},
     {stq_11_bits_addr_bits},
     {stq_10_bits_addr_bits},
     {stq_9_bits_addr_bits},
     {stq_8_bits_addr_bits},
     {stq_7_bits_addr_bits},
     {stq_6_bits_addr_bits},
     {stq_5_bits_addr_bits},
     {stq_4_bits_addr_bits},
     {stq_3_bits_addr_bits},
     {stq_2_bits_addr_bits},
     {stq_1_bits_addr_bits},
     {stq_0_bits_addr_bits}};	// lsu.scala:211:16, :224:42
  wire [39:0]       _GEN_89 = _GEN_88[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [31:0]       _GEN_90 =
    {{stq_0_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual},
     {stq_23_bits_addr_is_virtual},
     {stq_22_bits_addr_is_virtual},
     {stq_21_bits_addr_is_virtual},
     {stq_20_bits_addr_is_virtual},
     {stq_19_bits_addr_is_virtual},
     {stq_18_bits_addr_is_virtual},
     {stq_17_bits_addr_is_virtual},
     {stq_16_bits_addr_is_virtual},
     {stq_15_bits_addr_is_virtual},
     {stq_14_bits_addr_is_virtual},
     {stq_13_bits_addr_is_virtual},
     {stq_12_bits_addr_is_virtual},
     {stq_11_bits_addr_is_virtual},
     {stq_10_bits_addr_is_virtual},
     {stq_9_bits_addr_is_virtual},
     {stq_8_bits_addr_is_virtual},
     {stq_7_bits_addr_is_virtual},
     {stq_6_bits_addr_is_virtual},
     {stq_5_bits_addr_is_virtual},
     {stq_4_bits_addr_is_virtual},
     {stq_3_bits_addr_is_virtual},
     {stq_2_bits_addr_is_virtual},
     {stq_1_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual}};	// lsu.scala:211:16, :224:42
  wire [31:0]       _GEN_91 =
    {{stq_0_bits_data_valid},
     {stq_0_bits_data_valid},
     {stq_0_bits_data_valid},
     {stq_0_bits_data_valid},
     {stq_0_bits_data_valid},
     {stq_0_bits_data_valid},
     {stq_0_bits_data_valid},
     {stq_0_bits_data_valid},
     {stq_23_bits_data_valid},
     {stq_22_bits_data_valid},
     {stq_21_bits_data_valid},
     {stq_20_bits_data_valid},
     {stq_19_bits_data_valid},
     {stq_18_bits_data_valid},
     {stq_17_bits_data_valid},
     {stq_16_bits_data_valid},
     {stq_15_bits_data_valid},
     {stq_14_bits_data_valid},
     {stq_13_bits_data_valid},
     {stq_12_bits_data_valid},
     {stq_11_bits_data_valid},
     {stq_10_bits_data_valid},
     {stq_9_bits_data_valid},
     {stq_8_bits_data_valid},
     {stq_7_bits_data_valid},
     {stq_6_bits_data_valid},
     {stq_5_bits_data_valid},
     {stq_4_bits_data_valid},
     {stq_3_bits_data_valid},
     {stq_2_bits_data_valid},
     {stq_1_bits_data_valid},
     {stq_0_bits_data_valid}};	// lsu.scala:211:16, :224:42
  wire [31:0][63:0] _GEN_92 =
    {{stq_0_bits_data_bits},
     {stq_0_bits_data_bits},
     {stq_0_bits_data_bits},
     {stq_0_bits_data_bits},
     {stq_0_bits_data_bits},
     {stq_0_bits_data_bits},
     {stq_0_bits_data_bits},
     {stq_0_bits_data_bits},
     {stq_23_bits_data_bits},
     {stq_22_bits_data_bits},
     {stq_21_bits_data_bits},
     {stq_20_bits_data_bits},
     {stq_19_bits_data_bits},
     {stq_18_bits_data_bits},
     {stq_17_bits_data_bits},
     {stq_16_bits_data_bits},
     {stq_15_bits_data_bits},
     {stq_14_bits_data_bits},
     {stq_13_bits_data_bits},
     {stq_12_bits_data_bits},
     {stq_11_bits_data_bits},
     {stq_10_bits_data_bits},
     {stq_9_bits_data_bits},
     {stq_8_bits_data_bits},
     {stq_7_bits_data_bits},
     {stq_6_bits_data_bits},
     {stq_5_bits_data_bits},
     {stq_4_bits_data_bits},
     {stq_3_bits_data_bits},
     {stq_2_bits_data_bits},
     {stq_1_bits_data_bits},
     {stq_0_bits_data_bits}};	// lsu.scala:211:16, :224:42
  wire [63:0]       _GEN_93 = _GEN_92[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [31:0]       _GEN_94 =
    {{stq_0_bits_committed},
     {stq_0_bits_committed},
     {stq_0_bits_committed},
     {stq_0_bits_committed},
     {stq_0_bits_committed},
     {stq_0_bits_committed},
     {stq_0_bits_committed},
     {stq_0_bits_committed},
     {stq_23_bits_committed},
     {stq_22_bits_committed},
     {stq_21_bits_committed},
     {stq_20_bits_committed},
     {stq_19_bits_committed},
     {stq_18_bits_committed},
     {stq_17_bits_committed},
     {stq_16_bits_committed},
     {stq_15_bits_committed},
     {stq_14_bits_committed},
     {stq_13_bits_committed},
     {stq_12_bits_committed},
     {stq_11_bits_committed},
     {stq_10_bits_committed},
     {stq_9_bits_committed},
     {stq_8_bits_committed},
     {stq_7_bits_committed},
     {stq_6_bits_committed},
     {stq_5_bits_committed},
     {stq_4_bits_committed},
     {stq_3_bits_committed},
     {stq_2_bits_committed},
     {stq_1_bits_committed},
     {stq_0_bits_committed}};	// lsu.scala:211:16, :224:42
  reg  [2:0]        hella_state;	// lsu.scala:242:38
  reg  [39:0]       hella_req_addr;	// lsu.scala:243:34
  reg  [4:0]        hella_req_cmd;	// lsu.scala:243:34
  reg  [1:0]        hella_req_size;	// lsu.scala:243:34
  reg               hella_req_signed;	// lsu.scala:243:34
  reg               hella_req_phys;	// lsu.scala:243:34
  reg  [63:0]       hella_data_data;	// lsu.scala:244:34
  reg  [31:0]       hella_paddr;	// lsu.scala:245:34
  reg               hella_xcpt_ma_ld;	// lsu.scala:246:34
  reg               hella_xcpt_ma_st;	// lsu.scala:246:34
  reg               hella_xcpt_pf_ld;	// lsu.scala:246:34
  reg               hella_xcpt_pf_st;	// lsu.scala:246:34
  reg               hella_xcpt_ae_ld;	// lsu.scala:246:34
  reg               hella_xcpt_ae_st;	// lsu.scala:246:34
  reg  [23:0]       live_store_mask;	// lsu.scala:259:32
  wire              wrap = ldq_tail == 5'h17;	// lsu.scala:216:29, util.scala:205:25
  wire [4:0]        _GEN_95 = ldq_tail + 5'h1;	// lsu.scala:216:29, :305:44, util.scala:206:28
  wire [4:0]        _GEN_96 = wrap ? 5'h0 : _GEN_95;	// util.scala:205:25, :206:{10,28}
  wire              wrap_1 = stq_tail == 5'h17;	// lsu.scala:218:29, util.scala:205:25
  wire [4:0]        _GEN_97 = stq_tail + 5'h1;	// lsu.scala:218:29, :305:44, util.scala:206:28
  wire [4:0]        _GEN_98 = wrap_1 ? 5'h0 : _GEN_97;	// util.scala:205:25, :206:{10,28}
  wire              dis_ld_val =
    io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_ldq
    & ~io_core_dis_uops_0_bits_exception;	// lsu.scala:301:{85,88}
  wire              dis_st_val =
    io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_stq
    & ~io_core_dis_uops_0_bits_exception;	// lsu.scala:301:88, :302:85
  wire [31:0]       _GEN_99 =
    {{ldq_0_valid},
     {ldq_0_valid},
     {ldq_0_valid},
     {ldq_0_valid},
     {ldq_0_valid},
     {ldq_0_valid},
     {ldq_0_valid},
     {ldq_0_valid},
     {ldq_23_valid},
     {ldq_22_valid},
     {ldq_21_valid},
     {ldq_20_valid},
     {ldq_19_valid},
     {ldq_18_valid},
     {ldq_17_valid},
     {ldq_16_valid},
     {ldq_15_valid},
     {ldq_14_valid},
     {ldq_13_valid},
     {ldq_12_valid},
     {ldq_11_valid},
     {ldq_10_valid},
     {ldq_9_valid},
     {ldq_8_valid},
     {ldq_7_valid},
     {ldq_6_valid},
     {ldq_5_valid},
     {ldq_4_valid},
     {ldq_3_valid},
     {ldq_2_valid},
     {ldq_1_valid},
     {ldq_0_valid}};	// lsu.scala:210:16, :305:44
  wire [4:0]        _GEN_100 = dis_ld_val ? _GEN_96 : ldq_tail;	// lsu.scala:216:29, :301:85, :333:21, util.scala:206:10
  wire [4:0]        _GEN_101 = dis_st_val ? _GEN_98 : stq_tail;	// lsu.scala:218:29, :302:85, :338:21, util.scala:206:10
  wire              wrap_4 = _GEN_100 == 5'h17;	// lsu.scala:333:21, util.scala:205:25
  wire [4:0]        _GEN_102 = _GEN_100 + 5'h1;	// lsu.scala:305:44, :333:21, util.scala:206:28
  wire [4:0]        _GEN_103 = wrap_4 ? 5'h0 : _GEN_102;	// util.scala:205:25, :206:{10,28}
  wire              wrap_5 = _GEN_101 == 5'h17;	// lsu.scala:338:21, util.scala:205:25
  wire [4:0]        _GEN_104 = _GEN_101 + 5'h1;	// lsu.scala:305:44, :338:21, util.scala:206:28
  wire [4:0]        _GEN_105 = wrap_5 ? 5'h0 : _GEN_104;	// util.scala:205:25, :206:{10,28}
  wire              dis_ld_val_1 =
    io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_ldq
    & ~io_core_dis_uops_1_bits_exception;	// lsu.scala:301:{85,88}
  wire              dis_st_val_1 =
    io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_stq
    & ~io_core_dis_uops_1_bits_exception;	// lsu.scala:301:88, :302:85
  wire [4:0]        _GEN_106 = dis_ld_val_1 ? _GEN_103 : _GEN_100;	// lsu.scala:301:85, :333:21, util.scala:206:10
  wire [4:0]        _GEN_107 = dis_st_val_1 ? _GEN_105 : _GEN_101;	// lsu.scala:302:85, :338:21, util.scala:206:10
  wire              wrap_8 = _GEN_106 == 5'h17;	// lsu.scala:333:21, util.scala:205:25
  wire [4:0]        _GEN_108 = _GEN_106 + 5'h1;	// lsu.scala:305:44, :333:21, util.scala:206:28
  wire              wrap_9 = _GEN_107 == 5'h17;	// lsu.scala:338:21, util.scala:205:25
  wire [4:0]        _GEN_109 = _GEN_107 + 5'h1;	// lsu.scala:305:44, :338:21, util.scala:206:28
  wire              dis_ld_val_2 =
    io_core_dis_uops_2_valid & io_core_dis_uops_2_bits_uses_ldq
    & ~io_core_dis_uops_2_bits_exception;	// lsu.scala:301:{85,88}
  wire              dis_st_val_2 =
    io_core_dis_uops_2_valid & io_core_dis_uops_2_bits_uses_stq
    & ~io_core_dis_uops_2_bits_exception;	// lsu.scala:301:88, :302:85
  reg               p1_block_load_mask_0;	// lsu.scala:398:35
  reg               p1_block_load_mask_1;	// lsu.scala:398:35
  reg               p1_block_load_mask_2;	// lsu.scala:398:35
  reg               p1_block_load_mask_3;	// lsu.scala:398:35
  reg               p1_block_load_mask_4;	// lsu.scala:398:35
  reg               p1_block_load_mask_5;	// lsu.scala:398:35
  reg               p1_block_load_mask_6;	// lsu.scala:398:35
  reg               p1_block_load_mask_7;	// lsu.scala:398:35
  reg               p1_block_load_mask_8;	// lsu.scala:398:35
  reg               p1_block_load_mask_9;	// lsu.scala:398:35
  reg               p1_block_load_mask_10;	// lsu.scala:398:35
  reg               p1_block_load_mask_11;	// lsu.scala:398:35
  reg               p1_block_load_mask_12;	// lsu.scala:398:35
  reg               p1_block_load_mask_13;	// lsu.scala:398:35
  reg               p1_block_load_mask_14;	// lsu.scala:398:35
  reg               p1_block_load_mask_15;	// lsu.scala:398:35
  reg               p1_block_load_mask_16;	// lsu.scala:398:35
  reg               p1_block_load_mask_17;	// lsu.scala:398:35
  reg               p1_block_load_mask_18;	// lsu.scala:398:35
  reg               p1_block_load_mask_19;	// lsu.scala:398:35
  reg               p1_block_load_mask_20;	// lsu.scala:398:35
  reg               p1_block_load_mask_21;	// lsu.scala:398:35
  reg               p1_block_load_mask_22;	// lsu.scala:398:35
  reg               p1_block_load_mask_23;	// lsu.scala:398:35
  reg               p2_block_load_mask_0;	// lsu.scala:399:35
  reg               p2_block_load_mask_1;	// lsu.scala:399:35
  reg               p2_block_load_mask_2;	// lsu.scala:399:35
  reg               p2_block_load_mask_3;	// lsu.scala:399:35
  reg               p2_block_load_mask_4;	// lsu.scala:399:35
  reg               p2_block_load_mask_5;	// lsu.scala:399:35
  reg               p2_block_load_mask_6;	// lsu.scala:399:35
  reg               p2_block_load_mask_7;	// lsu.scala:399:35
  reg               p2_block_load_mask_8;	// lsu.scala:399:35
  reg               p2_block_load_mask_9;	// lsu.scala:399:35
  reg               p2_block_load_mask_10;	// lsu.scala:399:35
  reg               p2_block_load_mask_11;	// lsu.scala:399:35
  reg               p2_block_load_mask_12;	// lsu.scala:399:35
  reg               p2_block_load_mask_13;	// lsu.scala:399:35
  reg               p2_block_load_mask_14;	// lsu.scala:399:35
  reg               p2_block_load_mask_15;	// lsu.scala:399:35
  reg               p2_block_load_mask_16;	// lsu.scala:399:35
  reg               p2_block_load_mask_17;	// lsu.scala:399:35
  reg               p2_block_load_mask_18;	// lsu.scala:399:35
  reg               p2_block_load_mask_19;	// lsu.scala:399:35
  reg               p2_block_load_mask_20;	// lsu.scala:399:35
  reg               p2_block_load_mask_21;	// lsu.scala:399:35
  reg               p2_block_load_mask_22;	// lsu.scala:399:35
  reg               p2_block_load_mask_23;	// lsu.scala:399:35
  wire [31:0][15:0] _GEN_110 =
    {{ldq_0_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask},
     {ldq_23_bits_uop_br_mask},
     {ldq_22_bits_uop_br_mask},
     {ldq_21_bits_uop_br_mask},
     {ldq_20_bits_uop_br_mask},
     {ldq_19_bits_uop_br_mask},
     {ldq_18_bits_uop_br_mask},
     {ldq_17_bits_uop_br_mask},
     {ldq_16_bits_uop_br_mask},
     {ldq_15_bits_uop_br_mask},
     {ldq_14_bits_uop_br_mask},
     {ldq_13_bits_uop_br_mask},
     {ldq_12_bits_uop_br_mask},
     {ldq_11_bits_uop_br_mask},
     {ldq_10_bits_uop_br_mask},
     {ldq_9_bits_uop_br_mask},
     {ldq_8_bits_uop_br_mask},
     {ldq_7_bits_uop_br_mask},
     {ldq_6_bits_uop_br_mask},
     {ldq_5_bits_uop_br_mask},
     {ldq_4_bits_uop_br_mask},
     {ldq_3_bits_uop_br_mask},
     {ldq_2_bits_uop_br_mask},
     {ldq_1_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask}};	// lsu.scala:210:16, :264:49
  wire [31:0][4:0]  _GEN_111 =
    {{ldq_0_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx},
     {ldq_23_bits_uop_stq_idx},
     {ldq_22_bits_uop_stq_idx},
     {ldq_21_bits_uop_stq_idx},
     {ldq_20_bits_uop_stq_idx},
     {ldq_19_bits_uop_stq_idx},
     {ldq_18_bits_uop_stq_idx},
     {ldq_17_bits_uop_stq_idx},
     {ldq_16_bits_uop_stq_idx},
     {ldq_15_bits_uop_stq_idx},
     {ldq_14_bits_uop_stq_idx},
     {ldq_13_bits_uop_stq_idx},
     {ldq_12_bits_uop_stq_idx},
     {ldq_11_bits_uop_stq_idx},
     {ldq_10_bits_uop_stq_idx},
     {ldq_9_bits_uop_stq_idx},
     {ldq_8_bits_uop_stq_idx},
     {ldq_7_bits_uop_stq_idx},
     {ldq_6_bits_uop_stq_idx},
     {ldq_5_bits_uop_stq_idx},
     {ldq_4_bits_uop_stq_idx},
     {ldq_3_bits_uop_stq_idx},
     {ldq_2_bits_uop_stq_idx},
     {ldq_1_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx}};	// lsu.scala:210:16, :264:49
  wire [31:0][1:0]  _GEN_112 =
    {{ldq_0_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size},
     {ldq_23_bits_uop_mem_size},
     {ldq_22_bits_uop_mem_size},
     {ldq_21_bits_uop_mem_size},
     {ldq_20_bits_uop_mem_size},
     {ldq_19_bits_uop_mem_size},
     {ldq_18_bits_uop_mem_size},
     {ldq_17_bits_uop_mem_size},
     {ldq_16_bits_uop_mem_size},
     {ldq_15_bits_uop_mem_size},
     {ldq_14_bits_uop_mem_size},
     {ldq_13_bits_uop_mem_size},
     {ldq_12_bits_uop_mem_size},
     {ldq_11_bits_uop_mem_size},
     {ldq_10_bits_uop_mem_size},
     {ldq_9_bits_uop_mem_size},
     {ldq_8_bits_uop_mem_size},
     {ldq_7_bits_uop_mem_size},
     {ldq_6_bits_uop_mem_size},
     {ldq_5_bits_uop_mem_size},
     {ldq_4_bits_uop_mem_size},
     {ldq_3_bits_uop_mem_size},
     {ldq_2_bits_uop_mem_size},
     {ldq_1_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size}};	// lsu.scala:210:16, :264:49
  wire [31:0]       _GEN_113 =
    {{ldq_0_bits_addr_valid},
     {ldq_0_bits_addr_valid},
     {ldq_0_bits_addr_valid},
     {ldq_0_bits_addr_valid},
     {ldq_0_bits_addr_valid},
     {ldq_0_bits_addr_valid},
     {ldq_0_bits_addr_valid},
     {ldq_0_bits_addr_valid},
     {ldq_23_bits_addr_valid},
     {ldq_22_bits_addr_valid},
     {ldq_21_bits_addr_valid},
     {ldq_20_bits_addr_valid},
     {ldq_19_bits_addr_valid},
     {ldq_18_bits_addr_valid},
     {ldq_17_bits_addr_valid},
     {ldq_16_bits_addr_valid},
     {ldq_15_bits_addr_valid},
     {ldq_14_bits_addr_valid},
     {ldq_13_bits_addr_valid},
     {ldq_12_bits_addr_valid},
     {ldq_11_bits_addr_valid},
     {ldq_10_bits_addr_valid},
     {ldq_9_bits_addr_valid},
     {ldq_8_bits_addr_valid},
     {ldq_7_bits_addr_valid},
     {ldq_6_bits_addr_valid},
     {ldq_5_bits_addr_valid},
     {ldq_4_bits_addr_valid},
     {ldq_3_bits_addr_valid},
     {ldq_2_bits_addr_valid},
     {ldq_1_bits_addr_valid},
     {ldq_0_bits_addr_valid}};	// lsu.scala:210:16, :264:49
  wire [31:0]       _GEN_114 =
    {{ldq_0_bits_executed},
     {ldq_0_bits_executed},
     {ldq_0_bits_executed},
     {ldq_0_bits_executed},
     {ldq_0_bits_executed},
     {ldq_0_bits_executed},
     {ldq_0_bits_executed},
     {ldq_0_bits_executed},
     {ldq_23_bits_executed},
     {ldq_22_bits_executed},
     {ldq_21_bits_executed},
     {ldq_20_bits_executed},
     {ldq_19_bits_executed},
     {ldq_18_bits_executed},
     {ldq_17_bits_executed},
     {ldq_16_bits_executed},
     {ldq_15_bits_executed},
     {ldq_14_bits_executed},
     {ldq_13_bits_executed},
     {ldq_12_bits_executed},
     {ldq_11_bits_executed},
     {ldq_10_bits_executed},
     {ldq_9_bits_executed},
     {ldq_8_bits_executed},
     {ldq_7_bits_executed},
     {ldq_6_bits_executed},
     {ldq_5_bits_executed},
     {ldq_4_bits_executed},
     {ldq_3_bits_executed},
     {ldq_2_bits_executed},
     {ldq_1_bits_executed},
     {ldq_0_bits_executed}};	// lsu.scala:210:16, :264:49
  wire [31:0][23:0] _GEN_115 =
    {{ldq_0_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask},
     {ldq_23_bits_st_dep_mask},
     {ldq_22_bits_st_dep_mask},
     {ldq_21_bits_st_dep_mask},
     {ldq_20_bits_st_dep_mask},
     {ldq_19_bits_st_dep_mask},
     {ldq_18_bits_st_dep_mask},
     {ldq_17_bits_st_dep_mask},
     {ldq_16_bits_st_dep_mask},
     {ldq_15_bits_st_dep_mask},
     {ldq_14_bits_st_dep_mask},
     {ldq_13_bits_st_dep_mask},
     {ldq_12_bits_st_dep_mask},
     {ldq_11_bits_st_dep_mask},
     {ldq_10_bits_st_dep_mask},
     {ldq_9_bits_st_dep_mask},
     {ldq_8_bits_st_dep_mask},
     {ldq_7_bits_st_dep_mask},
     {ldq_6_bits_st_dep_mask},
     {ldq_5_bits_st_dep_mask},
     {ldq_4_bits_st_dep_mask},
     {ldq_3_bits_st_dep_mask},
     {ldq_2_bits_st_dep_mask},
     {ldq_1_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask}};	// lsu.scala:210:16, :264:49
  reg  [4:0]        ldq_retry_idx;	// lsu.scala:415:30
  reg  [4:0]        stq_retry_idx;	// lsu.scala:422:30
  reg  [4:0]        ldq_wakeup_idx;	// lsu.scala:430:31
  wire              can_fire_load_incoming_0 =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_ctrl_is_load;	// lsu.scala:441:63
  wire              _can_fire_sta_incoming_T =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_ctrl_is_sta;	// lsu.scala:444:63
  wire [31:0][6:0]  _GEN_116 =
    {{ldq_0_bits_uop_uopc},
     {ldq_0_bits_uop_uopc},
     {ldq_0_bits_uop_uopc},
     {ldq_0_bits_uop_uopc},
     {ldq_0_bits_uop_uopc},
     {ldq_0_bits_uop_uopc},
     {ldq_0_bits_uop_uopc},
     {ldq_0_bits_uop_uopc},
     {ldq_23_bits_uop_uopc},
     {ldq_22_bits_uop_uopc},
     {ldq_21_bits_uop_uopc},
     {ldq_20_bits_uop_uopc},
     {ldq_19_bits_uop_uopc},
     {ldq_18_bits_uop_uopc},
     {ldq_17_bits_uop_uopc},
     {ldq_16_bits_uop_uopc},
     {ldq_15_bits_uop_uopc},
     {ldq_14_bits_uop_uopc},
     {ldq_13_bits_uop_uopc},
     {ldq_12_bits_uop_uopc},
     {ldq_11_bits_uop_uopc},
     {ldq_10_bits_uop_uopc},
     {ldq_9_bits_uop_uopc},
     {ldq_8_bits_uop_uopc},
     {ldq_7_bits_uop_uopc},
     {ldq_6_bits_uop_uopc},
     {ldq_5_bits_uop_uopc},
     {ldq_4_bits_uop_uopc},
     {ldq_3_bits_uop_uopc},
     {ldq_2_bits_uop_uopc},
     {ldq_1_bits_uop_uopc},
     {ldq_0_bits_uop_uopc}};	// lsu.scala:210:16, :465:79
  wire [31:0][31:0] _GEN_117 =
    {{ldq_0_bits_uop_inst},
     {ldq_0_bits_uop_inst},
     {ldq_0_bits_uop_inst},
     {ldq_0_bits_uop_inst},
     {ldq_0_bits_uop_inst},
     {ldq_0_bits_uop_inst},
     {ldq_0_bits_uop_inst},
     {ldq_0_bits_uop_inst},
     {ldq_23_bits_uop_inst},
     {ldq_22_bits_uop_inst},
     {ldq_21_bits_uop_inst},
     {ldq_20_bits_uop_inst},
     {ldq_19_bits_uop_inst},
     {ldq_18_bits_uop_inst},
     {ldq_17_bits_uop_inst},
     {ldq_16_bits_uop_inst},
     {ldq_15_bits_uop_inst},
     {ldq_14_bits_uop_inst},
     {ldq_13_bits_uop_inst},
     {ldq_12_bits_uop_inst},
     {ldq_11_bits_uop_inst},
     {ldq_10_bits_uop_inst},
     {ldq_9_bits_uop_inst},
     {ldq_8_bits_uop_inst},
     {ldq_7_bits_uop_inst},
     {ldq_6_bits_uop_inst},
     {ldq_5_bits_uop_inst},
     {ldq_4_bits_uop_inst},
     {ldq_3_bits_uop_inst},
     {ldq_2_bits_uop_inst},
     {ldq_1_bits_uop_inst},
     {ldq_0_bits_uop_inst}};	// lsu.scala:210:16, :465:79
  wire [31:0][31:0] _GEN_118 =
    {{ldq_0_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst},
     {ldq_23_bits_uop_debug_inst},
     {ldq_22_bits_uop_debug_inst},
     {ldq_21_bits_uop_debug_inst},
     {ldq_20_bits_uop_debug_inst},
     {ldq_19_bits_uop_debug_inst},
     {ldq_18_bits_uop_debug_inst},
     {ldq_17_bits_uop_debug_inst},
     {ldq_16_bits_uop_debug_inst},
     {ldq_15_bits_uop_debug_inst},
     {ldq_14_bits_uop_debug_inst},
     {ldq_13_bits_uop_debug_inst},
     {ldq_12_bits_uop_debug_inst},
     {ldq_11_bits_uop_debug_inst},
     {ldq_10_bits_uop_debug_inst},
     {ldq_9_bits_uop_debug_inst},
     {ldq_8_bits_uop_debug_inst},
     {ldq_7_bits_uop_debug_inst},
     {ldq_6_bits_uop_debug_inst},
     {ldq_5_bits_uop_debug_inst},
     {ldq_4_bits_uop_debug_inst},
     {ldq_3_bits_uop_debug_inst},
     {ldq_2_bits_uop_debug_inst},
     {ldq_1_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_119 =
    {{ldq_0_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc},
     {ldq_23_bits_uop_is_rvc},
     {ldq_22_bits_uop_is_rvc},
     {ldq_21_bits_uop_is_rvc},
     {ldq_20_bits_uop_is_rvc},
     {ldq_19_bits_uop_is_rvc},
     {ldq_18_bits_uop_is_rvc},
     {ldq_17_bits_uop_is_rvc},
     {ldq_16_bits_uop_is_rvc},
     {ldq_15_bits_uop_is_rvc},
     {ldq_14_bits_uop_is_rvc},
     {ldq_13_bits_uop_is_rvc},
     {ldq_12_bits_uop_is_rvc},
     {ldq_11_bits_uop_is_rvc},
     {ldq_10_bits_uop_is_rvc},
     {ldq_9_bits_uop_is_rvc},
     {ldq_8_bits_uop_is_rvc},
     {ldq_7_bits_uop_is_rvc},
     {ldq_6_bits_uop_is_rvc},
     {ldq_5_bits_uop_is_rvc},
     {ldq_4_bits_uop_is_rvc},
     {ldq_3_bits_uop_is_rvc},
     {ldq_2_bits_uop_is_rvc},
     {ldq_1_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc}};	// lsu.scala:210:16, :465:79
  wire [31:0][39:0] _GEN_120 =
    {{ldq_0_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc},
     {ldq_23_bits_uop_debug_pc},
     {ldq_22_bits_uop_debug_pc},
     {ldq_21_bits_uop_debug_pc},
     {ldq_20_bits_uop_debug_pc},
     {ldq_19_bits_uop_debug_pc},
     {ldq_18_bits_uop_debug_pc},
     {ldq_17_bits_uop_debug_pc},
     {ldq_16_bits_uop_debug_pc},
     {ldq_15_bits_uop_debug_pc},
     {ldq_14_bits_uop_debug_pc},
     {ldq_13_bits_uop_debug_pc},
     {ldq_12_bits_uop_debug_pc},
     {ldq_11_bits_uop_debug_pc},
     {ldq_10_bits_uop_debug_pc},
     {ldq_9_bits_uop_debug_pc},
     {ldq_8_bits_uop_debug_pc},
     {ldq_7_bits_uop_debug_pc},
     {ldq_6_bits_uop_debug_pc},
     {ldq_5_bits_uop_debug_pc},
     {ldq_4_bits_uop_debug_pc},
     {ldq_3_bits_uop_debug_pc},
     {ldq_2_bits_uop_debug_pc},
     {ldq_1_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc}};	// lsu.scala:210:16, :465:79
  wire [31:0][2:0]  _GEN_121 =
    {{ldq_0_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type},
     {ldq_23_bits_uop_iq_type},
     {ldq_22_bits_uop_iq_type},
     {ldq_21_bits_uop_iq_type},
     {ldq_20_bits_uop_iq_type},
     {ldq_19_bits_uop_iq_type},
     {ldq_18_bits_uop_iq_type},
     {ldq_17_bits_uop_iq_type},
     {ldq_16_bits_uop_iq_type},
     {ldq_15_bits_uop_iq_type},
     {ldq_14_bits_uop_iq_type},
     {ldq_13_bits_uop_iq_type},
     {ldq_12_bits_uop_iq_type},
     {ldq_11_bits_uop_iq_type},
     {ldq_10_bits_uop_iq_type},
     {ldq_9_bits_uop_iq_type},
     {ldq_8_bits_uop_iq_type},
     {ldq_7_bits_uop_iq_type},
     {ldq_6_bits_uop_iq_type},
     {ldq_5_bits_uop_iq_type},
     {ldq_4_bits_uop_iq_type},
     {ldq_3_bits_uop_iq_type},
     {ldq_2_bits_uop_iq_type},
     {ldq_1_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type}};	// lsu.scala:210:16, :465:79
  wire [31:0][9:0]  _GEN_122 =
    {{ldq_0_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code},
     {ldq_23_bits_uop_fu_code},
     {ldq_22_bits_uop_fu_code},
     {ldq_21_bits_uop_fu_code},
     {ldq_20_bits_uop_fu_code},
     {ldq_19_bits_uop_fu_code},
     {ldq_18_bits_uop_fu_code},
     {ldq_17_bits_uop_fu_code},
     {ldq_16_bits_uop_fu_code},
     {ldq_15_bits_uop_fu_code},
     {ldq_14_bits_uop_fu_code},
     {ldq_13_bits_uop_fu_code},
     {ldq_12_bits_uop_fu_code},
     {ldq_11_bits_uop_fu_code},
     {ldq_10_bits_uop_fu_code},
     {ldq_9_bits_uop_fu_code},
     {ldq_8_bits_uop_fu_code},
     {ldq_7_bits_uop_fu_code},
     {ldq_6_bits_uop_fu_code},
     {ldq_5_bits_uop_fu_code},
     {ldq_4_bits_uop_fu_code},
     {ldq_3_bits_uop_fu_code},
     {ldq_2_bits_uop_fu_code},
     {ldq_1_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code}};	// lsu.scala:210:16, :465:79
  wire [31:0][3:0]  _GEN_123 =
    {{ldq_0_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type},
     {ldq_23_bits_uop_ctrl_br_type},
     {ldq_22_bits_uop_ctrl_br_type},
     {ldq_21_bits_uop_ctrl_br_type},
     {ldq_20_bits_uop_ctrl_br_type},
     {ldq_19_bits_uop_ctrl_br_type},
     {ldq_18_bits_uop_ctrl_br_type},
     {ldq_17_bits_uop_ctrl_br_type},
     {ldq_16_bits_uop_ctrl_br_type},
     {ldq_15_bits_uop_ctrl_br_type},
     {ldq_14_bits_uop_ctrl_br_type},
     {ldq_13_bits_uop_ctrl_br_type},
     {ldq_12_bits_uop_ctrl_br_type},
     {ldq_11_bits_uop_ctrl_br_type},
     {ldq_10_bits_uop_ctrl_br_type},
     {ldq_9_bits_uop_ctrl_br_type},
     {ldq_8_bits_uop_ctrl_br_type},
     {ldq_7_bits_uop_ctrl_br_type},
     {ldq_6_bits_uop_ctrl_br_type},
     {ldq_5_bits_uop_ctrl_br_type},
     {ldq_4_bits_uop_ctrl_br_type},
     {ldq_3_bits_uop_ctrl_br_type},
     {ldq_2_bits_uop_ctrl_br_type},
     {ldq_1_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type}};	// lsu.scala:210:16, :465:79
  wire [31:0][1:0]  _GEN_124 =
    {{ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel},
     {ldq_23_bits_uop_ctrl_op1_sel},
     {ldq_22_bits_uop_ctrl_op1_sel},
     {ldq_21_bits_uop_ctrl_op1_sel},
     {ldq_20_bits_uop_ctrl_op1_sel},
     {ldq_19_bits_uop_ctrl_op1_sel},
     {ldq_18_bits_uop_ctrl_op1_sel},
     {ldq_17_bits_uop_ctrl_op1_sel},
     {ldq_16_bits_uop_ctrl_op1_sel},
     {ldq_15_bits_uop_ctrl_op1_sel},
     {ldq_14_bits_uop_ctrl_op1_sel},
     {ldq_13_bits_uop_ctrl_op1_sel},
     {ldq_12_bits_uop_ctrl_op1_sel},
     {ldq_11_bits_uop_ctrl_op1_sel},
     {ldq_10_bits_uop_ctrl_op1_sel},
     {ldq_9_bits_uop_ctrl_op1_sel},
     {ldq_8_bits_uop_ctrl_op1_sel},
     {ldq_7_bits_uop_ctrl_op1_sel},
     {ldq_6_bits_uop_ctrl_op1_sel},
     {ldq_5_bits_uop_ctrl_op1_sel},
     {ldq_4_bits_uop_ctrl_op1_sel},
     {ldq_3_bits_uop_ctrl_op1_sel},
     {ldq_2_bits_uop_ctrl_op1_sel},
     {ldq_1_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel}};	// lsu.scala:210:16, :465:79
  wire [31:0][2:0]  _GEN_125 =
    {{ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel},
     {ldq_23_bits_uop_ctrl_op2_sel},
     {ldq_22_bits_uop_ctrl_op2_sel},
     {ldq_21_bits_uop_ctrl_op2_sel},
     {ldq_20_bits_uop_ctrl_op2_sel},
     {ldq_19_bits_uop_ctrl_op2_sel},
     {ldq_18_bits_uop_ctrl_op2_sel},
     {ldq_17_bits_uop_ctrl_op2_sel},
     {ldq_16_bits_uop_ctrl_op2_sel},
     {ldq_15_bits_uop_ctrl_op2_sel},
     {ldq_14_bits_uop_ctrl_op2_sel},
     {ldq_13_bits_uop_ctrl_op2_sel},
     {ldq_12_bits_uop_ctrl_op2_sel},
     {ldq_11_bits_uop_ctrl_op2_sel},
     {ldq_10_bits_uop_ctrl_op2_sel},
     {ldq_9_bits_uop_ctrl_op2_sel},
     {ldq_8_bits_uop_ctrl_op2_sel},
     {ldq_7_bits_uop_ctrl_op2_sel},
     {ldq_6_bits_uop_ctrl_op2_sel},
     {ldq_5_bits_uop_ctrl_op2_sel},
     {ldq_4_bits_uop_ctrl_op2_sel},
     {ldq_3_bits_uop_ctrl_op2_sel},
     {ldq_2_bits_uop_ctrl_op2_sel},
     {ldq_1_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel}};	// lsu.scala:210:16, :465:79
  wire [31:0][2:0]  _GEN_126 =
    {{ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel},
     {ldq_23_bits_uop_ctrl_imm_sel},
     {ldq_22_bits_uop_ctrl_imm_sel},
     {ldq_21_bits_uop_ctrl_imm_sel},
     {ldq_20_bits_uop_ctrl_imm_sel},
     {ldq_19_bits_uop_ctrl_imm_sel},
     {ldq_18_bits_uop_ctrl_imm_sel},
     {ldq_17_bits_uop_ctrl_imm_sel},
     {ldq_16_bits_uop_ctrl_imm_sel},
     {ldq_15_bits_uop_ctrl_imm_sel},
     {ldq_14_bits_uop_ctrl_imm_sel},
     {ldq_13_bits_uop_ctrl_imm_sel},
     {ldq_12_bits_uop_ctrl_imm_sel},
     {ldq_11_bits_uop_ctrl_imm_sel},
     {ldq_10_bits_uop_ctrl_imm_sel},
     {ldq_9_bits_uop_ctrl_imm_sel},
     {ldq_8_bits_uop_ctrl_imm_sel},
     {ldq_7_bits_uop_ctrl_imm_sel},
     {ldq_6_bits_uop_ctrl_imm_sel},
     {ldq_5_bits_uop_ctrl_imm_sel},
     {ldq_4_bits_uop_ctrl_imm_sel},
     {ldq_3_bits_uop_ctrl_imm_sel},
     {ldq_2_bits_uop_ctrl_imm_sel},
     {ldq_1_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel}};	// lsu.scala:210:16, :465:79
  wire [31:0][3:0]  _GEN_127 =
    {{ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn},
     {ldq_23_bits_uop_ctrl_op_fcn},
     {ldq_22_bits_uop_ctrl_op_fcn},
     {ldq_21_bits_uop_ctrl_op_fcn},
     {ldq_20_bits_uop_ctrl_op_fcn},
     {ldq_19_bits_uop_ctrl_op_fcn},
     {ldq_18_bits_uop_ctrl_op_fcn},
     {ldq_17_bits_uop_ctrl_op_fcn},
     {ldq_16_bits_uop_ctrl_op_fcn},
     {ldq_15_bits_uop_ctrl_op_fcn},
     {ldq_14_bits_uop_ctrl_op_fcn},
     {ldq_13_bits_uop_ctrl_op_fcn},
     {ldq_12_bits_uop_ctrl_op_fcn},
     {ldq_11_bits_uop_ctrl_op_fcn},
     {ldq_10_bits_uop_ctrl_op_fcn},
     {ldq_9_bits_uop_ctrl_op_fcn},
     {ldq_8_bits_uop_ctrl_op_fcn},
     {ldq_7_bits_uop_ctrl_op_fcn},
     {ldq_6_bits_uop_ctrl_op_fcn},
     {ldq_5_bits_uop_ctrl_op_fcn},
     {ldq_4_bits_uop_ctrl_op_fcn},
     {ldq_3_bits_uop_ctrl_op_fcn},
     {ldq_2_bits_uop_ctrl_op_fcn},
     {ldq_1_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_128 =
    {{ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw},
     {ldq_23_bits_uop_ctrl_fcn_dw},
     {ldq_22_bits_uop_ctrl_fcn_dw},
     {ldq_21_bits_uop_ctrl_fcn_dw},
     {ldq_20_bits_uop_ctrl_fcn_dw},
     {ldq_19_bits_uop_ctrl_fcn_dw},
     {ldq_18_bits_uop_ctrl_fcn_dw},
     {ldq_17_bits_uop_ctrl_fcn_dw},
     {ldq_16_bits_uop_ctrl_fcn_dw},
     {ldq_15_bits_uop_ctrl_fcn_dw},
     {ldq_14_bits_uop_ctrl_fcn_dw},
     {ldq_13_bits_uop_ctrl_fcn_dw},
     {ldq_12_bits_uop_ctrl_fcn_dw},
     {ldq_11_bits_uop_ctrl_fcn_dw},
     {ldq_10_bits_uop_ctrl_fcn_dw},
     {ldq_9_bits_uop_ctrl_fcn_dw},
     {ldq_8_bits_uop_ctrl_fcn_dw},
     {ldq_7_bits_uop_ctrl_fcn_dw},
     {ldq_6_bits_uop_ctrl_fcn_dw},
     {ldq_5_bits_uop_ctrl_fcn_dw},
     {ldq_4_bits_uop_ctrl_fcn_dw},
     {ldq_3_bits_uop_ctrl_fcn_dw},
     {ldq_2_bits_uop_ctrl_fcn_dw},
     {ldq_1_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw}};	// lsu.scala:210:16, :465:79
  wire [31:0][2:0]  _GEN_129 =
    {{ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd},
     {ldq_23_bits_uop_ctrl_csr_cmd},
     {ldq_22_bits_uop_ctrl_csr_cmd},
     {ldq_21_bits_uop_ctrl_csr_cmd},
     {ldq_20_bits_uop_ctrl_csr_cmd},
     {ldq_19_bits_uop_ctrl_csr_cmd},
     {ldq_18_bits_uop_ctrl_csr_cmd},
     {ldq_17_bits_uop_ctrl_csr_cmd},
     {ldq_16_bits_uop_ctrl_csr_cmd},
     {ldq_15_bits_uop_ctrl_csr_cmd},
     {ldq_14_bits_uop_ctrl_csr_cmd},
     {ldq_13_bits_uop_ctrl_csr_cmd},
     {ldq_12_bits_uop_ctrl_csr_cmd},
     {ldq_11_bits_uop_ctrl_csr_cmd},
     {ldq_10_bits_uop_ctrl_csr_cmd},
     {ldq_9_bits_uop_ctrl_csr_cmd},
     {ldq_8_bits_uop_ctrl_csr_cmd},
     {ldq_7_bits_uop_ctrl_csr_cmd},
     {ldq_6_bits_uop_ctrl_csr_cmd},
     {ldq_5_bits_uop_ctrl_csr_cmd},
     {ldq_4_bits_uop_ctrl_csr_cmd},
     {ldq_3_bits_uop_ctrl_csr_cmd},
     {ldq_2_bits_uop_ctrl_csr_cmd},
     {ldq_1_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_130 =
    {{ldq_0_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load},
     {ldq_23_bits_uop_ctrl_is_load},
     {ldq_22_bits_uop_ctrl_is_load},
     {ldq_21_bits_uop_ctrl_is_load},
     {ldq_20_bits_uop_ctrl_is_load},
     {ldq_19_bits_uop_ctrl_is_load},
     {ldq_18_bits_uop_ctrl_is_load},
     {ldq_17_bits_uop_ctrl_is_load},
     {ldq_16_bits_uop_ctrl_is_load},
     {ldq_15_bits_uop_ctrl_is_load},
     {ldq_14_bits_uop_ctrl_is_load},
     {ldq_13_bits_uop_ctrl_is_load},
     {ldq_12_bits_uop_ctrl_is_load},
     {ldq_11_bits_uop_ctrl_is_load},
     {ldq_10_bits_uop_ctrl_is_load},
     {ldq_9_bits_uop_ctrl_is_load},
     {ldq_8_bits_uop_ctrl_is_load},
     {ldq_7_bits_uop_ctrl_is_load},
     {ldq_6_bits_uop_ctrl_is_load},
     {ldq_5_bits_uop_ctrl_is_load},
     {ldq_4_bits_uop_ctrl_is_load},
     {ldq_3_bits_uop_ctrl_is_load},
     {ldq_2_bits_uop_ctrl_is_load},
     {ldq_1_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_131 =
    {{ldq_0_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta},
     {ldq_23_bits_uop_ctrl_is_sta},
     {ldq_22_bits_uop_ctrl_is_sta},
     {ldq_21_bits_uop_ctrl_is_sta},
     {ldq_20_bits_uop_ctrl_is_sta},
     {ldq_19_bits_uop_ctrl_is_sta},
     {ldq_18_bits_uop_ctrl_is_sta},
     {ldq_17_bits_uop_ctrl_is_sta},
     {ldq_16_bits_uop_ctrl_is_sta},
     {ldq_15_bits_uop_ctrl_is_sta},
     {ldq_14_bits_uop_ctrl_is_sta},
     {ldq_13_bits_uop_ctrl_is_sta},
     {ldq_12_bits_uop_ctrl_is_sta},
     {ldq_11_bits_uop_ctrl_is_sta},
     {ldq_10_bits_uop_ctrl_is_sta},
     {ldq_9_bits_uop_ctrl_is_sta},
     {ldq_8_bits_uop_ctrl_is_sta},
     {ldq_7_bits_uop_ctrl_is_sta},
     {ldq_6_bits_uop_ctrl_is_sta},
     {ldq_5_bits_uop_ctrl_is_sta},
     {ldq_4_bits_uop_ctrl_is_sta},
     {ldq_3_bits_uop_ctrl_is_sta},
     {ldq_2_bits_uop_ctrl_is_sta},
     {ldq_1_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_132 =
    {{ldq_0_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std},
     {ldq_23_bits_uop_ctrl_is_std},
     {ldq_22_bits_uop_ctrl_is_std},
     {ldq_21_bits_uop_ctrl_is_std},
     {ldq_20_bits_uop_ctrl_is_std},
     {ldq_19_bits_uop_ctrl_is_std},
     {ldq_18_bits_uop_ctrl_is_std},
     {ldq_17_bits_uop_ctrl_is_std},
     {ldq_16_bits_uop_ctrl_is_std},
     {ldq_15_bits_uop_ctrl_is_std},
     {ldq_14_bits_uop_ctrl_is_std},
     {ldq_13_bits_uop_ctrl_is_std},
     {ldq_12_bits_uop_ctrl_is_std},
     {ldq_11_bits_uop_ctrl_is_std},
     {ldq_10_bits_uop_ctrl_is_std},
     {ldq_9_bits_uop_ctrl_is_std},
     {ldq_8_bits_uop_ctrl_is_std},
     {ldq_7_bits_uop_ctrl_is_std},
     {ldq_6_bits_uop_ctrl_is_std},
     {ldq_5_bits_uop_ctrl_is_std},
     {ldq_4_bits_uop_ctrl_is_std},
     {ldq_3_bits_uop_ctrl_is_std},
     {ldq_2_bits_uop_ctrl_is_std},
     {ldq_1_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std}};	// lsu.scala:210:16, :465:79
  wire [31:0][1:0]  _GEN_133 =
    {{ldq_0_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state},
     {ldq_23_bits_uop_iw_state},
     {ldq_22_bits_uop_iw_state},
     {ldq_21_bits_uop_iw_state},
     {ldq_20_bits_uop_iw_state},
     {ldq_19_bits_uop_iw_state},
     {ldq_18_bits_uop_iw_state},
     {ldq_17_bits_uop_iw_state},
     {ldq_16_bits_uop_iw_state},
     {ldq_15_bits_uop_iw_state},
     {ldq_14_bits_uop_iw_state},
     {ldq_13_bits_uop_iw_state},
     {ldq_12_bits_uop_iw_state},
     {ldq_11_bits_uop_iw_state},
     {ldq_10_bits_uop_iw_state},
     {ldq_9_bits_uop_iw_state},
     {ldq_8_bits_uop_iw_state},
     {ldq_7_bits_uop_iw_state},
     {ldq_6_bits_uop_iw_state},
     {ldq_5_bits_uop_iw_state},
     {ldq_4_bits_uop_iw_state},
     {ldq_3_bits_uop_iw_state},
     {ldq_2_bits_uop_iw_state},
     {ldq_1_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_134 =
    {{ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned},
     {ldq_23_bits_uop_iw_p1_poisoned},
     {ldq_22_bits_uop_iw_p1_poisoned},
     {ldq_21_bits_uop_iw_p1_poisoned},
     {ldq_20_bits_uop_iw_p1_poisoned},
     {ldq_19_bits_uop_iw_p1_poisoned},
     {ldq_18_bits_uop_iw_p1_poisoned},
     {ldq_17_bits_uop_iw_p1_poisoned},
     {ldq_16_bits_uop_iw_p1_poisoned},
     {ldq_15_bits_uop_iw_p1_poisoned},
     {ldq_14_bits_uop_iw_p1_poisoned},
     {ldq_13_bits_uop_iw_p1_poisoned},
     {ldq_12_bits_uop_iw_p1_poisoned},
     {ldq_11_bits_uop_iw_p1_poisoned},
     {ldq_10_bits_uop_iw_p1_poisoned},
     {ldq_9_bits_uop_iw_p1_poisoned},
     {ldq_8_bits_uop_iw_p1_poisoned},
     {ldq_7_bits_uop_iw_p1_poisoned},
     {ldq_6_bits_uop_iw_p1_poisoned},
     {ldq_5_bits_uop_iw_p1_poisoned},
     {ldq_4_bits_uop_iw_p1_poisoned},
     {ldq_3_bits_uop_iw_p1_poisoned},
     {ldq_2_bits_uop_iw_p1_poisoned},
     {ldq_1_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_135 =
    {{ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned},
     {ldq_23_bits_uop_iw_p2_poisoned},
     {ldq_22_bits_uop_iw_p2_poisoned},
     {ldq_21_bits_uop_iw_p2_poisoned},
     {ldq_20_bits_uop_iw_p2_poisoned},
     {ldq_19_bits_uop_iw_p2_poisoned},
     {ldq_18_bits_uop_iw_p2_poisoned},
     {ldq_17_bits_uop_iw_p2_poisoned},
     {ldq_16_bits_uop_iw_p2_poisoned},
     {ldq_15_bits_uop_iw_p2_poisoned},
     {ldq_14_bits_uop_iw_p2_poisoned},
     {ldq_13_bits_uop_iw_p2_poisoned},
     {ldq_12_bits_uop_iw_p2_poisoned},
     {ldq_11_bits_uop_iw_p2_poisoned},
     {ldq_10_bits_uop_iw_p2_poisoned},
     {ldq_9_bits_uop_iw_p2_poisoned},
     {ldq_8_bits_uop_iw_p2_poisoned},
     {ldq_7_bits_uop_iw_p2_poisoned},
     {ldq_6_bits_uop_iw_p2_poisoned},
     {ldq_5_bits_uop_iw_p2_poisoned},
     {ldq_4_bits_uop_iw_p2_poisoned},
     {ldq_3_bits_uop_iw_p2_poisoned},
     {ldq_2_bits_uop_iw_p2_poisoned},
     {ldq_1_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_136 =
    {{ldq_0_bits_uop_is_br},
     {ldq_0_bits_uop_is_br},
     {ldq_0_bits_uop_is_br},
     {ldq_0_bits_uop_is_br},
     {ldq_0_bits_uop_is_br},
     {ldq_0_bits_uop_is_br},
     {ldq_0_bits_uop_is_br},
     {ldq_0_bits_uop_is_br},
     {ldq_23_bits_uop_is_br},
     {ldq_22_bits_uop_is_br},
     {ldq_21_bits_uop_is_br},
     {ldq_20_bits_uop_is_br},
     {ldq_19_bits_uop_is_br},
     {ldq_18_bits_uop_is_br},
     {ldq_17_bits_uop_is_br},
     {ldq_16_bits_uop_is_br},
     {ldq_15_bits_uop_is_br},
     {ldq_14_bits_uop_is_br},
     {ldq_13_bits_uop_is_br},
     {ldq_12_bits_uop_is_br},
     {ldq_11_bits_uop_is_br},
     {ldq_10_bits_uop_is_br},
     {ldq_9_bits_uop_is_br},
     {ldq_8_bits_uop_is_br},
     {ldq_7_bits_uop_is_br},
     {ldq_6_bits_uop_is_br},
     {ldq_5_bits_uop_is_br},
     {ldq_4_bits_uop_is_br},
     {ldq_3_bits_uop_is_br},
     {ldq_2_bits_uop_is_br},
     {ldq_1_bits_uop_is_br},
     {ldq_0_bits_uop_is_br}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_137 =
    {{ldq_0_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr},
     {ldq_23_bits_uop_is_jalr},
     {ldq_22_bits_uop_is_jalr},
     {ldq_21_bits_uop_is_jalr},
     {ldq_20_bits_uop_is_jalr},
     {ldq_19_bits_uop_is_jalr},
     {ldq_18_bits_uop_is_jalr},
     {ldq_17_bits_uop_is_jalr},
     {ldq_16_bits_uop_is_jalr},
     {ldq_15_bits_uop_is_jalr},
     {ldq_14_bits_uop_is_jalr},
     {ldq_13_bits_uop_is_jalr},
     {ldq_12_bits_uop_is_jalr},
     {ldq_11_bits_uop_is_jalr},
     {ldq_10_bits_uop_is_jalr},
     {ldq_9_bits_uop_is_jalr},
     {ldq_8_bits_uop_is_jalr},
     {ldq_7_bits_uop_is_jalr},
     {ldq_6_bits_uop_is_jalr},
     {ldq_5_bits_uop_is_jalr},
     {ldq_4_bits_uop_is_jalr},
     {ldq_3_bits_uop_is_jalr},
     {ldq_2_bits_uop_is_jalr},
     {ldq_1_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_138 =
    {{ldq_0_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal},
     {ldq_23_bits_uop_is_jal},
     {ldq_22_bits_uop_is_jal},
     {ldq_21_bits_uop_is_jal},
     {ldq_20_bits_uop_is_jal},
     {ldq_19_bits_uop_is_jal},
     {ldq_18_bits_uop_is_jal},
     {ldq_17_bits_uop_is_jal},
     {ldq_16_bits_uop_is_jal},
     {ldq_15_bits_uop_is_jal},
     {ldq_14_bits_uop_is_jal},
     {ldq_13_bits_uop_is_jal},
     {ldq_12_bits_uop_is_jal},
     {ldq_11_bits_uop_is_jal},
     {ldq_10_bits_uop_is_jal},
     {ldq_9_bits_uop_is_jal},
     {ldq_8_bits_uop_is_jal},
     {ldq_7_bits_uop_is_jal},
     {ldq_6_bits_uop_is_jal},
     {ldq_5_bits_uop_is_jal},
     {ldq_4_bits_uop_is_jal},
     {ldq_3_bits_uop_is_jal},
     {ldq_2_bits_uop_is_jal},
     {ldq_1_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_139 =
    {{ldq_0_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb},
     {ldq_23_bits_uop_is_sfb},
     {ldq_22_bits_uop_is_sfb},
     {ldq_21_bits_uop_is_sfb},
     {ldq_20_bits_uop_is_sfb},
     {ldq_19_bits_uop_is_sfb},
     {ldq_18_bits_uop_is_sfb},
     {ldq_17_bits_uop_is_sfb},
     {ldq_16_bits_uop_is_sfb},
     {ldq_15_bits_uop_is_sfb},
     {ldq_14_bits_uop_is_sfb},
     {ldq_13_bits_uop_is_sfb},
     {ldq_12_bits_uop_is_sfb},
     {ldq_11_bits_uop_is_sfb},
     {ldq_10_bits_uop_is_sfb},
     {ldq_9_bits_uop_is_sfb},
     {ldq_8_bits_uop_is_sfb},
     {ldq_7_bits_uop_is_sfb},
     {ldq_6_bits_uop_is_sfb},
     {ldq_5_bits_uop_is_sfb},
     {ldq_4_bits_uop_is_sfb},
     {ldq_3_bits_uop_is_sfb},
     {ldq_2_bits_uop_is_sfb},
     {ldq_1_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_140 = _GEN_110[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79
  wire [31:0][3:0]  _GEN_141 =
    {{ldq_0_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag},
     {ldq_23_bits_uop_br_tag},
     {ldq_22_bits_uop_br_tag},
     {ldq_21_bits_uop_br_tag},
     {ldq_20_bits_uop_br_tag},
     {ldq_19_bits_uop_br_tag},
     {ldq_18_bits_uop_br_tag},
     {ldq_17_bits_uop_br_tag},
     {ldq_16_bits_uop_br_tag},
     {ldq_15_bits_uop_br_tag},
     {ldq_14_bits_uop_br_tag},
     {ldq_13_bits_uop_br_tag},
     {ldq_12_bits_uop_br_tag},
     {ldq_11_bits_uop_br_tag},
     {ldq_10_bits_uop_br_tag},
     {ldq_9_bits_uop_br_tag},
     {ldq_8_bits_uop_br_tag},
     {ldq_7_bits_uop_br_tag},
     {ldq_6_bits_uop_br_tag},
     {ldq_5_bits_uop_br_tag},
     {ldq_4_bits_uop_br_tag},
     {ldq_3_bits_uop_br_tag},
     {ldq_2_bits_uop_br_tag},
     {ldq_1_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag}};	// lsu.scala:210:16, :465:79
  wire [31:0][4:0]  _GEN_142 =
    {{ldq_0_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx},
     {ldq_23_bits_uop_ftq_idx},
     {ldq_22_bits_uop_ftq_idx},
     {ldq_21_bits_uop_ftq_idx},
     {ldq_20_bits_uop_ftq_idx},
     {ldq_19_bits_uop_ftq_idx},
     {ldq_18_bits_uop_ftq_idx},
     {ldq_17_bits_uop_ftq_idx},
     {ldq_16_bits_uop_ftq_idx},
     {ldq_15_bits_uop_ftq_idx},
     {ldq_14_bits_uop_ftq_idx},
     {ldq_13_bits_uop_ftq_idx},
     {ldq_12_bits_uop_ftq_idx},
     {ldq_11_bits_uop_ftq_idx},
     {ldq_10_bits_uop_ftq_idx},
     {ldq_9_bits_uop_ftq_idx},
     {ldq_8_bits_uop_ftq_idx},
     {ldq_7_bits_uop_ftq_idx},
     {ldq_6_bits_uop_ftq_idx},
     {ldq_5_bits_uop_ftq_idx},
     {ldq_4_bits_uop_ftq_idx},
     {ldq_3_bits_uop_ftq_idx},
     {ldq_2_bits_uop_ftq_idx},
     {ldq_1_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_143 =
    {{ldq_0_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst},
     {ldq_23_bits_uop_edge_inst},
     {ldq_22_bits_uop_edge_inst},
     {ldq_21_bits_uop_edge_inst},
     {ldq_20_bits_uop_edge_inst},
     {ldq_19_bits_uop_edge_inst},
     {ldq_18_bits_uop_edge_inst},
     {ldq_17_bits_uop_edge_inst},
     {ldq_16_bits_uop_edge_inst},
     {ldq_15_bits_uop_edge_inst},
     {ldq_14_bits_uop_edge_inst},
     {ldq_13_bits_uop_edge_inst},
     {ldq_12_bits_uop_edge_inst},
     {ldq_11_bits_uop_edge_inst},
     {ldq_10_bits_uop_edge_inst},
     {ldq_9_bits_uop_edge_inst},
     {ldq_8_bits_uop_edge_inst},
     {ldq_7_bits_uop_edge_inst},
     {ldq_6_bits_uop_edge_inst},
     {ldq_5_bits_uop_edge_inst},
     {ldq_4_bits_uop_edge_inst},
     {ldq_3_bits_uop_edge_inst},
     {ldq_2_bits_uop_edge_inst},
     {ldq_1_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst}};	// lsu.scala:210:16, :465:79
  wire [31:0][5:0]  _GEN_144 =
    {{ldq_0_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob},
     {ldq_23_bits_uop_pc_lob},
     {ldq_22_bits_uop_pc_lob},
     {ldq_21_bits_uop_pc_lob},
     {ldq_20_bits_uop_pc_lob},
     {ldq_19_bits_uop_pc_lob},
     {ldq_18_bits_uop_pc_lob},
     {ldq_17_bits_uop_pc_lob},
     {ldq_16_bits_uop_pc_lob},
     {ldq_15_bits_uop_pc_lob},
     {ldq_14_bits_uop_pc_lob},
     {ldq_13_bits_uop_pc_lob},
     {ldq_12_bits_uop_pc_lob},
     {ldq_11_bits_uop_pc_lob},
     {ldq_10_bits_uop_pc_lob},
     {ldq_9_bits_uop_pc_lob},
     {ldq_8_bits_uop_pc_lob},
     {ldq_7_bits_uop_pc_lob},
     {ldq_6_bits_uop_pc_lob},
     {ldq_5_bits_uop_pc_lob},
     {ldq_4_bits_uop_pc_lob},
     {ldq_3_bits_uop_pc_lob},
     {ldq_2_bits_uop_pc_lob},
     {ldq_1_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_145 =
    {{ldq_0_bits_uop_taken},
     {ldq_0_bits_uop_taken},
     {ldq_0_bits_uop_taken},
     {ldq_0_bits_uop_taken},
     {ldq_0_bits_uop_taken},
     {ldq_0_bits_uop_taken},
     {ldq_0_bits_uop_taken},
     {ldq_0_bits_uop_taken},
     {ldq_23_bits_uop_taken},
     {ldq_22_bits_uop_taken},
     {ldq_21_bits_uop_taken},
     {ldq_20_bits_uop_taken},
     {ldq_19_bits_uop_taken},
     {ldq_18_bits_uop_taken},
     {ldq_17_bits_uop_taken},
     {ldq_16_bits_uop_taken},
     {ldq_15_bits_uop_taken},
     {ldq_14_bits_uop_taken},
     {ldq_13_bits_uop_taken},
     {ldq_12_bits_uop_taken},
     {ldq_11_bits_uop_taken},
     {ldq_10_bits_uop_taken},
     {ldq_9_bits_uop_taken},
     {ldq_8_bits_uop_taken},
     {ldq_7_bits_uop_taken},
     {ldq_6_bits_uop_taken},
     {ldq_5_bits_uop_taken},
     {ldq_4_bits_uop_taken},
     {ldq_3_bits_uop_taken},
     {ldq_2_bits_uop_taken},
     {ldq_1_bits_uop_taken},
     {ldq_0_bits_uop_taken}};	// lsu.scala:210:16, :465:79
  wire [31:0][19:0] _GEN_146 =
    {{ldq_0_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed},
     {ldq_23_bits_uop_imm_packed},
     {ldq_22_bits_uop_imm_packed},
     {ldq_21_bits_uop_imm_packed},
     {ldq_20_bits_uop_imm_packed},
     {ldq_19_bits_uop_imm_packed},
     {ldq_18_bits_uop_imm_packed},
     {ldq_17_bits_uop_imm_packed},
     {ldq_16_bits_uop_imm_packed},
     {ldq_15_bits_uop_imm_packed},
     {ldq_14_bits_uop_imm_packed},
     {ldq_13_bits_uop_imm_packed},
     {ldq_12_bits_uop_imm_packed},
     {ldq_11_bits_uop_imm_packed},
     {ldq_10_bits_uop_imm_packed},
     {ldq_9_bits_uop_imm_packed},
     {ldq_8_bits_uop_imm_packed},
     {ldq_7_bits_uop_imm_packed},
     {ldq_6_bits_uop_imm_packed},
     {ldq_5_bits_uop_imm_packed},
     {ldq_4_bits_uop_imm_packed},
     {ldq_3_bits_uop_imm_packed},
     {ldq_2_bits_uop_imm_packed},
     {ldq_1_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed}};	// lsu.scala:210:16, :465:79
  wire [31:0][11:0] _GEN_147 =
    {{ldq_0_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr},
     {ldq_23_bits_uop_csr_addr},
     {ldq_22_bits_uop_csr_addr},
     {ldq_21_bits_uop_csr_addr},
     {ldq_20_bits_uop_csr_addr},
     {ldq_19_bits_uop_csr_addr},
     {ldq_18_bits_uop_csr_addr},
     {ldq_17_bits_uop_csr_addr},
     {ldq_16_bits_uop_csr_addr},
     {ldq_15_bits_uop_csr_addr},
     {ldq_14_bits_uop_csr_addr},
     {ldq_13_bits_uop_csr_addr},
     {ldq_12_bits_uop_csr_addr},
     {ldq_11_bits_uop_csr_addr},
     {ldq_10_bits_uop_csr_addr},
     {ldq_9_bits_uop_csr_addr},
     {ldq_8_bits_uop_csr_addr},
     {ldq_7_bits_uop_csr_addr},
     {ldq_6_bits_uop_csr_addr},
     {ldq_5_bits_uop_csr_addr},
     {ldq_4_bits_uop_csr_addr},
     {ldq_3_bits_uop_csr_addr},
     {ldq_2_bits_uop_csr_addr},
     {ldq_1_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr}};	// lsu.scala:210:16, :465:79
  wire [31:0][6:0]  _GEN_148 =
    {{ldq_0_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx},
     {ldq_23_bits_uop_rob_idx},
     {ldq_22_bits_uop_rob_idx},
     {ldq_21_bits_uop_rob_idx},
     {ldq_20_bits_uop_rob_idx},
     {ldq_19_bits_uop_rob_idx},
     {ldq_18_bits_uop_rob_idx},
     {ldq_17_bits_uop_rob_idx},
     {ldq_16_bits_uop_rob_idx},
     {ldq_15_bits_uop_rob_idx},
     {ldq_14_bits_uop_rob_idx},
     {ldq_13_bits_uop_rob_idx},
     {ldq_12_bits_uop_rob_idx},
     {ldq_11_bits_uop_rob_idx},
     {ldq_10_bits_uop_rob_idx},
     {ldq_9_bits_uop_rob_idx},
     {ldq_8_bits_uop_rob_idx},
     {ldq_7_bits_uop_rob_idx},
     {ldq_6_bits_uop_rob_idx},
     {ldq_5_bits_uop_rob_idx},
     {ldq_4_bits_uop_rob_idx},
     {ldq_3_bits_uop_rob_idx},
     {ldq_2_bits_uop_rob_idx},
     {ldq_1_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx}};	// lsu.scala:210:16, :465:79
  wire [6:0]        _GEN_149 = _GEN_148[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [31:0][4:0]  _GEN_150 =
    {{ldq_0_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx},
     {ldq_23_bits_uop_ldq_idx},
     {ldq_22_bits_uop_ldq_idx},
     {ldq_21_bits_uop_ldq_idx},
     {ldq_20_bits_uop_ldq_idx},
     {ldq_19_bits_uop_ldq_idx},
     {ldq_18_bits_uop_ldq_idx},
     {ldq_17_bits_uop_ldq_idx},
     {ldq_16_bits_uop_ldq_idx},
     {ldq_15_bits_uop_ldq_idx},
     {ldq_14_bits_uop_ldq_idx},
     {ldq_13_bits_uop_ldq_idx},
     {ldq_12_bits_uop_ldq_idx},
     {ldq_11_bits_uop_ldq_idx},
     {ldq_10_bits_uop_ldq_idx},
     {ldq_9_bits_uop_ldq_idx},
     {ldq_8_bits_uop_ldq_idx},
     {ldq_7_bits_uop_ldq_idx},
     {ldq_6_bits_uop_ldq_idx},
     {ldq_5_bits_uop_ldq_idx},
     {ldq_4_bits_uop_ldq_idx},
     {ldq_3_bits_uop_ldq_idx},
     {ldq_2_bits_uop_ldq_idx},
     {ldq_1_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx}};	// lsu.scala:210:16, :465:79
  wire [4:0]        _GEN_151 = _GEN_150[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [4:0]        mem_ldq_retry_e_out_bits_uop_stq_idx = _GEN_111[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79
  wire [31:0][1:0]  _GEN_152 =
    {{ldq_0_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx},
     {ldq_23_bits_uop_rxq_idx},
     {ldq_22_bits_uop_rxq_idx},
     {ldq_21_bits_uop_rxq_idx},
     {ldq_20_bits_uop_rxq_idx},
     {ldq_19_bits_uop_rxq_idx},
     {ldq_18_bits_uop_rxq_idx},
     {ldq_17_bits_uop_rxq_idx},
     {ldq_16_bits_uop_rxq_idx},
     {ldq_15_bits_uop_rxq_idx},
     {ldq_14_bits_uop_rxq_idx},
     {ldq_13_bits_uop_rxq_idx},
     {ldq_12_bits_uop_rxq_idx},
     {ldq_11_bits_uop_rxq_idx},
     {ldq_10_bits_uop_rxq_idx},
     {ldq_9_bits_uop_rxq_idx},
     {ldq_8_bits_uop_rxq_idx},
     {ldq_7_bits_uop_rxq_idx},
     {ldq_6_bits_uop_rxq_idx},
     {ldq_5_bits_uop_rxq_idx},
     {ldq_4_bits_uop_rxq_idx},
     {ldq_3_bits_uop_rxq_idx},
     {ldq_2_bits_uop_rxq_idx},
     {ldq_1_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx}};	// lsu.scala:210:16, :465:79
  wire [31:0][6:0]  _GEN_153 =
    {{ldq_0_bits_uop_pdst},
     {ldq_0_bits_uop_pdst},
     {ldq_0_bits_uop_pdst},
     {ldq_0_bits_uop_pdst},
     {ldq_0_bits_uop_pdst},
     {ldq_0_bits_uop_pdst},
     {ldq_0_bits_uop_pdst},
     {ldq_0_bits_uop_pdst},
     {ldq_23_bits_uop_pdst},
     {ldq_22_bits_uop_pdst},
     {ldq_21_bits_uop_pdst},
     {ldq_20_bits_uop_pdst},
     {ldq_19_bits_uop_pdst},
     {ldq_18_bits_uop_pdst},
     {ldq_17_bits_uop_pdst},
     {ldq_16_bits_uop_pdst},
     {ldq_15_bits_uop_pdst},
     {ldq_14_bits_uop_pdst},
     {ldq_13_bits_uop_pdst},
     {ldq_12_bits_uop_pdst},
     {ldq_11_bits_uop_pdst},
     {ldq_10_bits_uop_pdst},
     {ldq_9_bits_uop_pdst},
     {ldq_8_bits_uop_pdst},
     {ldq_7_bits_uop_pdst},
     {ldq_6_bits_uop_pdst},
     {ldq_5_bits_uop_pdst},
     {ldq_4_bits_uop_pdst},
     {ldq_3_bits_uop_pdst},
     {ldq_2_bits_uop_pdst},
     {ldq_1_bits_uop_pdst},
     {ldq_0_bits_uop_pdst}};	// lsu.scala:210:16, :465:79
  wire [6:0]        _GEN_154 = _GEN_153[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [31:0][6:0]  _GEN_155 =
    {{ldq_0_bits_uop_prs1},
     {ldq_0_bits_uop_prs1},
     {ldq_0_bits_uop_prs1},
     {ldq_0_bits_uop_prs1},
     {ldq_0_bits_uop_prs1},
     {ldq_0_bits_uop_prs1},
     {ldq_0_bits_uop_prs1},
     {ldq_0_bits_uop_prs1},
     {ldq_23_bits_uop_prs1},
     {ldq_22_bits_uop_prs1},
     {ldq_21_bits_uop_prs1},
     {ldq_20_bits_uop_prs1},
     {ldq_19_bits_uop_prs1},
     {ldq_18_bits_uop_prs1},
     {ldq_17_bits_uop_prs1},
     {ldq_16_bits_uop_prs1},
     {ldq_15_bits_uop_prs1},
     {ldq_14_bits_uop_prs1},
     {ldq_13_bits_uop_prs1},
     {ldq_12_bits_uop_prs1},
     {ldq_11_bits_uop_prs1},
     {ldq_10_bits_uop_prs1},
     {ldq_9_bits_uop_prs1},
     {ldq_8_bits_uop_prs1},
     {ldq_7_bits_uop_prs1},
     {ldq_6_bits_uop_prs1},
     {ldq_5_bits_uop_prs1},
     {ldq_4_bits_uop_prs1},
     {ldq_3_bits_uop_prs1},
     {ldq_2_bits_uop_prs1},
     {ldq_1_bits_uop_prs1},
     {ldq_0_bits_uop_prs1}};	// lsu.scala:210:16, :465:79
  wire [31:0][6:0]  _GEN_156 =
    {{ldq_0_bits_uop_prs2},
     {ldq_0_bits_uop_prs2},
     {ldq_0_bits_uop_prs2},
     {ldq_0_bits_uop_prs2},
     {ldq_0_bits_uop_prs2},
     {ldq_0_bits_uop_prs2},
     {ldq_0_bits_uop_prs2},
     {ldq_0_bits_uop_prs2},
     {ldq_23_bits_uop_prs2},
     {ldq_22_bits_uop_prs2},
     {ldq_21_bits_uop_prs2},
     {ldq_20_bits_uop_prs2},
     {ldq_19_bits_uop_prs2},
     {ldq_18_bits_uop_prs2},
     {ldq_17_bits_uop_prs2},
     {ldq_16_bits_uop_prs2},
     {ldq_15_bits_uop_prs2},
     {ldq_14_bits_uop_prs2},
     {ldq_13_bits_uop_prs2},
     {ldq_12_bits_uop_prs2},
     {ldq_11_bits_uop_prs2},
     {ldq_10_bits_uop_prs2},
     {ldq_9_bits_uop_prs2},
     {ldq_8_bits_uop_prs2},
     {ldq_7_bits_uop_prs2},
     {ldq_6_bits_uop_prs2},
     {ldq_5_bits_uop_prs2},
     {ldq_4_bits_uop_prs2},
     {ldq_3_bits_uop_prs2},
     {ldq_2_bits_uop_prs2},
     {ldq_1_bits_uop_prs2},
     {ldq_0_bits_uop_prs2}};	// lsu.scala:210:16, :465:79
  wire [31:0][6:0]  _GEN_157 =
    {{ldq_0_bits_uop_prs3},
     {ldq_0_bits_uop_prs3},
     {ldq_0_bits_uop_prs3},
     {ldq_0_bits_uop_prs3},
     {ldq_0_bits_uop_prs3},
     {ldq_0_bits_uop_prs3},
     {ldq_0_bits_uop_prs3},
     {ldq_0_bits_uop_prs3},
     {ldq_23_bits_uop_prs3},
     {ldq_22_bits_uop_prs3},
     {ldq_21_bits_uop_prs3},
     {ldq_20_bits_uop_prs3},
     {ldq_19_bits_uop_prs3},
     {ldq_18_bits_uop_prs3},
     {ldq_17_bits_uop_prs3},
     {ldq_16_bits_uop_prs3},
     {ldq_15_bits_uop_prs3},
     {ldq_14_bits_uop_prs3},
     {ldq_13_bits_uop_prs3},
     {ldq_12_bits_uop_prs3},
     {ldq_11_bits_uop_prs3},
     {ldq_10_bits_uop_prs3},
     {ldq_9_bits_uop_prs3},
     {ldq_8_bits_uop_prs3},
     {ldq_7_bits_uop_prs3},
     {ldq_6_bits_uop_prs3},
     {ldq_5_bits_uop_prs3},
     {ldq_4_bits_uop_prs3},
     {ldq_3_bits_uop_prs3},
     {ldq_2_bits_uop_prs3},
     {ldq_1_bits_uop_prs3},
     {ldq_0_bits_uop_prs3}};	// lsu.scala:210:16, :465:79
  wire [31:0][4:0]  _GEN_158 =
    {{ldq_0_bits_uop_ppred},
     {ldq_0_bits_uop_ppred},
     {ldq_0_bits_uop_ppred},
     {ldq_0_bits_uop_ppred},
     {ldq_0_bits_uop_ppred},
     {ldq_0_bits_uop_ppred},
     {ldq_0_bits_uop_ppred},
     {ldq_0_bits_uop_ppred},
     {ldq_23_bits_uop_ppred},
     {ldq_22_bits_uop_ppred},
     {ldq_21_bits_uop_ppred},
     {ldq_20_bits_uop_ppred},
     {ldq_19_bits_uop_ppred},
     {ldq_18_bits_uop_ppred},
     {ldq_17_bits_uop_ppred},
     {ldq_16_bits_uop_ppred},
     {ldq_15_bits_uop_ppred},
     {ldq_14_bits_uop_ppred},
     {ldq_13_bits_uop_ppred},
     {ldq_12_bits_uop_ppred},
     {ldq_11_bits_uop_ppred},
     {ldq_10_bits_uop_ppred},
     {ldq_9_bits_uop_ppred},
     {ldq_8_bits_uop_ppred},
     {ldq_7_bits_uop_ppred},
     {ldq_6_bits_uop_ppred},
     {ldq_5_bits_uop_ppred},
     {ldq_4_bits_uop_ppred},
     {ldq_3_bits_uop_ppred},
     {ldq_2_bits_uop_ppred},
     {ldq_1_bits_uop_ppred},
     {ldq_0_bits_uop_ppred}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_159 =
    {{ldq_0_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy},
     {ldq_23_bits_uop_prs1_busy},
     {ldq_22_bits_uop_prs1_busy},
     {ldq_21_bits_uop_prs1_busy},
     {ldq_20_bits_uop_prs1_busy},
     {ldq_19_bits_uop_prs1_busy},
     {ldq_18_bits_uop_prs1_busy},
     {ldq_17_bits_uop_prs1_busy},
     {ldq_16_bits_uop_prs1_busy},
     {ldq_15_bits_uop_prs1_busy},
     {ldq_14_bits_uop_prs1_busy},
     {ldq_13_bits_uop_prs1_busy},
     {ldq_12_bits_uop_prs1_busy},
     {ldq_11_bits_uop_prs1_busy},
     {ldq_10_bits_uop_prs1_busy},
     {ldq_9_bits_uop_prs1_busy},
     {ldq_8_bits_uop_prs1_busy},
     {ldq_7_bits_uop_prs1_busy},
     {ldq_6_bits_uop_prs1_busy},
     {ldq_5_bits_uop_prs1_busy},
     {ldq_4_bits_uop_prs1_busy},
     {ldq_3_bits_uop_prs1_busy},
     {ldq_2_bits_uop_prs1_busy},
     {ldq_1_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_160 =
    {{ldq_0_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy},
     {ldq_23_bits_uop_prs2_busy},
     {ldq_22_bits_uop_prs2_busy},
     {ldq_21_bits_uop_prs2_busy},
     {ldq_20_bits_uop_prs2_busy},
     {ldq_19_bits_uop_prs2_busy},
     {ldq_18_bits_uop_prs2_busy},
     {ldq_17_bits_uop_prs2_busy},
     {ldq_16_bits_uop_prs2_busy},
     {ldq_15_bits_uop_prs2_busy},
     {ldq_14_bits_uop_prs2_busy},
     {ldq_13_bits_uop_prs2_busy},
     {ldq_12_bits_uop_prs2_busy},
     {ldq_11_bits_uop_prs2_busy},
     {ldq_10_bits_uop_prs2_busy},
     {ldq_9_bits_uop_prs2_busy},
     {ldq_8_bits_uop_prs2_busy},
     {ldq_7_bits_uop_prs2_busy},
     {ldq_6_bits_uop_prs2_busy},
     {ldq_5_bits_uop_prs2_busy},
     {ldq_4_bits_uop_prs2_busy},
     {ldq_3_bits_uop_prs2_busy},
     {ldq_2_bits_uop_prs2_busy},
     {ldq_1_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_161 =
    {{ldq_0_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy},
     {ldq_23_bits_uop_prs3_busy},
     {ldq_22_bits_uop_prs3_busy},
     {ldq_21_bits_uop_prs3_busy},
     {ldq_20_bits_uop_prs3_busy},
     {ldq_19_bits_uop_prs3_busy},
     {ldq_18_bits_uop_prs3_busy},
     {ldq_17_bits_uop_prs3_busy},
     {ldq_16_bits_uop_prs3_busy},
     {ldq_15_bits_uop_prs3_busy},
     {ldq_14_bits_uop_prs3_busy},
     {ldq_13_bits_uop_prs3_busy},
     {ldq_12_bits_uop_prs3_busy},
     {ldq_11_bits_uop_prs3_busy},
     {ldq_10_bits_uop_prs3_busy},
     {ldq_9_bits_uop_prs3_busy},
     {ldq_8_bits_uop_prs3_busy},
     {ldq_7_bits_uop_prs3_busy},
     {ldq_6_bits_uop_prs3_busy},
     {ldq_5_bits_uop_prs3_busy},
     {ldq_4_bits_uop_prs3_busy},
     {ldq_3_bits_uop_prs3_busy},
     {ldq_2_bits_uop_prs3_busy},
     {ldq_1_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_162 =
    {{ldq_0_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy},
     {ldq_23_bits_uop_ppred_busy},
     {ldq_22_bits_uop_ppred_busy},
     {ldq_21_bits_uop_ppred_busy},
     {ldq_20_bits_uop_ppred_busy},
     {ldq_19_bits_uop_ppred_busy},
     {ldq_18_bits_uop_ppred_busy},
     {ldq_17_bits_uop_ppred_busy},
     {ldq_16_bits_uop_ppred_busy},
     {ldq_15_bits_uop_ppred_busy},
     {ldq_14_bits_uop_ppred_busy},
     {ldq_13_bits_uop_ppred_busy},
     {ldq_12_bits_uop_ppred_busy},
     {ldq_11_bits_uop_ppred_busy},
     {ldq_10_bits_uop_ppred_busy},
     {ldq_9_bits_uop_ppred_busy},
     {ldq_8_bits_uop_ppred_busy},
     {ldq_7_bits_uop_ppred_busy},
     {ldq_6_bits_uop_ppred_busy},
     {ldq_5_bits_uop_ppred_busy},
     {ldq_4_bits_uop_ppred_busy},
     {ldq_3_bits_uop_ppred_busy},
     {ldq_2_bits_uop_ppred_busy},
     {ldq_1_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy}};	// lsu.scala:210:16, :465:79
  wire [31:0][6:0]  _GEN_163 =
    {{ldq_0_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst},
     {ldq_23_bits_uop_stale_pdst},
     {ldq_22_bits_uop_stale_pdst},
     {ldq_21_bits_uop_stale_pdst},
     {ldq_20_bits_uop_stale_pdst},
     {ldq_19_bits_uop_stale_pdst},
     {ldq_18_bits_uop_stale_pdst},
     {ldq_17_bits_uop_stale_pdst},
     {ldq_16_bits_uop_stale_pdst},
     {ldq_15_bits_uop_stale_pdst},
     {ldq_14_bits_uop_stale_pdst},
     {ldq_13_bits_uop_stale_pdst},
     {ldq_12_bits_uop_stale_pdst},
     {ldq_11_bits_uop_stale_pdst},
     {ldq_10_bits_uop_stale_pdst},
     {ldq_9_bits_uop_stale_pdst},
     {ldq_8_bits_uop_stale_pdst},
     {ldq_7_bits_uop_stale_pdst},
     {ldq_6_bits_uop_stale_pdst},
     {ldq_5_bits_uop_stale_pdst},
     {ldq_4_bits_uop_stale_pdst},
     {ldq_3_bits_uop_stale_pdst},
     {ldq_2_bits_uop_stale_pdst},
     {ldq_1_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_164 =
    {{ldq_0_bits_uop_exception},
     {ldq_0_bits_uop_exception},
     {ldq_0_bits_uop_exception},
     {ldq_0_bits_uop_exception},
     {ldq_0_bits_uop_exception},
     {ldq_0_bits_uop_exception},
     {ldq_0_bits_uop_exception},
     {ldq_0_bits_uop_exception},
     {ldq_23_bits_uop_exception},
     {ldq_22_bits_uop_exception},
     {ldq_21_bits_uop_exception},
     {ldq_20_bits_uop_exception},
     {ldq_19_bits_uop_exception},
     {ldq_18_bits_uop_exception},
     {ldq_17_bits_uop_exception},
     {ldq_16_bits_uop_exception},
     {ldq_15_bits_uop_exception},
     {ldq_14_bits_uop_exception},
     {ldq_13_bits_uop_exception},
     {ldq_12_bits_uop_exception},
     {ldq_11_bits_uop_exception},
     {ldq_10_bits_uop_exception},
     {ldq_9_bits_uop_exception},
     {ldq_8_bits_uop_exception},
     {ldq_7_bits_uop_exception},
     {ldq_6_bits_uop_exception},
     {ldq_5_bits_uop_exception},
     {ldq_4_bits_uop_exception},
     {ldq_3_bits_uop_exception},
     {ldq_2_bits_uop_exception},
     {ldq_1_bits_uop_exception},
     {ldq_0_bits_uop_exception}};	// lsu.scala:210:16, :465:79
  wire [31:0][63:0] _GEN_165 =
    {{ldq_0_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause},
     {ldq_23_bits_uop_exc_cause},
     {ldq_22_bits_uop_exc_cause},
     {ldq_21_bits_uop_exc_cause},
     {ldq_20_bits_uop_exc_cause},
     {ldq_19_bits_uop_exc_cause},
     {ldq_18_bits_uop_exc_cause},
     {ldq_17_bits_uop_exc_cause},
     {ldq_16_bits_uop_exc_cause},
     {ldq_15_bits_uop_exc_cause},
     {ldq_14_bits_uop_exc_cause},
     {ldq_13_bits_uop_exc_cause},
     {ldq_12_bits_uop_exc_cause},
     {ldq_11_bits_uop_exc_cause},
     {ldq_10_bits_uop_exc_cause},
     {ldq_9_bits_uop_exc_cause},
     {ldq_8_bits_uop_exc_cause},
     {ldq_7_bits_uop_exc_cause},
     {ldq_6_bits_uop_exc_cause},
     {ldq_5_bits_uop_exc_cause},
     {ldq_4_bits_uop_exc_cause},
     {ldq_3_bits_uop_exc_cause},
     {ldq_2_bits_uop_exc_cause},
     {ldq_1_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_166 =
    {{ldq_0_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable},
     {ldq_23_bits_uop_bypassable},
     {ldq_22_bits_uop_bypassable},
     {ldq_21_bits_uop_bypassable},
     {ldq_20_bits_uop_bypassable},
     {ldq_19_bits_uop_bypassable},
     {ldq_18_bits_uop_bypassable},
     {ldq_17_bits_uop_bypassable},
     {ldq_16_bits_uop_bypassable},
     {ldq_15_bits_uop_bypassable},
     {ldq_14_bits_uop_bypassable},
     {ldq_13_bits_uop_bypassable},
     {ldq_12_bits_uop_bypassable},
     {ldq_11_bits_uop_bypassable},
     {ldq_10_bits_uop_bypassable},
     {ldq_9_bits_uop_bypassable},
     {ldq_8_bits_uop_bypassable},
     {ldq_7_bits_uop_bypassable},
     {ldq_6_bits_uop_bypassable},
     {ldq_5_bits_uop_bypassable},
     {ldq_4_bits_uop_bypassable},
     {ldq_3_bits_uop_bypassable},
     {ldq_2_bits_uop_bypassable},
     {ldq_1_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable}};	// lsu.scala:210:16, :465:79
  wire [31:0][4:0]  _GEN_167 =
    {{ldq_0_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd},
     {ldq_23_bits_uop_mem_cmd},
     {ldq_22_bits_uop_mem_cmd},
     {ldq_21_bits_uop_mem_cmd},
     {ldq_20_bits_uop_mem_cmd},
     {ldq_19_bits_uop_mem_cmd},
     {ldq_18_bits_uop_mem_cmd},
     {ldq_17_bits_uop_mem_cmd},
     {ldq_16_bits_uop_mem_cmd},
     {ldq_15_bits_uop_mem_cmd},
     {ldq_14_bits_uop_mem_cmd},
     {ldq_13_bits_uop_mem_cmd},
     {ldq_12_bits_uop_mem_cmd},
     {ldq_11_bits_uop_mem_cmd},
     {ldq_10_bits_uop_mem_cmd},
     {ldq_9_bits_uop_mem_cmd},
     {ldq_8_bits_uop_mem_cmd},
     {ldq_7_bits_uop_mem_cmd},
     {ldq_6_bits_uop_mem_cmd},
     {ldq_5_bits_uop_mem_cmd},
     {ldq_4_bits_uop_mem_cmd},
     {ldq_3_bits_uop_mem_cmd},
     {ldq_2_bits_uop_mem_cmd},
     {ldq_1_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd}};	// lsu.scala:210:16, :465:79
  wire [1:0]        mem_ldq_retry_e_out_bits_uop_mem_size = _GEN_112[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79
  wire [31:0]       _GEN_168 =
    {{ldq_0_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed},
     {ldq_23_bits_uop_mem_signed},
     {ldq_22_bits_uop_mem_signed},
     {ldq_21_bits_uop_mem_signed},
     {ldq_20_bits_uop_mem_signed},
     {ldq_19_bits_uop_mem_signed},
     {ldq_18_bits_uop_mem_signed},
     {ldq_17_bits_uop_mem_signed},
     {ldq_16_bits_uop_mem_signed},
     {ldq_15_bits_uop_mem_signed},
     {ldq_14_bits_uop_mem_signed},
     {ldq_13_bits_uop_mem_signed},
     {ldq_12_bits_uop_mem_signed},
     {ldq_11_bits_uop_mem_signed},
     {ldq_10_bits_uop_mem_signed},
     {ldq_9_bits_uop_mem_signed},
     {ldq_8_bits_uop_mem_signed},
     {ldq_7_bits_uop_mem_signed},
     {ldq_6_bits_uop_mem_signed},
     {ldq_5_bits_uop_mem_signed},
     {ldq_4_bits_uop_mem_signed},
     {ldq_3_bits_uop_mem_signed},
     {ldq_2_bits_uop_mem_signed},
     {ldq_1_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_169 =
    {{ldq_0_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence},
     {ldq_23_bits_uop_is_fence},
     {ldq_22_bits_uop_is_fence},
     {ldq_21_bits_uop_is_fence},
     {ldq_20_bits_uop_is_fence},
     {ldq_19_bits_uop_is_fence},
     {ldq_18_bits_uop_is_fence},
     {ldq_17_bits_uop_is_fence},
     {ldq_16_bits_uop_is_fence},
     {ldq_15_bits_uop_is_fence},
     {ldq_14_bits_uop_is_fence},
     {ldq_13_bits_uop_is_fence},
     {ldq_12_bits_uop_is_fence},
     {ldq_11_bits_uop_is_fence},
     {ldq_10_bits_uop_is_fence},
     {ldq_9_bits_uop_is_fence},
     {ldq_8_bits_uop_is_fence},
     {ldq_7_bits_uop_is_fence},
     {ldq_6_bits_uop_is_fence},
     {ldq_5_bits_uop_is_fence},
     {ldq_4_bits_uop_is_fence},
     {ldq_3_bits_uop_is_fence},
     {ldq_2_bits_uop_is_fence},
     {ldq_1_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_170 =
    {{ldq_0_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei},
     {ldq_23_bits_uop_is_fencei},
     {ldq_22_bits_uop_is_fencei},
     {ldq_21_bits_uop_is_fencei},
     {ldq_20_bits_uop_is_fencei},
     {ldq_19_bits_uop_is_fencei},
     {ldq_18_bits_uop_is_fencei},
     {ldq_17_bits_uop_is_fencei},
     {ldq_16_bits_uop_is_fencei},
     {ldq_15_bits_uop_is_fencei},
     {ldq_14_bits_uop_is_fencei},
     {ldq_13_bits_uop_is_fencei},
     {ldq_12_bits_uop_is_fencei},
     {ldq_11_bits_uop_is_fencei},
     {ldq_10_bits_uop_is_fencei},
     {ldq_9_bits_uop_is_fencei},
     {ldq_8_bits_uop_is_fencei},
     {ldq_7_bits_uop_is_fencei},
     {ldq_6_bits_uop_is_fencei},
     {ldq_5_bits_uop_is_fencei},
     {ldq_4_bits_uop_is_fencei},
     {ldq_3_bits_uop_is_fencei},
     {ldq_2_bits_uop_is_fencei},
     {ldq_1_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_171 =
    {{ldq_0_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo},
     {ldq_23_bits_uop_is_amo},
     {ldq_22_bits_uop_is_amo},
     {ldq_21_bits_uop_is_amo},
     {ldq_20_bits_uop_is_amo},
     {ldq_19_bits_uop_is_amo},
     {ldq_18_bits_uop_is_amo},
     {ldq_17_bits_uop_is_amo},
     {ldq_16_bits_uop_is_amo},
     {ldq_15_bits_uop_is_amo},
     {ldq_14_bits_uop_is_amo},
     {ldq_13_bits_uop_is_amo},
     {ldq_12_bits_uop_is_amo},
     {ldq_11_bits_uop_is_amo},
     {ldq_10_bits_uop_is_amo},
     {ldq_9_bits_uop_is_amo},
     {ldq_8_bits_uop_is_amo},
     {ldq_7_bits_uop_is_amo},
     {ldq_6_bits_uop_is_amo},
     {ldq_5_bits_uop_is_amo},
     {ldq_4_bits_uop_is_amo},
     {ldq_3_bits_uop_is_amo},
     {ldq_2_bits_uop_is_amo},
     {ldq_1_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_172 =
    {{ldq_0_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq},
     {ldq_23_bits_uop_uses_ldq},
     {ldq_22_bits_uop_uses_ldq},
     {ldq_21_bits_uop_uses_ldq},
     {ldq_20_bits_uop_uses_ldq},
     {ldq_19_bits_uop_uses_ldq},
     {ldq_18_bits_uop_uses_ldq},
     {ldq_17_bits_uop_uses_ldq},
     {ldq_16_bits_uop_uses_ldq},
     {ldq_15_bits_uop_uses_ldq},
     {ldq_14_bits_uop_uses_ldq},
     {ldq_13_bits_uop_uses_ldq},
     {ldq_12_bits_uop_uses_ldq},
     {ldq_11_bits_uop_uses_ldq},
     {ldq_10_bits_uop_uses_ldq},
     {ldq_9_bits_uop_uses_ldq},
     {ldq_8_bits_uop_uses_ldq},
     {ldq_7_bits_uop_uses_ldq},
     {ldq_6_bits_uop_uses_ldq},
     {ldq_5_bits_uop_uses_ldq},
     {ldq_4_bits_uop_uses_ldq},
     {ldq_3_bits_uop_uses_ldq},
     {ldq_2_bits_uop_uses_ldq},
     {ldq_1_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq}};	// lsu.scala:210:16, :465:79
  wire              _GEN_173 = _GEN_172[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [31:0]       _GEN_174 =
    {{ldq_0_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq},
     {ldq_23_bits_uop_uses_stq},
     {ldq_22_bits_uop_uses_stq},
     {ldq_21_bits_uop_uses_stq},
     {ldq_20_bits_uop_uses_stq},
     {ldq_19_bits_uop_uses_stq},
     {ldq_18_bits_uop_uses_stq},
     {ldq_17_bits_uop_uses_stq},
     {ldq_16_bits_uop_uses_stq},
     {ldq_15_bits_uop_uses_stq},
     {ldq_14_bits_uop_uses_stq},
     {ldq_13_bits_uop_uses_stq},
     {ldq_12_bits_uop_uses_stq},
     {ldq_11_bits_uop_uses_stq},
     {ldq_10_bits_uop_uses_stq},
     {ldq_9_bits_uop_uses_stq},
     {ldq_8_bits_uop_uses_stq},
     {ldq_7_bits_uop_uses_stq},
     {ldq_6_bits_uop_uses_stq},
     {ldq_5_bits_uop_uses_stq},
     {ldq_4_bits_uop_uses_stq},
     {ldq_3_bits_uop_uses_stq},
     {ldq_2_bits_uop_uses_stq},
     {ldq_1_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq}};	// lsu.scala:210:16, :465:79
  wire              _GEN_175 = _GEN_174[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [31:0]       _GEN_176 =
    {{ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc},
     {ldq_23_bits_uop_is_sys_pc2epc},
     {ldq_22_bits_uop_is_sys_pc2epc},
     {ldq_21_bits_uop_is_sys_pc2epc},
     {ldq_20_bits_uop_is_sys_pc2epc},
     {ldq_19_bits_uop_is_sys_pc2epc},
     {ldq_18_bits_uop_is_sys_pc2epc},
     {ldq_17_bits_uop_is_sys_pc2epc},
     {ldq_16_bits_uop_is_sys_pc2epc},
     {ldq_15_bits_uop_is_sys_pc2epc},
     {ldq_14_bits_uop_is_sys_pc2epc},
     {ldq_13_bits_uop_is_sys_pc2epc},
     {ldq_12_bits_uop_is_sys_pc2epc},
     {ldq_11_bits_uop_is_sys_pc2epc},
     {ldq_10_bits_uop_is_sys_pc2epc},
     {ldq_9_bits_uop_is_sys_pc2epc},
     {ldq_8_bits_uop_is_sys_pc2epc},
     {ldq_7_bits_uop_is_sys_pc2epc},
     {ldq_6_bits_uop_is_sys_pc2epc},
     {ldq_5_bits_uop_is_sys_pc2epc},
     {ldq_4_bits_uop_is_sys_pc2epc},
     {ldq_3_bits_uop_is_sys_pc2epc},
     {ldq_2_bits_uop_is_sys_pc2epc},
     {ldq_1_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_177 =
    {{ldq_0_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique},
     {ldq_23_bits_uop_is_unique},
     {ldq_22_bits_uop_is_unique},
     {ldq_21_bits_uop_is_unique},
     {ldq_20_bits_uop_is_unique},
     {ldq_19_bits_uop_is_unique},
     {ldq_18_bits_uop_is_unique},
     {ldq_17_bits_uop_is_unique},
     {ldq_16_bits_uop_is_unique},
     {ldq_15_bits_uop_is_unique},
     {ldq_14_bits_uop_is_unique},
     {ldq_13_bits_uop_is_unique},
     {ldq_12_bits_uop_is_unique},
     {ldq_11_bits_uop_is_unique},
     {ldq_10_bits_uop_is_unique},
     {ldq_9_bits_uop_is_unique},
     {ldq_8_bits_uop_is_unique},
     {ldq_7_bits_uop_is_unique},
     {ldq_6_bits_uop_is_unique},
     {ldq_5_bits_uop_is_unique},
     {ldq_4_bits_uop_is_unique},
     {ldq_3_bits_uop_is_unique},
     {ldq_2_bits_uop_is_unique},
     {ldq_1_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_178 =
    {{ldq_0_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit},
     {ldq_23_bits_uop_flush_on_commit},
     {ldq_22_bits_uop_flush_on_commit},
     {ldq_21_bits_uop_flush_on_commit},
     {ldq_20_bits_uop_flush_on_commit},
     {ldq_19_bits_uop_flush_on_commit},
     {ldq_18_bits_uop_flush_on_commit},
     {ldq_17_bits_uop_flush_on_commit},
     {ldq_16_bits_uop_flush_on_commit},
     {ldq_15_bits_uop_flush_on_commit},
     {ldq_14_bits_uop_flush_on_commit},
     {ldq_13_bits_uop_flush_on_commit},
     {ldq_12_bits_uop_flush_on_commit},
     {ldq_11_bits_uop_flush_on_commit},
     {ldq_10_bits_uop_flush_on_commit},
     {ldq_9_bits_uop_flush_on_commit},
     {ldq_8_bits_uop_flush_on_commit},
     {ldq_7_bits_uop_flush_on_commit},
     {ldq_6_bits_uop_flush_on_commit},
     {ldq_5_bits_uop_flush_on_commit},
     {ldq_4_bits_uop_flush_on_commit},
     {ldq_3_bits_uop_flush_on_commit},
     {ldq_2_bits_uop_flush_on_commit},
     {ldq_1_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_179 =
    {{ldq_0_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1},
     {ldq_23_bits_uop_ldst_is_rs1},
     {ldq_22_bits_uop_ldst_is_rs1},
     {ldq_21_bits_uop_ldst_is_rs1},
     {ldq_20_bits_uop_ldst_is_rs1},
     {ldq_19_bits_uop_ldst_is_rs1},
     {ldq_18_bits_uop_ldst_is_rs1},
     {ldq_17_bits_uop_ldst_is_rs1},
     {ldq_16_bits_uop_ldst_is_rs1},
     {ldq_15_bits_uop_ldst_is_rs1},
     {ldq_14_bits_uop_ldst_is_rs1},
     {ldq_13_bits_uop_ldst_is_rs1},
     {ldq_12_bits_uop_ldst_is_rs1},
     {ldq_11_bits_uop_ldst_is_rs1},
     {ldq_10_bits_uop_ldst_is_rs1},
     {ldq_9_bits_uop_ldst_is_rs1},
     {ldq_8_bits_uop_ldst_is_rs1},
     {ldq_7_bits_uop_ldst_is_rs1},
     {ldq_6_bits_uop_ldst_is_rs1},
     {ldq_5_bits_uop_ldst_is_rs1},
     {ldq_4_bits_uop_ldst_is_rs1},
     {ldq_3_bits_uop_ldst_is_rs1},
     {ldq_2_bits_uop_ldst_is_rs1},
     {ldq_1_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1}};	// lsu.scala:210:16, :465:79
  wire [31:0][5:0]  _GEN_180 =
    {{ldq_0_bits_uop_ldst},
     {ldq_0_bits_uop_ldst},
     {ldq_0_bits_uop_ldst},
     {ldq_0_bits_uop_ldst},
     {ldq_0_bits_uop_ldst},
     {ldq_0_bits_uop_ldst},
     {ldq_0_bits_uop_ldst},
     {ldq_0_bits_uop_ldst},
     {ldq_23_bits_uop_ldst},
     {ldq_22_bits_uop_ldst},
     {ldq_21_bits_uop_ldst},
     {ldq_20_bits_uop_ldst},
     {ldq_19_bits_uop_ldst},
     {ldq_18_bits_uop_ldst},
     {ldq_17_bits_uop_ldst},
     {ldq_16_bits_uop_ldst},
     {ldq_15_bits_uop_ldst},
     {ldq_14_bits_uop_ldst},
     {ldq_13_bits_uop_ldst},
     {ldq_12_bits_uop_ldst},
     {ldq_11_bits_uop_ldst},
     {ldq_10_bits_uop_ldst},
     {ldq_9_bits_uop_ldst},
     {ldq_8_bits_uop_ldst},
     {ldq_7_bits_uop_ldst},
     {ldq_6_bits_uop_ldst},
     {ldq_5_bits_uop_ldst},
     {ldq_4_bits_uop_ldst},
     {ldq_3_bits_uop_ldst},
     {ldq_2_bits_uop_ldst},
     {ldq_1_bits_uop_ldst},
     {ldq_0_bits_uop_ldst}};	// lsu.scala:210:16, :465:79
  wire [31:0][5:0]  _GEN_181 =
    {{ldq_0_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1},
     {ldq_23_bits_uop_lrs1},
     {ldq_22_bits_uop_lrs1},
     {ldq_21_bits_uop_lrs1},
     {ldq_20_bits_uop_lrs1},
     {ldq_19_bits_uop_lrs1},
     {ldq_18_bits_uop_lrs1},
     {ldq_17_bits_uop_lrs1},
     {ldq_16_bits_uop_lrs1},
     {ldq_15_bits_uop_lrs1},
     {ldq_14_bits_uop_lrs1},
     {ldq_13_bits_uop_lrs1},
     {ldq_12_bits_uop_lrs1},
     {ldq_11_bits_uop_lrs1},
     {ldq_10_bits_uop_lrs1},
     {ldq_9_bits_uop_lrs1},
     {ldq_8_bits_uop_lrs1},
     {ldq_7_bits_uop_lrs1},
     {ldq_6_bits_uop_lrs1},
     {ldq_5_bits_uop_lrs1},
     {ldq_4_bits_uop_lrs1},
     {ldq_3_bits_uop_lrs1},
     {ldq_2_bits_uop_lrs1},
     {ldq_1_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1}};	// lsu.scala:210:16, :465:79
  wire [31:0][5:0]  _GEN_182 =
    {{ldq_0_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2},
     {ldq_23_bits_uop_lrs2},
     {ldq_22_bits_uop_lrs2},
     {ldq_21_bits_uop_lrs2},
     {ldq_20_bits_uop_lrs2},
     {ldq_19_bits_uop_lrs2},
     {ldq_18_bits_uop_lrs2},
     {ldq_17_bits_uop_lrs2},
     {ldq_16_bits_uop_lrs2},
     {ldq_15_bits_uop_lrs2},
     {ldq_14_bits_uop_lrs2},
     {ldq_13_bits_uop_lrs2},
     {ldq_12_bits_uop_lrs2},
     {ldq_11_bits_uop_lrs2},
     {ldq_10_bits_uop_lrs2},
     {ldq_9_bits_uop_lrs2},
     {ldq_8_bits_uop_lrs2},
     {ldq_7_bits_uop_lrs2},
     {ldq_6_bits_uop_lrs2},
     {ldq_5_bits_uop_lrs2},
     {ldq_4_bits_uop_lrs2},
     {ldq_3_bits_uop_lrs2},
     {ldq_2_bits_uop_lrs2},
     {ldq_1_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2}};	// lsu.scala:210:16, :465:79
  wire [31:0][5:0]  _GEN_183 =
    {{ldq_0_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3},
     {ldq_23_bits_uop_lrs3},
     {ldq_22_bits_uop_lrs3},
     {ldq_21_bits_uop_lrs3},
     {ldq_20_bits_uop_lrs3},
     {ldq_19_bits_uop_lrs3},
     {ldq_18_bits_uop_lrs3},
     {ldq_17_bits_uop_lrs3},
     {ldq_16_bits_uop_lrs3},
     {ldq_15_bits_uop_lrs3},
     {ldq_14_bits_uop_lrs3},
     {ldq_13_bits_uop_lrs3},
     {ldq_12_bits_uop_lrs3},
     {ldq_11_bits_uop_lrs3},
     {ldq_10_bits_uop_lrs3},
     {ldq_9_bits_uop_lrs3},
     {ldq_8_bits_uop_lrs3},
     {ldq_7_bits_uop_lrs3},
     {ldq_6_bits_uop_lrs3},
     {ldq_5_bits_uop_lrs3},
     {ldq_4_bits_uop_lrs3},
     {ldq_3_bits_uop_lrs3},
     {ldq_2_bits_uop_lrs3},
     {ldq_1_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_184 =
    {{ldq_0_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val},
     {ldq_23_bits_uop_ldst_val},
     {ldq_22_bits_uop_ldst_val},
     {ldq_21_bits_uop_ldst_val},
     {ldq_20_bits_uop_ldst_val},
     {ldq_19_bits_uop_ldst_val},
     {ldq_18_bits_uop_ldst_val},
     {ldq_17_bits_uop_ldst_val},
     {ldq_16_bits_uop_ldst_val},
     {ldq_15_bits_uop_ldst_val},
     {ldq_14_bits_uop_ldst_val},
     {ldq_13_bits_uop_ldst_val},
     {ldq_12_bits_uop_ldst_val},
     {ldq_11_bits_uop_ldst_val},
     {ldq_10_bits_uop_ldst_val},
     {ldq_9_bits_uop_ldst_val},
     {ldq_8_bits_uop_ldst_val},
     {ldq_7_bits_uop_ldst_val},
     {ldq_6_bits_uop_ldst_val},
     {ldq_5_bits_uop_ldst_val},
     {ldq_4_bits_uop_ldst_val},
     {ldq_3_bits_uop_ldst_val},
     {ldq_2_bits_uop_ldst_val},
     {ldq_1_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val}};	// lsu.scala:210:16, :465:79
  wire [31:0][1:0]  _GEN_185 =
    {{ldq_0_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype},
     {ldq_23_bits_uop_dst_rtype},
     {ldq_22_bits_uop_dst_rtype},
     {ldq_21_bits_uop_dst_rtype},
     {ldq_20_bits_uop_dst_rtype},
     {ldq_19_bits_uop_dst_rtype},
     {ldq_18_bits_uop_dst_rtype},
     {ldq_17_bits_uop_dst_rtype},
     {ldq_16_bits_uop_dst_rtype},
     {ldq_15_bits_uop_dst_rtype},
     {ldq_14_bits_uop_dst_rtype},
     {ldq_13_bits_uop_dst_rtype},
     {ldq_12_bits_uop_dst_rtype},
     {ldq_11_bits_uop_dst_rtype},
     {ldq_10_bits_uop_dst_rtype},
     {ldq_9_bits_uop_dst_rtype},
     {ldq_8_bits_uop_dst_rtype},
     {ldq_7_bits_uop_dst_rtype},
     {ldq_6_bits_uop_dst_rtype},
     {ldq_5_bits_uop_dst_rtype},
     {ldq_4_bits_uop_dst_rtype},
     {ldq_3_bits_uop_dst_rtype},
     {ldq_2_bits_uop_dst_rtype},
     {ldq_1_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype}};	// lsu.scala:210:16, :465:79
  wire [31:0][1:0]  _GEN_186 =
    {{ldq_0_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype},
     {ldq_23_bits_uop_lrs1_rtype},
     {ldq_22_bits_uop_lrs1_rtype},
     {ldq_21_bits_uop_lrs1_rtype},
     {ldq_20_bits_uop_lrs1_rtype},
     {ldq_19_bits_uop_lrs1_rtype},
     {ldq_18_bits_uop_lrs1_rtype},
     {ldq_17_bits_uop_lrs1_rtype},
     {ldq_16_bits_uop_lrs1_rtype},
     {ldq_15_bits_uop_lrs1_rtype},
     {ldq_14_bits_uop_lrs1_rtype},
     {ldq_13_bits_uop_lrs1_rtype},
     {ldq_12_bits_uop_lrs1_rtype},
     {ldq_11_bits_uop_lrs1_rtype},
     {ldq_10_bits_uop_lrs1_rtype},
     {ldq_9_bits_uop_lrs1_rtype},
     {ldq_8_bits_uop_lrs1_rtype},
     {ldq_7_bits_uop_lrs1_rtype},
     {ldq_6_bits_uop_lrs1_rtype},
     {ldq_5_bits_uop_lrs1_rtype},
     {ldq_4_bits_uop_lrs1_rtype},
     {ldq_3_bits_uop_lrs1_rtype},
     {ldq_2_bits_uop_lrs1_rtype},
     {ldq_1_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype}};	// lsu.scala:210:16, :465:79
  wire [31:0][1:0]  _GEN_187 =
    {{ldq_0_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype},
     {ldq_23_bits_uop_lrs2_rtype},
     {ldq_22_bits_uop_lrs2_rtype},
     {ldq_21_bits_uop_lrs2_rtype},
     {ldq_20_bits_uop_lrs2_rtype},
     {ldq_19_bits_uop_lrs2_rtype},
     {ldq_18_bits_uop_lrs2_rtype},
     {ldq_17_bits_uop_lrs2_rtype},
     {ldq_16_bits_uop_lrs2_rtype},
     {ldq_15_bits_uop_lrs2_rtype},
     {ldq_14_bits_uop_lrs2_rtype},
     {ldq_13_bits_uop_lrs2_rtype},
     {ldq_12_bits_uop_lrs2_rtype},
     {ldq_11_bits_uop_lrs2_rtype},
     {ldq_10_bits_uop_lrs2_rtype},
     {ldq_9_bits_uop_lrs2_rtype},
     {ldq_8_bits_uop_lrs2_rtype},
     {ldq_7_bits_uop_lrs2_rtype},
     {ldq_6_bits_uop_lrs2_rtype},
     {ldq_5_bits_uop_lrs2_rtype},
     {ldq_4_bits_uop_lrs2_rtype},
     {ldq_3_bits_uop_lrs2_rtype},
     {ldq_2_bits_uop_lrs2_rtype},
     {ldq_1_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_188 =
    {{ldq_0_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en},
     {ldq_23_bits_uop_frs3_en},
     {ldq_22_bits_uop_frs3_en},
     {ldq_21_bits_uop_frs3_en},
     {ldq_20_bits_uop_frs3_en},
     {ldq_19_bits_uop_frs3_en},
     {ldq_18_bits_uop_frs3_en},
     {ldq_17_bits_uop_frs3_en},
     {ldq_16_bits_uop_frs3_en},
     {ldq_15_bits_uop_frs3_en},
     {ldq_14_bits_uop_frs3_en},
     {ldq_13_bits_uop_frs3_en},
     {ldq_12_bits_uop_frs3_en},
     {ldq_11_bits_uop_frs3_en},
     {ldq_10_bits_uop_frs3_en},
     {ldq_9_bits_uop_frs3_en},
     {ldq_8_bits_uop_frs3_en},
     {ldq_7_bits_uop_frs3_en},
     {ldq_6_bits_uop_frs3_en},
     {ldq_5_bits_uop_frs3_en},
     {ldq_4_bits_uop_frs3_en},
     {ldq_3_bits_uop_frs3_en},
     {ldq_2_bits_uop_frs3_en},
     {ldq_1_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_189 =
    {{ldq_0_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val},
     {ldq_23_bits_uop_fp_val},
     {ldq_22_bits_uop_fp_val},
     {ldq_21_bits_uop_fp_val},
     {ldq_20_bits_uop_fp_val},
     {ldq_19_bits_uop_fp_val},
     {ldq_18_bits_uop_fp_val},
     {ldq_17_bits_uop_fp_val},
     {ldq_16_bits_uop_fp_val},
     {ldq_15_bits_uop_fp_val},
     {ldq_14_bits_uop_fp_val},
     {ldq_13_bits_uop_fp_val},
     {ldq_12_bits_uop_fp_val},
     {ldq_11_bits_uop_fp_val},
     {ldq_10_bits_uop_fp_val},
     {ldq_9_bits_uop_fp_val},
     {ldq_8_bits_uop_fp_val},
     {ldq_7_bits_uop_fp_val},
     {ldq_6_bits_uop_fp_val},
     {ldq_5_bits_uop_fp_val},
     {ldq_4_bits_uop_fp_val},
     {ldq_3_bits_uop_fp_val},
     {ldq_2_bits_uop_fp_val},
     {ldq_1_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_190 =
    {{ldq_0_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single},
     {ldq_23_bits_uop_fp_single},
     {ldq_22_bits_uop_fp_single},
     {ldq_21_bits_uop_fp_single},
     {ldq_20_bits_uop_fp_single},
     {ldq_19_bits_uop_fp_single},
     {ldq_18_bits_uop_fp_single},
     {ldq_17_bits_uop_fp_single},
     {ldq_16_bits_uop_fp_single},
     {ldq_15_bits_uop_fp_single},
     {ldq_14_bits_uop_fp_single},
     {ldq_13_bits_uop_fp_single},
     {ldq_12_bits_uop_fp_single},
     {ldq_11_bits_uop_fp_single},
     {ldq_10_bits_uop_fp_single},
     {ldq_9_bits_uop_fp_single},
     {ldq_8_bits_uop_fp_single},
     {ldq_7_bits_uop_fp_single},
     {ldq_6_bits_uop_fp_single},
     {ldq_5_bits_uop_fp_single},
     {ldq_4_bits_uop_fp_single},
     {ldq_3_bits_uop_fp_single},
     {ldq_2_bits_uop_fp_single},
     {ldq_1_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_191 =
    {{ldq_0_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if},
     {ldq_23_bits_uop_xcpt_pf_if},
     {ldq_22_bits_uop_xcpt_pf_if},
     {ldq_21_bits_uop_xcpt_pf_if},
     {ldq_20_bits_uop_xcpt_pf_if},
     {ldq_19_bits_uop_xcpt_pf_if},
     {ldq_18_bits_uop_xcpt_pf_if},
     {ldq_17_bits_uop_xcpt_pf_if},
     {ldq_16_bits_uop_xcpt_pf_if},
     {ldq_15_bits_uop_xcpt_pf_if},
     {ldq_14_bits_uop_xcpt_pf_if},
     {ldq_13_bits_uop_xcpt_pf_if},
     {ldq_12_bits_uop_xcpt_pf_if},
     {ldq_11_bits_uop_xcpt_pf_if},
     {ldq_10_bits_uop_xcpt_pf_if},
     {ldq_9_bits_uop_xcpt_pf_if},
     {ldq_8_bits_uop_xcpt_pf_if},
     {ldq_7_bits_uop_xcpt_pf_if},
     {ldq_6_bits_uop_xcpt_pf_if},
     {ldq_5_bits_uop_xcpt_pf_if},
     {ldq_4_bits_uop_xcpt_pf_if},
     {ldq_3_bits_uop_xcpt_pf_if},
     {ldq_2_bits_uop_xcpt_pf_if},
     {ldq_1_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_192 =
    {{ldq_0_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if},
     {ldq_23_bits_uop_xcpt_ae_if},
     {ldq_22_bits_uop_xcpt_ae_if},
     {ldq_21_bits_uop_xcpt_ae_if},
     {ldq_20_bits_uop_xcpt_ae_if},
     {ldq_19_bits_uop_xcpt_ae_if},
     {ldq_18_bits_uop_xcpt_ae_if},
     {ldq_17_bits_uop_xcpt_ae_if},
     {ldq_16_bits_uop_xcpt_ae_if},
     {ldq_15_bits_uop_xcpt_ae_if},
     {ldq_14_bits_uop_xcpt_ae_if},
     {ldq_13_bits_uop_xcpt_ae_if},
     {ldq_12_bits_uop_xcpt_ae_if},
     {ldq_11_bits_uop_xcpt_ae_if},
     {ldq_10_bits_uop_xcpt_ae_if},
     {ldq_9_bits_uop_xcpt_ae_if},
     {ldq_8_bits_uop_xcpt_ae_if},
     {ldq_7_bits_uop_xcpt_ae_if},
     {ldq_6_bits_uop_xcpt_ae_if},
     {ldq_5_bits_uop_xcpt_ae_if},
     {ldq_4_bits_uop_xcpt_ae_if},
     {ldq_3_bits_uop_xcpt_ae_if},
     {ldq_2_bits_uop_xcpt_ae_if},
     {ldq_1_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_193 =
    {{ldq_0_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if},
     {ldq_23_bits_uop_xcpt_ma_if},
     {ldq_22_bits_uop_xcpt_ma_if},
     {ldq_21_bits_uop_xcpt_ma_if},
     {ldq_20_bits_uop_xcpt_ma_if},
     {ldq_19_bits_uop_xcpt_ma_if},
     {ldq_18_bits_uop_xcpt_ma_if},
     {ldq_17_bits_uop_xcpt_ma_if},
     {ldq_16_bits_uop_xcpt_ma_if},
     {ldq_15_bits_uop_xcpt_ma_if},
     {ldq_14_bits_uop_xcpt_ma_if},
     {ldq_13_bits_uop_xcpt_ma_if},
     {ldq_12_bits_uop_xcpt_ma_if},
     {ldq_11_bits_uop_xcpt_ma_if},
     {ldq_10_bits_uop_xcpt_ma_if},
     {ldq_9_bits_uop_xcpt_ma_if},
     {ldq_8_bits_uop_xcpt_ma_if},
     {ldq_7_bits_uop_xcpt_ma_if},
     {ldq_6_bits_uop_xcpt_ma_if},
     {ldq_5_bits_uop_xcpt_ma_if},
     {ldq_4_bits_uop_xcpt_ma_if},
     {ldq_3_bits_uop_xcpt_ma_if},
     {ldq_2_bits_uop_xcpt_ma_if},
     {ldq_1_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_194 =
    {{ldq_0_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if},
     {ldq_23_bits_uop_bp_debug_if},
     {ldq_22_bits_uop_bp_debug_if},
     {ldq_21_bits_uop_bp_debug_if},
     {ldq_20_bits_uop_bp_debug_if},
     {ldq_19_bits_uop_bp_debug_if},
     {ldq_18_bits_uop_bp_debug_if},
     {ldq_17_bits_uop_bp_debug_if},
     {ldq_16_bits_uop_bp_debug_if},
     {ldq_15_bits_uop_bp_debug_if},
     {ldq_14_bits_uop_bp_debug_if},
     {ldq_13_bits_uop_bp_debug_if},
     {ldq_12_bits_uop_bp_debug_if},
     {ldq_11_bits_uop_bp_debug_if},
     {ldq_10_bits_uop_bp_debug_if},
     {ldq_9_bits_uop_bp_debug_if},
     {ldq_8_bits_uop_bp_debug_if},
     {ldq_7_bits_uop_bp_debug_if},
     {ldq_6_bits_uop_bp_debug_if},
     {ldq_5_bits_uop_bp_debug_if},
     {ldq_4_bits_uop_bp_debug_if},
     {ldq_3_bits_uop_bp_debug_if},
     {ldq_2_bits_uop_bp_debug_if},
     {ldq_1_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_195 =
    {{ldq_0_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if},
     {ldq_23_bits_uop_bp_xcpt_if},
     {ldq_22_bits_uop_bp_xcpt_if},
     {ldq_21_bits_uop_bp_xcpt_if},
     {ldq_20_bits_uop_bp_xcpt_if},
     {ldq_19_bits_uop_bp_xcpt_if},
     {ldq_18_bits_uop_bp_xcpt_if},
     {ldq_17_bits_uop_bp_xcpt_if},
     {ldq_16_bits_uop_bp_xcpt_if},
     {ldq_15_bits_uop_bp_xcpt_if},
     {ldq_14_bits_uop_bp_xcpt_if},
     {ldq_13_bits_uop_bp_xcpt_if},
     {ldq_12_bits_uop_bp_xcpt_if},
     {ldq_11_bits_uop_bp_xcpt_if},
     {ldq_10_bits_uop_bp_xcpt_if},
     {ldq_9_bits_uop_bp_xcpt_if},
     {ldq_8_bits_uop_bp_xcpt_if},
     {ldq_7_bits_uop_bp_xcpt_if},
     {ldq_6_bits_uop_bp_xcpt_if},
     {ldq_5_bits_uop_bp_xcpt_if},
     {ldq_4_bits_uop_bp_xcpt_if},
     {ldq_3_bits_uop_bp_xcpt_if},
     {ldq_2_bits_uop_bp_xcpt_if},
     {ldq_1_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if}};	// lsu.scala:210:16, :465:79
  wire [31:0][1:0]  _GEN_196 =
    {{ldq_0_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc},
     {ldq_23_bits_uop_debug_fsrc},
     {ldq_22_bits_uop_debug_fsrc},
     {ldq_21_bits_uop_debug_fsrc},
     {ldq_20_bits_uop_debug_fsrc},
     {ldq_19_bits_uop_debug_fsrc},
     {ldq_18_bits_uop_debug_fsrc},
     {ldq_17_bits_uop_debug_fsrc},
     {ldq_16_bits_uop_debug_fsrc},
     {ldq_15_bits_uop_debug_fsrc},
     {ldq_14_bits_uop_debug_fsrc},
     {ldq_13_bits_uop_debug_fsrc},
     {ldq_12_bits_uop_debug_fsrc},
     {ldq_11_bits_uop_debug_fsrc},
     {ldq_10_bits_uop_debug_fsrc},
     {ldq_9_bits_uop_debug_fsrc},
     {ldq_8_bits_uop_debug_fsrc},
     {ldq_7_bits_uop_debug_fsrc},
     {ldq_6_bits_uop_debug_fsrc},
     {ldq_5_bits_uop_debug_fsrc},
     {ldq_4_bits_uop_debug_fsrc},
     {ldq_3_bits_uop_debug_fsrc},
     {ldq_2_bits_uop_debug_fsrc},
     {ldq_1_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc}};	// lsu.scala:210:16, :465:79
  wire [31:0][1:0]  _GEN_197 =
    {{ldq_0_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc},
     {ldq_23_bits_uop_debug_tsrc},
     {ldq_22_bits_uop_debug_tsrc},
     {ldq_21_bits_uop_debug_tsrc},
     {ldq_20_bits_uop_debug_tsrc},
     {ldq_19_bits_uop_debug_tsrc},
     {ldq_18_bits_uop_debug_tsrc},
     {ldq_17_bits_uop_debug_tsrc},
     {ldq_16_bits_uop_debug_tsrc},
     {ldq_15_bits_uop_debug_tsrc},
     {ldq_14_bits_uop_debug_tsrc},
     {ldq_13_bits_uop_debug_tsrc},
     {ldq_12_bits_uop_debug_tsrc},
     {ldq_11_bits_uop_debug_tsrc},
     {ldq_10_bits_uop_debug_tsrc},
     {ldq_9_bits_uop_debug_tsrc},
     {ldq_8_bits_uop_debug_tsrc},
     {ldq_7_bits_uop_debug_tsrc},
     {ldq_6_bits_uop_debug_tsrc},
     {ldq_5_bits_uop_debug_tsrc},
     {ldq_4_bits_uop_debug_tsrc},
     {ldq_3_bits_uop_debug_tsrc},
     {ldq_2_bits_uop_debug_tsrc},
     {ldq_1_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc}};	// lsu.scala:210:16, :465:79
  wire [31:0][39:0] _GEN_198 =
    {{ldq_0_bits_addr_bits},
     {ldq_0_bits_addr_bits},
     {ldq_0_bits_addr_bits},
     {ldq_0_bits_addr_bits},
     {ldq_0_bits_addr_bits},
     {ldq_0_bits_addr_bits},
     {ldq_0_bits_addr_bits},
     {ldq_0_bits_addr_bits},
     {ldq_23_bits_addr_bits},
     {ldq_22_bits_addr_bits},
     {ldq_21_bits_addr_bits},
     {ldq_20_bits_addr_bits},
     {ldq_19_bits_addr_bits},
     {ldq_18_bits_addr_bits},
     {ldq_17_bits_addr_bits},
     {ldq_16_bits_addr_bits},
     {ldq_15_bits_addr_bits},
     {ldq_14_bits_addr_bits},
     {ldq_13_bits_addr_bits},
     {ldq_12_bits_addr_bits},
     {ldq_11_bits_addr_bits},
     {ldq_10_bits_addr_bits},
     {ldq_9_bits_addr_bits},
     {ldq_8_bits_addr_bits},
     {ldq_7_bits_addr_bits},
     {ldq_6_bits_addr_bits},
     {ldq_5_bits_addr_bits},
     {ldq_4_bits_addr_bits},
     {ldq_3_bits_addr_bits},
     {ldq_2_bits_addr_bits},
     {ldq_1_bits_addr_bits},
     {ldq_0_bits_addr_bits}};	// lsu.scala:210:16, :465:79
  wire [39:0]       _GEN_199 = _GEN_198[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [31:0]       _GEN_200 =
    {{ldq_0_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual},
     {ldq_23_bits_addr_is_virtual},
     {ldq_22_bits_addr_is_virtual},
     {ldq_21_bits_addr_is_virtual},
     {ldq_20_bits_addr_is_virtual},
     {ldq_19_bits_addr_is_virtual},
     {ldq_18_bits_addr_is_virtual},
     {ldq_17_bits_addr_is_virtual},
     {ldq_16_bits_addr_is_virtual},
     {ldq_15_bits_addr_is_virtual},
     {ldq_14_bits_addr_is_virtual},
     {ldq_13_bits_addr_is_virtual},
     {ldq_12_bits_addr_is_virtual},
     {ldq_11_bits_addr_is_virtual},
     {ldq_10_bits_addr_is_virtual},
     {ldq_9_bits_addr_is_virtual},
     {ldq_8_bits_addr_is_virtual},
     {ldq_7_bits_addr_is_virtual},
     {ldq_6_bits_addr_is_virtual},
     {ldq_5_bits_addr_is_virtual},
     {ldq_4_bits_addr_is_virtual},
     {ldq_3_bits_addr_is_virtual},
     {ldq_2_bits_addr_is_virtual},
     {ldq_1_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_201 =
    {{ldq_0_bits_order_fail},
     {ldq_0_bits_order_fail},
     {ldq_0_bits_order_fail},
     {ldq_0_bits_order_fail},
     {ldq_0_bits_order_fail},
     {ldq_0_bits_order_fail},
     {ldq_0_bits_order_fail},
     {ldq_0_bits_order_fail},
     {ldq_23_bits_order_fail},
     {ldq_22_bits_order_fail},
     {ldq_21_bits_order_fail},
     {ldq_20_bits_order_fail},
     {ldq_19_bits_order_fail},
     {ldq_18_bits_order_fail},
     {ldq_17_bits_order_fail},
     {ldq_16_bits_order_fail},
     {ldq_15_bits_order_fail},
     {ldq_14_bits_order_fail},
     {ldq_13_bits_order_fail},
     {ldq_12_bits_order_fail},
     {ldq_11_bits_order_fail},
     {ldq_10_bits_order_fail},
     {ldq_9_bits_order_fail},
     {ldq_8_bits_order_fail},
     {ldq_7_bits_order_fail},
     {ldq_6_bits_order_fail},
     {ldq_5_bits_order_fail},
     {ldq_4_bits_order_fail},
     {ldq_3_bits_order_fail},
     {ldq_2_bits_order_fail},
     {ldq_1_bits_order_fail},
     {ldq_0_bits_order_fail}};	// lsu.scala:210:16, :465:79
  wire [31:0]       _GEN_202 =
    {{p1_block_load_mask_0},
     {p1_block_load_mask_0},
     {p1_block_load_mask_0},
     {p1_block_load_mask_0},
     {p1_block_load_mask_0},
     {p1_block_load_mask_0},
     {p1_block_load_mask_0},
     {p1_block_load_mask_0},
     {p1_block_load_mask_23},
     {p1_block_load_mask_22},
     {p1_block_load_mask_21},
     {p1_block_load_mask_20},
     {p1_block_load_mask_19},
     {p1_block_load_mask_18},
     {p1_block_load_mask_17},
     {p1_block_load_mask_16},
     {p1_block_load_mask_15},
     {p1_block_load_mask_14},
     {p1_block_load_mask_13},
     {p1_block_load_mask_12},
     {p1_block_load_mask_11},
     {p1_block_load_mask_10},
     {p1_block_load_mask_9},
     {p1_block_load_mask_8},
     {p1_block_load_mask_7},
     {p1_block_load_mask_6},
     {p1_block_load_mask_5},
     {p1_block_load_mask_4},
     {p1_block_load_mask_3},
     {p1_block_load_mask_2},
     {p1_block_load_mask_1},
     {p1_block_load_mask_0}};	// lsu.scala:398:35, :468:33
  wire [31:0]       _GEN_203 =
    {{p2_block_load_mask_0},
     {p2_block_load_mask_0},
     {p2_block_load_mask_0},
     {p2_block_load_mask_0},
     {p2_block_load_mask_0},
     {p2_block_load_mask_0},
     {p2_block_load_mask_0},
     {p2_block_load_mask_0},
     {p2_block_load_mask_23},
     {p2_block_load_mask_22},
     {p2_block_load_mask_21},
     {p2_block_load_mask_20},
     {p2_block_load_mask_19},
     {p2_block_load_mask_18},
     {p2_block_load_mask_17},
     {p2_block_load_mask_16},
     {p2_block_load_mask_15},
     {p2_block_load_mask_14},
     {p2_block_load_mask_13},
     {p2_block_load_mask_12},
     {p2_block_load_mask_11},
     {p2_block_load_mask_10},
     {p2_block_load_mask_9},
     {p2_block_load_mask_8},
     {p2_block_load_mask_7},
     {p2_block_load_mask_6},
     {p2_block_load_mask_5},
     {p2_block_load_mask_4},
     {p2_block_load_mask_3},
     {p2_block_load_mask_2},
     {p2_block_load_mask_1},
     {p2_block_load_mask_0}};	// lsu.scala:399:35, :469:33
  reg               can_fire_load_retry_REG;	// lsu.scala:470:40
  wire              _GEN_204 = _GEN_2[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [15:0]       _GEN_205 = _GEN_28[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [6:0]        mem_stq_retry_e_out_bits_uop_rob_idx = _GEN_36[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [4:0]        _GEN_206 = _GEN_37[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [4:0]        mem_stq_retry_e_out_bits_uop_stq_idx = _GEN_38[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [6:0]        _GEN_207 = _GEN_40[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [1:0]        mem_stq_retry_e_out_bits_uop_mem_size = _GEN_55[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire              mem_stq_retry_e_out_bits_uop_is_amo = _GEN_61[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [39:0]       _GEN_208 = _GEN_88[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  reg               can_fire_sta_retry_REG;	// lsu.scala:482:41
  wire              can_fire_store_commit_0 =
    _GEN_3 & ~_GEN_59 & ~mem_xcpt_valids_0 & ~_GEN_51
    & (_GEN_94[stq_execute_head] | _GEN_62 & _GEN_87[stq_execute_head]
       & ~_GEN_90[stq_execute_head] & _GEN_91[stq_execute_head]);	// lsu.scala:220:29, :224:42, :490:33, :491:33, :492:33, :493:79, :494:62, :496:{66,101}, :667:32
  wire [15:0]       _GEN_209 = _GEN_110[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [4:0]        mem_ldq_wakeup_e_out_bits_uop_stq_idx = _GEN_111[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [1:0]        mem_ldq_wakeup_e_out_bits_uop_mem_size = _GEN_112[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [39:0]       _GEN_210 = _GEN_198[ldq_wakeup_idx];	// lsu.scala:430:31, :465:79, :502:88
  wire              _GEN_211 = _GEN_200[ldq_wakeup_idx];	// lsu.scala:430:31, :465:79, :502:88
  wire [31:0]       _GEN_212 =
    {{ldq_0_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable},
     {ldq_23_bits_addr_is_uncacheable},
     {ldq_22_bits_addr_is_uncacheable},
     {ldq_21_bits_addr_is_uncacheable},
     {ldq_20_bits_addr_is_uncacheable},
     {ldq_19_bits_addr_is_uncacheable},
     {ldq_18_bits_addr_is_uncacheable},
     {ldq_17_bits_addr_is_uncacheable},
     {ldq_16_bits_addr_is_uncacheable},
     {ldq_15_bits_addr_is_uncacheable},
     {ldq_14_bits_addr_is_uncacheable},
     {ldq_13_bits_addr_is_uncacheable},
     {ldq_12_bits_addr_is_uncacheable},
     {ldq_11_bits_addr_is_uncacheable},
     {ldq_10_bits_addr_is_uncacheable},
     {ldq_9_bits_addr_is_uncacheable},
     {ldq_8_bits_addr_is_uncacheable},
     {ldq_7_bits_addr_is_uncacheable},
     {ldq_6_bits_addr_is_uncacheable},
     {ldq_5_bits_addr_is_uncacheable},
     {ldq_4_bits_addr_is_uncacheable},
     {ldq_3_bits_addr_is_uncacheable},
     {ldq_2_bits_addr_is_uncacheable},
     {ldq_1_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable}};	// lsu.scala:210:16, :502:88
  wire              _GEN_213 = _GEN_114[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [31:0]       _GEN_214 =
    {{ldq_0_bits_succeeded},
     {ldq_0_bits_succeeded},
     {ldq_0_bits_succeeded},
     {ldq_0_bits_succeeded},
     {ldq_0_bits_succeeded},
     {ldq_0_bits_succeeded},
     {ldq_0_bits_succeeded},
     {ldq_0_bits_succeeded},
     {ldq_23_bits_succeeded},
     {ldq_22_bits_succeeded},
     {ldq_21_bits_succeeded},
     {ldq_20_bits_succeeded},
     {ldq_19_bits_succeeded},
     {ldq_18_bits_succeeded},
     {ldq_17_bits_succeeded},
     {ldq_16_bits_succeeded},
     {ldq_15_bits_succeeded},
     {ldq_14_bits_succeeded},
     {ldq_13_bits_succeeded},
     {ldq_12_bits_succeeded},
     {ldq_11_bits_succeeded},
     {ldq_10_bits_succeeded},
     {ldq_9_bits_succeeded},
     {ldq_8_bits_succeeded},
     {ldq_7_bits_succeeded},
     {ldq_6_bits_succeeded},
     {ldq_5_bits_succeeded},
     {ldq_4_bits_succeeded},
     {ldq_3_bits_succeeded},
     {ldq_2_bits_succeeded},
     {ldq_1_bits_succeeded},
     {ldq_0_bits_succeeded}};	// lsu.scala:210:16, :502:88
  wire [23:0]       mem_ldq_wakeup_e_out_bits_st_dep_mask = _GEN_115[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire              will_fire_stad_incoming_0 =
    _can_fire_sta_incoming_T & io_core_exe_0_req_bits_uop_ctrl_is_std
    & ~can_fire_load_incoming_0 & ~can_fire_load_incoming_0;	// lsu.scala:441:63, :444:63, :534:{35,63}, :535:35
  wire              _will_fire_sta_incoming_0_will_fire_T_2 =
    ~can_fire_load_incoming_0 & ~will_fire_stad_incoming_0;	// lsu.scala:441:63, :534:63, :538:{31,34}
  wire              _will_fire_sta_incoming_0_will_fire_T_6 =
    ~can_fire_load_incoming_0 & ~will_fire_stad_incoming_0;	// lsu.scala:441:63, :534:63, :539:{31,34}
  wire              will_fire_sta_incoming_0 =
    _can_fire_sta_incoming_T & ~io_core_exe_0_req_bits_uop_ctrl_is_std
    & _will_fire_sta_incoming_0_will_fire_T_2 & _will_fire_sta_incoming_0_will_fire_T_6
    & ~will_fire_stad_incoming_0;	// lsu.scala:444:63, :449:66, :534:63, :536:61, :537:35, :538:31, :539:31
  wire              _will_fire_sfence_0_will_fire_T_2 =
    _will_fire_sta_incoming_0_will_fire_T_2 & ~will_fire_sta_incoming_0;	// lsu.scala:536:61, :538:{31,34}
  wire              _will_fire_release_0_will_fire_T_6 =
    _will_fire_sta_incoming_0_will_fire_T_6 & ~will_fire_sta_incoming_0;	// lsu.scala:536:61, :539:{31,34}
  wire              _will_fire_std_incoming_0_will_fire_T_14 =
    ~will_fire_stad_incoming_0 & ~will_fire_sta_incoming_0;	// lsu.scala:534:63, :536:61, :541:{31,34}
  wire              will_fire_std_incoming_0 =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_ctrl_is_std
    & ~io_core_exe_0_req_bits_uop_ctrl_is_sta & _will_fire_std_incoming_0_will_fire_T_14;	// lsu.scala:453:66, :536:61, :541:31
  wire              _will_fire_sfence_0_will_fire_T_14 =
    _will_fire_std_incoming_0_will_fire_T_14 & ~will_fire_std_incoming_0;	// lsu.scala:536:61, :541:{31,34}
  wire              will_fire_sfence_0 =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_sfence_valid
    & _will_fire_sfence_0_will_fire_T_2 & _will_fire_sfence_0_will_fire_T_14;	// lsu.scala:536:61, :538:31, :541:31
  wire              _will_fire_hella_incoming_0_will_fire_T_2 =
    _will_fire_sfence_0_will_fire_T_2 & ~will_fire_sfence_0;	// lsu.scala:536:61, :538:{31,34}
  wire              will_fire_release_0 =
    io_dmem_release_valid & _will_fire_release_0_will_fire_T_6;	// lsu.scala:534:63, :539:31
  wire              _will_fire_load_retry_0_will_fire_T_6 =
    _will_fire_release_0_will_fire_T_6 & ~will_fire_release_0;	// lsu.scala:534:63, :539:{31,34}
  wire              will_fire_hella_incoming_0 =
    (|hella_state) & _GEN_1 & _will_fire_hella_incoming_0_will_fire_T_2
    & ~can_fire_load_incoming_0;	// lsu.scala:242:38, :441:63, :535:65, :536:35, :538:31, :593:24, :803:26
  wire              _will_fire_load_retry_0_will_fire_T_2 =
    _will_fire_hella_incoming_0_will_fire_T_2 & ~will_fire_hella_incoming_0;	// lsu.scala:535:65, :538:{31,34}
  wire              _will_fire_hella_wakeup_0_will_fire_T_10 =
    ~can_fire_load_incoming_0 & ~will_fire_hella_incoming_0;	// lsu.scala:441:63, :535:65, :540:{31,34}
  wire              will_fire_hella_wakeup_0 =
    _GEN & _GEN_0 & _will_fire_hella_wakeup_0_will_fire_T_10;	// lsu.scala:535:65, :540:31, :820:26, :1527:34, :1533:38, :1550:43, :1553:38, :1560:40, :1576:42
  wire              _will_fire_load_retry_0_will_fire_T_10 =
    _will_fire_hella_wakeup_0_will_fire_T_10 & ~will_fire_hella_wakeup_0;	// lsu.scala:535:65, :540:{31,34}
  wire              will_fire_load_retry_0 =
    _GEN_99[ldq_retry_idx] & _GEN_113[ldq_retry_idx] & _GEN_200[ldq_retry_idx]
    & ~_GEN_202[ldq_retry_idx] & ~_GEN_203[ldq_retry_idx] & can_fire_load_retry_REG
    & ~store_needs_order & ~_GEN_201[ldq_retry_idx]
    & _will_fire_load_retry_0_will_fire_T_2 & _will_fire_load_retry_0_will_fire_T_6
    & _will_fire_load_retry_0_will_fire_T_10;	// lsu.scala:264:49, :305:44, :415:30, :465:79, :468:33, :469:33, :470:40, :471:33, :473:33, :535:65, :538:31, :539:31, :540:31, :1495:3, :1496:64
  wire              _will_fire_sta_retry_0_will_fire_T_2 =
    _will_fire_load_retry_0_will_fire_T_2 & ~will_fire_load_retry_0;	// lsu.scala:535:65, :538:{31,34}
  wire              _will_fire_sta_retry_0_will_fire_T_6 =
    _will_fire_load_retry_0_will_fire_T_6 & ~will_fire_load_retry_0;	// lsu.scala:535:65, :539:{31,34}
  wire              _will_fire_load_wakeup_0_will_fire_T_10 =
    _will_fire_load_retry_0_will_fire_T_10 & ~will_fire_load_retry_0;	// lsu.scala:535:65, :540:{31,34}
  wire              will_fire_sta_retry_0 =
    _GEN_204 & _GEN_87[stq_retry_idx] & _GEN_90[stq_retry_idx] & can_fire_sta_retry_REG
    & _will_fire_sta_retry_0_will_fire_T_2 & _will_fire_sta_retry_0_will_fire_T_6
    & _will_fire_sfence_0_will_fire_T_14 & ~will_fire_sfence_0;	// lsu.scala:224:42, :422:30, :478:79, :482:41, :536:61, :538:31, :539:31, :541:{31,34}
  assign _will_fire_store_commit_0_T_2 =
    _will_fire_sta_retry_0_will_fire_T_2 & ~will_fire_sta_retry_0;	// lsu.scala:536:61, :538:{31,34}
  wire              will_fire_load_wakeup_0 =
    _GEN_99[ldq_wakeup_idx] & _GEN_113[ldq_wakeup_idx] & ~_GEN_214[ldq_wakeup_idx]
    & ~_GEN_211 & ~_GEN_213 & ~_GEN_201[ldq_wakeup_idx] & ~_GEN_202[ldq_wakeup_idx]
    & ~_GEN_203[ldq_wakeup_idx] & ~store_needs_order & ~block_load_wakeup
    & (~_GEN_212[ldq_wakeup_idx] | io_core_commit_load_at_rob_head
       & ldq_head == ldq_wakeup_idx & mem_ldq_wakeup_e_out_bits_st_dep_mask == 24'h0)
    & _will_fire_sta_retry_0_will_fire_T_6 & ~will_fire_sta_retry_0
    & _will_fire_load_wakeup_0_will_fire_T_10;	// lsu.scala:215:29, :259:32, :264:49, :305:44, :430:31, :465:79, :468:33, :469:33, :471:33, :502:88, :504:31, :505:31, :506:31, :507:31, :508:31, :509:31, :511:31, :513:{32,71}, :514:{84,103}, :515:112, :535:65, :536:61, :539:{31,34}, :540:31, :1199:80, :1210:43, :1211:25, :1495:3, :1496:64
  wire              will_fire_store_commit_0 =
    can_fire_store_commit_0 & _will_fire_load_wakeup_0_will_fire_T_10
    & ~will_fire_load_wakeup_0;	// lsu.scala:493:79, :535:65, :540:{31,34}
  wire              _exe_cmd_T = can_fire_load_incoming_0 | will_fire_stad_incoming_0;	// lsu.scala:441:63, :534:63, :567:63
  wire              _GEN_215 = _exe_cmd_T | will_fire_sta_incoming_0;	// lsu.scala:536:61, :567:{63,93}
  wire              _GEN_216 = ldq_wakeup_idx == 5'h0;	// lsu.scala:430:31, :570:49
  wire              _GEN_217 = ldq_wakeup_idx == 5'h1;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_218 = ldq_wakeup_idx == 5'h2;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_219 = ldq_wakeup_idx == 5'h3;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_220 = ldq_wakeup_idx == 5'h4;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_221 = ldq_wakeup_idx == 5'h5;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_222 = ldq_wakeup_idx == 5'h6;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_223 = ldq_wakeup_idx == 5'h7;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_224 = ldq_wakeup_idx == 5'h8;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_225 = ldq_wakeup_idx == 5'h9;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_226 = ldq_wakeup_idx == 5'hA;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_227 = ldq_wakeup_idx == 5'hB;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_228 = ldq_wakeup_idx == 5'hC;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_229 = ldq_wakeup_idx == 5'hD;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_230 = ldq_wakeup_idx == 5'hE;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_231 = ldq_wakeup_idx == 5'hF;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_232 = ldq_wakeup_idx == 5'h10;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_233 = ldq_wakeup_idx == 5'h11;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_234 = ldq_wakeup_idx == 5'h12;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_235 = ldq_wakeup_idx == 5'h13;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_236 = ldq_wakeup_idx == 5'h14;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_237 = ldq_wakeup_idx == 5'h15;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_238 = ldq_wakeup_idx == 5'h16;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_239 = ldq_wakeup_idx == 5'h17;	// lsu.scala:430:31, :570:49, util.scala:205:25
  wire              _GEN_240 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h0;	// lsu.scala:572:52
  wire              _GEN_241 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h1;	// lsu.scala:305:44, :572:52
  wire              _GEN_242 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h2;	// lsu.scala:305:44, :572:52
  wire              _GEN_243 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h3;	// lsu.scala:305:44, :572:52
  wire              _GEN_244 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h4;	// lsu.scala:305:44, :572:52
  wire              _GEN_245 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h5;	// lsu.scala:305:44, :572:52
  wire              _GEN_246 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h6;	// lsu.scala:305:44, :572:52
  wire              _GEN_247 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h7;	// lsu.scala:305:44, :572:52
  wire              _GEN_248 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h8;	// lsu.scala:305:44, :572:52
  wire              _GEN_249 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h9;	// lsu.scala:305:44, :572:52
  wire              _GEN_250 = io_core_exe_0_req_bits_uop_ldq_idx == 5'hA;	// lsu.scala:305:44, :572:52
  wire              _GEN_251 = io_core_exe_0_req_bits_uop_ldq_idx == 5'hB;	// lsu.scala:305:44, :572:52
  wire              _GEN_252 = io_core_exe_0_req_bits_uop_ldq_idx == 5'hC;	// lsu.scala:305:44, :572:52
  wire              _GEN_253 = io_core_exe_0_req_bits_uop_ldq_idx == 5'hD;	// lsu.scala:305:44, :572:52
  wire              _GEN_254 = io_core_exe_0_req_bits_uop_ldq_idx == 5'hE;	// lsu.scala:305:44, :572:52
  wire              _GEN_255 = io_core_exe_0_req_bits_uop_ldq_idx == 5'hF;	// lsu.scala:305:44, :572:52
  wire              _GEN_256 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h10;	// lsu.scala:305:44, :572:52
  wire              _GEN_257 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h11;	// lsu.scala:305:44, :572:52
  wire              _GEN_258 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h12;	// lsu.scala:305:44, :572:52
  wire              _GEN_259 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h13;	// lsu.scala:305:44, :572:52
  wire              _GEN_260 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h14;	// lsu.scala:305:44, :572:52
  wire              _GEN_261 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h15;	// lsu.scala:305:44, :572:52
  wire              _GEN_262 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h16;	// lsu.scala:305:44, :572:52
  wire              _GEN_263 = io_core_exe_0_req_bits_uop_ldq_idx == 5'h17;	// lsu.scala:572:52, util.scala:205:25
  wire              _GEN_264 = ldq_retry_idx == 5'h0;	// lsu.scala:415:30, :574:49
  wire              _GEN_265 = will_fire_load_retry_0 & _GEN_264;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_266 = ldq_retry_idx == 5'h1;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_267 = will_fire_load_retry_0 & _GEN_266;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_268 = ldq_retry_idx == 5'h2;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_269 = will_fire_load_retry_0 & _GEN_268;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_270 = ldq_retry_idx == 5'h3;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_271 = will_fire_load_retry_0 & _GEN_270;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_272 = ldq_retry_idx == 5'h4;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_273 = will_fire_load_retry_0 & _GEN_272;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_274 = ldq_retry_idx == 5'h5;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_275 = will_fire_load_retry_0 & _GEN_274;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_276 = ldq_retry_idx == 5'h6;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_277 = will_fire_load_retry_0 & _GEN_276;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_278 = ldq_retry_idx == 5'h7;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_279 = will_fire_load_retry_0 & _GEN_278;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_280 = ldq_retry_idx == 5'h8;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_281 = will_fire_load_retry_0 & _GEN_280;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_282 = ldq_retry_idx == 5'h9;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_283 = will_fire_load_retry_0 & _GEN_282;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_284 = ldq_retry_idx == 5'hA;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_285 = will_fire_load_retry_0 & _GEN_284;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_286 = ldq_retry_idx == 5'hB;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_287 = will_fire_load_retry_0 & _GEN_286;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_288 = ldq_retry_idx == 5'hC;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_289 = will_fire_load_retry_0 & _GEN_288;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_290 = ldq_retry_idx == 5'hD;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_291 = will_fire_load_retry_0 & _GEN_290;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_292 = ldq_retry_idx == 5'hE;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_293 = will_fire_load_retry_0 & _GEN_292;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_294 = ldq_retry_idx == 5'hF;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_295 = will_fire_load_retry_0 & _GEN_294;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_296 = ldq_retry_idx == 5'h10;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_297 = will_fire_load_retry_0 & _GEN_296;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_298 = ldq_retry_idx == 5'h11;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_299 = will_fire_load_retry_0 & _GEN_298;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_300 = ldq_retry_idx == 5'h12;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_301 = will_fire_load_retry_0 & _GEN_300;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_302 = ldq_retry_idx == 5'h13;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_303 = will_fire_load_retry_0 & _GEN_302;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_304 = ldq_retry_idx == 5'h14;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_305 = will_fire_load_retry_0 & _GEN_304;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_306 = ldq_retry_idx == 5'h15;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_307 = will_fire_load_retry_0 & _GEN_306;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_308 = ldq_retry_idx == 5'h16;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_309 = will_fire_load_retry_0 & _GEN_308;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_310 = ldq_retry_idx == 5'h17;	// lsu.scala:415:30, :574:49, util.scala:205:25
  wire              _GEN_311 = will_fire_load_retry_0 & _GEN_310;	// lsu.scala:535:65, :573:43, :574:49
  wire              _exe_tlb_uop_T_2 =
    _exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0;	// lsu.scala:536:61, :567:63, :599:53
  wire              _exe_tlb_uop_T_4_uses_ldq =
    will_fire_sta_retry_0 & _GEN_63[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79, :536:61, :602:24
  wire              _exe_tlb_uop_T_4_uses_stq =
    will_fire_sta_retry_0 & _GEN_64[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79, :536:61, :602:24
  wire              exe_tlb_uop_0_ctrl_is_load =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_ctrl_is_load
      : will_fire_load_retry_0
          ? _GEN_130[ldq_retry_idx]
          : will_fire_sta_retry_0 & _GEN_18[stq_retry_idx];	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire              exe_tlb_uop_0_ctrl_is_sta =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_ctrl_is_sta
      : will_fire_load_retry_0
          ? _GEN_131[ldq_retry_idx]
          : will_fire_sta_retry_0 & _GEN_19[stq_retry_idx];	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire [15:0]       exe_tlb_uop_0_br_mask =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_br_mask
      : will_fire_load_retry_0 ? _GEN_140 : will_fire_sta_retry_0 ? _GEN_205 : 16'h0;	// lsu.scala:465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire [4:0]        exe_tlb_uop_0_mem_cmd =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_mem_cmd
      : will_fire_load_retry_0
          ? _GEN_167[ldq_retry_idx]
          : will_fire_sta_retry_0 ? _GEN_54[stq_retry_idx] : 5'h0;	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire [1:0]        exe_tlb_uop_0_mem_size =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_mem_size
      : will_fire_load_retry_0
          ? mem_ldq_retry_e_out_bits_uop_mem_size
          : will_fire_sta_retry_0 ? mem_stq_retry_e_out_bits_uop_mem_size : 2'h0;	// lsu.scala:465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire              exe_tlb_uop_0_is_fence =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_is_fence
      : will_fire_load_retry_0
          ? _GEN_169[ldq_retry_idx]
          : will_fire_sta_retry_0 & _GEN_58[stq_retry_idx];	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire              _mem_xcpt_uops_WIRE_0_uses_ldq =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_uses_ldq
      : will_fire_load_retry_0 ? _GEN_173 : _exe_tlb_uop_T_4_uses_ldq;	// lsu.scala:465:79, :535:65, :597:24, :599:53, :601:24, :602:24
  wire              _mem_xcpt_uops_WIRE_0_uses_stq =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_uses_stq
      : will_fire_load_retry_0 ? _GEN_175 : _exe_tlb_uop_T_4_uses_stq;	// lsu.scala:465:79, :535:65, :597:24, :599:53, :601:24, :602:24
  wire              _exe_tlb_vaddr_T_1 = _exe_cmd_T | will_fire_sta_incoming_0;	// lsu.scala:536:61, :567:63, :608:53
  wire [39:0]       _GEN_312 = {1'h0, io_core_exe_0_req_bits_sfence_bits_addr};	// lsu.scala:249:20, :610:24, :708:86
  wire [39:0]       exe_tlb_vaddr_0 =
    _exe_tlb_vaddr_T_1
      ? io_core_exe_0_req_bits_addr
      : will_fire_sfence_0
          ? _GEN_312
          : will_fire_load_retry_0
              ? _GEN_199
              : will_fire_sta_retry_0
                  ? _GEN_208
                  : will_fire_hella_incoming_0 ? hella_req_addr : 40'h0;	// lsu.scala:243:34, :465:79, :478:79, :535:65, :536:61, :607:24, :608:53, :610:24, :611:24, :612:24, :613:24
  wire              _stq_idx_T = will_fire_sta_incoming_0 | will_fire_stad_incoming_0;	// lsu.scala:534:63, :536:61, :660:56
  reg  [15:0]       mem_xcpt_uops_0_br_mask;	// lsu.scala:671:32
  reg  [6:0]        mem_xcpt_uops_0_rob_idx;	// lsu.scala:671:32
  reg  [4:0]        mem_xcpt_uops_0_ldq_idx;	// lsu.scala:671:32
  reg  [4:0]        mem_xcpt_uops_0_stq_idx;	// lsu.scala:671:32
  reg               mem_xcpt_uops_0_uses_ldq;	// lsu.scala:671:32
  reg               mem_xcpt_uops_0_uses_stq;	// lsu.scala:671:32
  reg  [3:0]        mem_xcpt_causes_0;	// lsu.scala:672:32
  reg  [39:0]       mem_xcpt_vaddrs_0;	// lsu.scala:679:32
  wire              exe_tlb_miss_0 =
    ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_miss;	// lsu.scala:249:20, :538:31, :576:25, :708:58
  wire [31:0]       exe_tlb_paddr_0 =
    {_dtlb_io_resp_0_paddr[31:12], exe_tlb_vaddr_0[11:0]};	// Cat.scala:30:58, lsu.scala:249:20, :607:24, :709:62, :710:57
  reg               REG;	// lsu.scala:718:21
  wire [39:0]       _GEN_313 =
    {8'h0, _dtlb_io_resp_0_paddr[31:12], exe_tlb_vaddr_0[11:0]};	// lsu.scala:249:20, :260:63, :607:24, :709:62, :710:57, :768:30
  wire [3:0][63:0]  _GEN_314 =
    {{_GEN_93},
     {{2{_GEN_93[31:0]}}},
     {{2{{2{_GEN_93[15:0]}}}}},
     {{2{{2{{2{_GEN_93[7:0]}}}}}}}};	// AMOALU.scala:26:{13,19,66}, Cat.scala:30:58, lsu.scala:224:42
  wire              _GEN_315 = can_fire_load_incoming_0 | will_fire_load_retry_0;	// lsu.scala:220:29, :441:63, :535:65, :766:39, :773:43, :780:45
  assign _GEN_1 = hella_state == 3'h1;	// lsu.scala:242:38, :803:26
  wire              _GEN_316 = will_fire_store_commit_0 | will_fire_load_wakeup_0;	// lsu.scala:245:34, :535:65, :780:45, :794:44, :802:47
  assign _GEN_0 = hella_state == 3'h5;	// lsu.scala:242:38, :820:26, util.scala:351:72
  wire              dmem_req_0_valid =
    can_fire_load_incoming_0
      ? ~exe_tlb_miss_0 & _dtlb_io_resp_0_cacheable
      : will_fire_load_retry_0
          ? ~exe_tlb_miss_0 & _dtlb_io_resp_0_cacheable
          : _GEN_316
            | (will_fire_hella_incoming_0
                 ? ~io_hellacache_s1_kill & (~exe_tlb_miss_0 | hella_req_phys)
                 : will_fire_hella_wakeup_0);	// lsu.scala:243:34, :245:34, :249:20, :441:63, :535:65, :708:58, :766:39, :767:{30,33,50}, :773:43, :774:{30,33,50}, :780:45, :781:33, :794:44, :795:30, :802:47, :805:{39,42,65,69,86}, :819:5
  wire [39:0]       _GEN_317 = {8'h0, hella_paddr};	// lsu.scala:245:34, :260:63, :822:39
  wire              _GEN_318 = can_fire_load_incoming_0 | will_fire_load_retry_0;	// lsu.scala:441:63, :535:65, :766:39, :768:30, :773:43
  wire [3:0][63:0]  _GEN_319 =
    {{hella_data_data},
     {{2{hella_data_data[31:0]}}},
     {{2{{2{hella_data_data[15:0]}}}}},
     {{2{{2{{2{hella_data_data[7:0]}}}}}}}};	// AMOALU.scala:26:{13,19,66}, Cat.scala:30:58, lsu.scala:244:34
  wire              _GEN_320 = will_fire_hella_incoming_0 | will_fire_hella_wakeup_0;	// lsu.scala:535:65, :759:28, :802:47, :811:39, :819:5, :827:39
  wire              _GEN_321 = _stq_idx_T | will_fire_sta_retry_0;	// lsu.scala:536:61, :660:56, :848:67
  wire              _io_core_fp_stdata_ready_output =
    ~will_fire_std_incoming_0 & ~will_fire_stad_incoming_0;	// lsu.scala:534:63, :536:61, :866:{34,61,64}
  wire              fp_stdata_fire =
    _io_core_fp_stdata_ready_output & io_core_fp_stdata_valid;	// Decoupled.scala:40:37, lsu.scala:866:61
  wire              _stq_bits_data_bits_T =
    will_fire_std_incoming_0 | will_fire_stad_incoming_0;	// lsu.scala:534:63, :536:61, :868:37
  wire              _GEN_322 = _stq_bits_data_bits_T | fp_stdata_fire;	// Decoupled.scala:40:37, lsu.scala:868:{37,67}
  wire [4:0]        sidx =
    _stq_bits_data_bits_T
      ? io_core_exe_0_req_bits_uop_stq_idx
      : io_core_fp_stdata_bits_uop_stq_idx;	// lsu.scala:868:37, :870:21
  reg               fired_load_incoming_REG;	// lsu.scala:894:51
  reg               fired_stad_incoming_REG;	// lsu.scala:895:51
  reg               fired_sta_incoming_REG;	// lsu.scala:896:51
  reg               fired_std_incoming_REG;	// lsu.scala:897:51
  reg               fired_stdf_incoming;	// lsu.scala:898:37
  reg               fired_sfence_0;	// lsu.scala:899:37
  reg               fired_release_0;	// lsu.scala:900:37
  reg               fired_load_retry_REG;	// lsu.scala:901:51
  reg               fired_sta_retry_REG;	// lsu.scala:902:51
  reg               fired_load_wakeup_REG;	// lsu.scala:904:51
  reg  [15:0]       mem_incoming_uop_0_br_mask;	// lsu.scala:908:37
  reg  [6:0]        mem_incoming_uop_0_rob_idx;	// lsu.scala:908:37
  reg  [4:0]        mem_incoming_uop_0_ldq_idx;	// lsu.scala:908:37
  reg  [4:0]        mem_incoming_uop_0_stq_idx;	// lsu.scala:908:37
  reg  [6:0]        mem_incoming_uop_0_pdst;	// lsu.scala:908:37
  reg               mem_incoming_uop_0_fp_val;	// lsu.scala:908:37
  reg  [15:0]       mem_ldq_incoming_e_0_bits_uop_br_mask;	// lsu.scala:909:37
  reg  [4:0]        mem_ldq_incoming_e_0_bits_uop_stq_idx;	// lsu.scala:909:37
  reg  [1:0]        mem_ldq_incoming_e_0_bits_uop_mem_size;	// lsu.scala:909:37
  reg  [23:0]       mem_ldq_incoming_e_0_bits_st_dep_mask;	// lsu.scala:909:37
  reg               mem_stq_incoming_e_0_valid;	// lsu.scala:910:37
  reg  [15:0]       mem_stq_incoming_e_0_bits_uop_br_mask;	// lsu.scala:910:37
  reg  [6:0]        mem_stq_incoming_e_0_bits_uop_rob_idx;	// lsu.scala:910:37
  reg  [4:0]        mem_stq_incoming_e_0_bits_uop_stq_idx;	// lsu.scala:910:37
  reg  [1:0]        mem_stq_incoming_e_0_bits_uop_mem_size;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_uop_is_amo;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_addr_valid;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_addr_is_virtual;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_data_valid;	// lsu.scala:910:37
  reg  [15:0]       mem_ldq_wakeup_e_bits_uop_br_mask;	// lsu.scala:911:37
  reg  [4:0]        mem_ldq_wakeup_e_bits_uop_stq_idx;	// lsu.scala:911:37
  reg  [1:0]        mem_ldq_wakeup_e_bits_uop_mem_size;	// lsu.scala:911:37
  reg  [23:0]       mem_ldq_wakeup_e_bits_st_dep_mask;	// lsu.scala:911:37
  reg  [15:0]       mem_ldq_retry_e_bits_uop_br_mask;	// lsu.scala:912:37
  reg  [4:0]        mem_ldq_retry_e_bits_uop_stq_idx;	// lsu.scala:912:37
  reg  [1:0]        mem_ldq_retry_e_bits_uop_mem_size;	// lsu.scala:912:37
  reg  [23:0]       mem_ldq_retry_e_bits_st_dep_mask;	// lsu.scala:912:37
  reg               mem_stq_retry_e_valid;	// lsu.scala:913:37
  reg  [15:0]       mem_stq_retry_e_bits_uop_br_mask;	// lsu.scala:913:37
  reg  [6:0]        mem_stq_retry_e_bits_uop_rob_idx;	// lsu.scala:913:37
  reg  [4:0]        mem_stq_retry_e_bits_uop_stq_idx;	// lsu.scala:913:37
  reg  [1:0]        mem_stq_retry_e_bits_uop_mem_size;	// lsu.scala:913:37
  reg               mem_stq_retry_e_bits_uop_is_amo;	// lsu.scala:913:37
  reg               mem_stq_retry_e_bits_data_valid;	// lsu.scala:913:37
  wire [23:0]       lcam_st_dep_mask_0 =
    fired_load_incoming_REG
      ? mem_ldq_incoming_e_0_bits_st_dep_mask
      : fired_load_retry_REG
          ? mem_ldq_retry_e_bits_st_dep_mask
          : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_st_dep_mask : 24'h0;	// lsu.scala:259:32, :894:51, :901:51, :904:51, :909:37, :911:37, :912:37, :915:33, :916:33, :917:33
  wire              _lcam_stq_idx_T = fired_stad_incoming_REG | fired_sta_incoming_REG;	// lsu.scala:895:51, :896:51, :919:57
  reg  [15:0]       mem_stdf_uop_br_mask;	// lsu.scala:922:37
  reg  [6:0]        mem_stdf_uop_rob_idx;	// lsu.scala:922:37
  reg  [4:0]        mem_stdf_uop_stq_idx;	// lsu.scala:922:37
  reg               mem_tlb_miss_0;	// lsu.scala:925:41
  reg               mem_tlb_uncacheable_0;	// lsu.scala:926:41
  reg  [39:0]       mem_paddr_0;	// lsu.scala:927:41
  reg               clr_bsy_valid_0;	// lsu.scala:930:32
  reg  [6:0]        clr_bsy_rob_idx_0;	// lsu.scala:931:28
  reg  [15:0]       clr_bsy_brmask_0;	// lsu.scala:932:28
  reg               io_core_clr_bsy_0_valid_REG;	// lsu.scala:979:62
  reg               io_core_clr_bsy_0_valid_REG_1;	// lsu.scala:979:101
  reg               io_core_clr_bsy_0_valid_REG_2;	// lsu.scala:979:93
  reg               stdf_clr_bsy_valid;	// lsu.scala:983:37
  reg  [6:0]        stdf_clr_bsy_rob_idx;	// lsu.scala:984:33
  reg  [15:0]       stdf_clr_bsy_brmask;	// lsu.scala:985:33
  reg               io_core_clr_bsy_1_valid_REG;	// lsu.scala:1004:67
  reg               io_core_clr_bsy_1_valid_REG_1;	// lsu.scala:1004:106
  reg               io_core_clr_bsy_1_valid_REG_2;	// lsu.scala:1004:98
  wire              do_st_search_0 =
    (_lcam_stq_idx_T | fired_sta_retry_REG) & ~mem_tlb_miss_0;	// lsu.scala:902:51, :919:57, :925:41, :1014:{85,108,111}
  wire              _can_forward_T = fired_load_incoming_REG | fired_load_retry_REG;	// lsu.scala:894:51, :901:51, :1016:61
  wire              do_ld_search_0 =
    _can_forward_T & ~mem_tlb_miss_0 | fired_load_wakeup_REG;	// lsu.scala:904:51, :925:41, :1014:111, :1016:{61,85,106}
  wire              _lcam_addr_T_1 = _lcam_stq_idx_T | fired_sta_retry_REG;	// lsu.scala:902:51, :919:57, :1025:86
  reg  [31:0]       lcam_addr_REG;	// lsu.scala:1026:45
  reg  [31:0]       lcam_addr_REG_1;	// lsu.scala:1027:67
  wire [39:0]       _GEN_323 = {8'h0, lcam_addr_REG_1};	// lsu.scala:260:63, :1027:{41,67}
  wire [39:0]       _GEN_324 = {8'h0, lcam_addr_REG};	// lsu.scala:260:63, :1025:37, :1026:45
  wire [39:0]       lcam_addr_0 =
    _lcam_addr_T_1 ? _GEN_324 : fired_release_0 ? _GEN_323 : mem_paddr_0;	// lsu.scala:900:37, :927:41, :1025:{37,86}, :1027:41
  wire [14:0]       _lcam_mask_mask_T_2 = 15'h1 << lcam_addr_0[2:0];	// lsu.scala:1025:37, :1663:{48,55}
  wire [14:0]       _lcam_mask_mask_T_6 = 15'h3 << {12'h0, lcam_addr_0[2:1], 1'h0};	// lsu.scala:249:20, :708:86, :1025:37, :1664:{48,56}
  wire [3:0][7:0]   _GEN_325 =
    {{8'hFF},
     {lcam_addr_0[2] ? 8'hF0 : 8'hF},
     {_lcam_mask_mask_T_6[7:0]},
     {_lcam_mask_mask_T_2[7:0]}};	// Mux.scala:98:16, lsu.scala:1025:37, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire [7:0]        lcam_mask_0 =
    _GEN_325[do_st_search_0
               ? (_lcam_stq_idx_T
                    ? mem_stq_incoming_e_0_bits_uop_mem_size
                    : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_mem_size : 2'h0)
               : do_ld_search_0
                   ? (fired_load_incoming_REG
                        ? mem_ldq_incoming_e_0_bits_uop_mem_size
                        : fired_load_retry_REG
                            ? mem_ldq_retry_e_bits_uop_mem_size
                            : fired_load_wakeup_REG
                                ? mem_ldq_wakeup_e_bits_uop_mem_size
                                : 2'h0)
                   : 2'h0];	// Mux.scala:98:16, lsu.scala:894:51, :901:51, :902:51, :904:51, :909:37, :910:37, :911:37, :912:37, :913:37, :915:33, :916:33, :917:33, :919:{33,57}, :921:33, :1014:108, :1016:106, :1029:37, :1030:37, :1663:26, :1664:26, :1665:26
  reg  [4:0]        lcam_ldq_idx_REG;	// lsu.scala:1037:58
  reg  [4:0]        lcam_ldq_idx_REG_1;	// lsu.scala:1038:58
  wire [4:0]        lcam_ldq_idx_0 =
    fired_load_incoming_REG
      ? mem_incoming_uop_0_ldq_idx
      : fired_load_wakeup_REG
          ? lcam_ldq_idx_REG
          : fired_load_retry_REG ? lcam_ldq_idx_REG_1 : 5'h0;	// lsu.scala:894:51, :901:51, :904:51, :908:37, :1036:26, :1037:{26,58}, :1038:{26,58}
  reg  [4:0]        lcam_stq_idx_REG;	// lsu.scala:1042:58
  wire [4:0]        lcam_stq_idx_0 =
    _lcam_stq_idx_T
      ? mem_incoming_uop_0_stq_idx
      : fired_sta_retry_REG ? lcam_stq_idx_REG : 5'h0;	// lsu.scala:902:51, :908:37, :919:57, :1040:26, :1042:{26,58}
  reg               s1_executing_loads_0;	// lsu.scala:1056:35
  reg               s1_executing_loads_1;	// lsu.scala:1056:35
  reg               s1_executing_loads_2;	// lsu.scala:1056:35
  reg               s1_executing_loads_3;	// lsu.scala:1056:35
  reg               s1_executing_loads_4;	// lsu.scala:1056:35
  reg               s1_executing_loads_5;	// lsu.scala:1056:35
  reg               s1_executing_loads_6;	// lsu.scala:1056:35
  reg               s1_executing_loads_7;	// lsu.scala:1056:35
  reg               s1_executing_loads_8;	// lsu.scala:1056:35
  reg               s1_executing_loads_9;	// lsu.scala:1056:35
  reg               s1_executing_loads_10;	// lsu.scala:1056:35
  reg               s1_executing_loads_11;	// lsu.scala:1056:35
  reg               s1_executing_loads_12;	// lsu.scala:1056:35
  reg               s1_executing_loads_13;	// lsu.scala:1056:35
  reg               s1_executing_loads_14;	// lsu.scala:1056:35
  reg               s1_executing_loads_15;	// lsu.scala:1056:35
  reg               s1_executing_loads_16;	// lsu.scala:1056:35
  reg               s1_executing_loads_17;	// lsu.scala:1056:35
  reg               s1_executing_loads_18;	// lsu.scala:1056:35
  reg               s1_executing_loads_19;	// lsu.scala:1056:35
  reg               s1_executing_loads_20;	// lsu.scala:1056:35
  reg               s1_executing_loads_21;	// lsu.scala:1056:35
  reg               s1_executing_loads_22;	// lsu.scala:1056:35
  reg               s1_executing_loads_23;	// lsu.scala:1056:35
  reg               wb_forward_valid_0;	// lsu.scala:1064:36
  reg  [4:0]        wb_forward_ldq_idx_0;	// lsu.scala:1065:36
  reg  [39:0]       wb_forward_ld_addr_0;	// lsu.scala:1066:36
  reg  [4:0]        wb_forward_stq_idx_0;	// lsu.scala:1067:36
  wire [14:0]       _l_mask_mask_T_2 = 15'h1 << ldq_0_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_6 = 15'h3 << {12'h0, ldq_0_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_326 =
    {{8'hFF},
     {ldq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_6[7:0]},
     {_l_mask_mask_T_2[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_0 = wb_forward_valid_0 & ~(|wb_forward_ldq_idx_0);	// lsu.scala:1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_0 =
    lcam_addr_0[39:6] == ldq_0_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_0 =
    block_addr_matches_0 & lcam_addr_0[5:3] == ldq_0_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T = _GEN_326[ldq_0_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_327 =
    fired_release_0 & ldq_0_valid & ldq_0_bits_addr_valid & block_addr_matches_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_328 = ldq_0_bits_executed | ldq_0_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_329 = _GEN_328 | l_forwarders_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_330 = {19'h0, lcam_stq_idx_0};	// lsu.scala:1040:26, :1100:38
  wire [23:0]       _GEN_331 = ldq_0_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_332 =
    do_st_search_0 & ldq_0_valid & ldq_0_bits_addr_valid & _GEN_329
    & ~ldq_0_bits_addr_is_virtual & _GEN_331[0] & dword_addr_matches_0
    & (|_mask_overlap_T);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_333 =
    do_ld_search_0 & ldq_0_valid & ldq_0_bits_addr_valid & ~ldq_0_bits_addr_is_virtual
    & dword_addr_matches_0 & (|_mask_overlap_T);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older = lcam_ldq_idx_0 < ldq_head ^ (|ldq_head);	// lsu.scala:215:29, :1036:26, util.scala:363:{64,72,78}
  reg               older_nacked_REG;	// lsu.scala:1128:57
  wire              _GEN_334 = ~_GEN_328 | nacking_loads_0 | older_nacked_REG;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_335 = _GEN_327 | _GEN_332;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG;	// lsu.scala:1131:58
  wire              _GEN_336 = (|lcam_ldq_idx_0) & _GEN_334;	// lsu.scala:764:24, :1036:26, :1125:{38,47}, :1129:{56,73}, :1131:48
  wire [14:0]       _l_mask_mask_T_17 = 15'h1 << ldq_1_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_21 = 15'h3 << {12'h0, ldq_1_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_337 =
    {{8'hFF},
     {ldq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_21[7:0]},
     {_l_mask_mask_T_17[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_1_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_1_0 =
    lcam_addr_0[39:6] == ldq_1_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_1_0 =
    block_addr_matches_1_0 & lcam_addr_0[5:3] == ldq_1_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_2 = _GEN_337[ldq_1_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_338 =
    fired_release_0 & ldq_1_valid & ldq_1_bits_addr_valid & block_addr_matches_1_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_339 = ldq_1_bits_executed | ldq_1_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_340 = _GEN_339 | l_forwarders_1_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_341 = ldq_1_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_342 =
    do_st_search_0 & ldq_1_valid & ldq_1_bits_addr_valid & _GEN_340
    & ~ldq_1_bits_addr_is_virtual & _GEN_341[0] & dword_addr_matches_1_0
    & (|_mask_overlap_T_2);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_343 =
    do_ld_search_0 & ldq_1_valid & ldq_1_bits_addr_valid & ~ldq_1_bits_addr_is_virtual
    & dword_addr_matches_1_0 & (|_mask_overlap_T_2);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_1 =
    lcam_ldq_idx_0 == 5'h0 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[4:1]));	// lsu.scala:215:29, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_344 = lcam_ldq_idx_0 != 5'h1;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_1;	// lsu.scala:1128:57
  wire              _GEN_345 = ~_GEN_339 | nacking_loads_1 | older_nacked_REG_1;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_346 = _GEN_338 | _GEN_342;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_1;	// lsu.scala:1131:58
  wire              _GEN_347 =
    _GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_32 = 15'h1 << ldq_2_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_36 = 15'h3 << {12'h0, ldq_2_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_348 =
    {{8'hFF},
     {ldq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_36[7:0]},
     {_l_mask_mask_T_32[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_2_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h2;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_2_0 =
    lcam_addr_0[39:6] == ldq_2_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_2_0 =
    block_addr_matches_2_0 & lcam_addr_0[5:3] == ldq_2_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_4 = _GEN_348[ldq_2_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_349 =
    fired_release_0 & ldq_2_valid & ldq_2_bits_addr_valid & block_addr_matches_2_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_350 = ldq_2_bits_executed | ldq_2_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_351 = _GEN_350 | l_forwarders_2_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_352 = ldq_2_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_353 =
    do_st_search_0 & ldq_2_valid & ldq_2_bits_addr_valid & _GEN_351
    & ~ldq_2_bits_addr_is_virtual & _GEN_352[0] & dword_addr_matches_2_0
    & (|_mask_overlap_T_4);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_354 =
    do_ld_search_0 & ldq_2_valid & ldq_2_bits_addr_valid & ~ldq_2_bits_addr_is_virtual
    & dword_addr_matches_2_0 & (|_mask_overlap_T_4);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_2 =
    lcam_ldq_idx_0 < 5'h2 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h2;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_355 = lcam_ldq_idx_0 != 5'h2;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_2;	// lsu.scala:1128:57
  wire              _GEN_356 = ~_GEN_350 | nacking_loads_2 | older_nacked_REG_2;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_357 = _GEN_349 | _GEN_353;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_2;	// lsu.scala:1131:58
  wire              _GEN_358 =
    _GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_47 = 15'h1 << ldq_3_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_51 = 15'h3 << {12'h0, ldq_3_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_359 =
    {{8'hFF},
     {ldq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_51[7:0]},
     {_l_mask_mask_T_47[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_3_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h3;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_3_0 =
    lcam_addr_0[39:6] == ldq_3_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_3_0 =
    block_addr_matches_3_0 & lcam_addr_0[5:3] == ldq_3_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_6 = _GEN_359[ldq_3_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_360 =
    fired_release_0 & ldq_3_valid & ldq_3_bits_addr_valid & block_addr_matches_3_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_361 = ldq_3_bits_executed | ldq_3_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_362 = _GEN_361 | l_forwarders_3_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_363 = ldq_3_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_364 =
    do_st_search_0 & ldq_3_valid & ldq_3_bits_addr_valid & _GEN_362
    & ~ldq_3_bits_addr_is_virtual & _GEN_363[0] & dword_addr_matches_3_0
    & (|_mask_overlap_T_6);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_365 =
    do_ld_search_0 & ldq_3_valid & ldq_3_bits_addr_valid & ~ldq_3_bits_addr_is_virtual
    & dword_addr_matches_3_0 & (|_mask_overlap_T_6);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_3 =
    lcam_ldq_idx_0 < 5'h3 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[4:2]));	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_366 = lcam_ldq_idx_0 != 5'h3;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_3;	// lsu.scala:1128:57
  wire              _GEN_367 = ~_GEN_361 | nacking_loads_3 | older_nacked_REG_3;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_368 = _GEN_360 | _GEN_364;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_3;	// lsu.scala:1131:58
  wire              _GEN_369 =
    _GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_62 = 15'h1 << ldq_4_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_66 = 15'h3 << {12'h0, ldq_4_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_370 =
    {{8'hFF},
     {ldq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_66[7:0]},
     {_l_mask_mask_T_62[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_4_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h4;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_4_0 =
    lcam_addr_0[39:6] == ldq_4_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_4_0 =
    block_addr_matches_4_0 & lcam_addr_0[5:3] == ldq_4_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_8 = _GEN_370[ldq_4_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_371 =
    fired_release_0 & ldq_4_valid & ldq_4_bits_addr_valid & block_addr_matches_4_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_372 = ldq_4_bits_executed | ldq_4_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_373 = _GEN_372 | l_forwarders_4_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_374 = ldq_4_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_375 =
    do_st_search_0 & ldq_4_valid & ldq_4_bits_addr_valid & _GEN_373
    & ~ldq_4_bits_addr_is_virtual & _GEN_374[0] & dword_addr_matches_4_0
    & (|_mask_overlap_T_8);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_376 =
    do_ld_search_0 & ldq_4_valid & ldq_4_bits_addr_valid & ~ldq_4_bits_addr_is_virtual
    & dword_addr_matches_4_0 & (|_mask_overlap_T_8);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_4 =
    lcam_ldq_idx_0 < 5'h4 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h4;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_377 = lcam_ldq_idx_0 != 5'h4;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_4;	// lsu.scala:1128:57
  wire              _GEN_378 = ~_GEN_372 | nacking_loads_4 | older_nacked_REG_4;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_379 = _GEN_371 | _GEN_375;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_4;	// lsu.scala:1131:58
  wire              _GEN_380 =
    _GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_77 = 15'h1 << ldq_5_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_81 = 15'h3 << {12'h0, ldq_5_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_381 =
    {{8'hFF},
     {ldq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_81[7:0]},
     {_l_mask_mask_T_77[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_5_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h5;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_5_0 =
    lcam_addr_0[39:6] == ldq_5_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_5_0 =
    block_addr_matches_5_0 & lcam_addr_0[5:3] == ldq_5_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_10 = _GEN_381[ldq_5_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_382 =
    fired_release_0 & ldq_5_valid & ldq_5_bits_addr_valid & block_addr_matches_5_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_383 = ldq_5_bits_executed | ldq_5_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_384 = _GEN_383 | l_forwarders_5_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_385 = ldq_5_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_386 =
    do_st_search_0 & ldq_5_valid & ldq_5_bits_addr_valid & _GEN_384
    & ~ldq_5_bits_addr_is_virtual & _GEN_385[0] & dword_addr_matches_5_0
    & (|_mask_overlap_T_10);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_387 =
    do_ld_search_0 & ldq_5_valid & ldq_5_bits_addr_valid & ~ldq_5_bits_addr_is_virtual
    & dword_addr_matches_5_0 & (|_mask_overlap_T_10);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_5 =
    lcam_ldq_idx_0 < 5'h5 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h5;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_388 = lcam_ldq_idx_0 != 5'h5;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_5;	// lsu.scala:1128:57
  wire              _GEN_389 = ~_GEN_383 | nacking_loads_5 | older_nacked_REG_5;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_390 = _GEN_382 | _GEN_386;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_5;	// lsu.scala:1131:58
  wire              _GEN_391 =
    _GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_92 = 15'h1 << ldq_6_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_96 = 15'h3 << {12'h0, ldq_6_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_392 =
    {{8'hFF},
     {ldq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_96[7:0]},
     {_l_mask_mask_T_92[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_6_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h6;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_6_0 =
    lcam_addr_0[39:6] == ldq_6_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_6_0 =
    block_addr_matches_6_0 & lcam_addr_0[5:3] == ldq_6_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_12 = _GEN_392[ldq_6_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_393 =
    fired_release_0 & ldq_6_valid & ldq_6_bits_addr_valid & block_addr_matches_6_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_394 = ldq_6_bits_executed | ldq_6_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_395 = _GEN_394 | l_forwarders_6_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_396 = ldq_6_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_397 =
    do_st_search_0 & ldq_6_valid & ldq_6_bits_addr_valid & _GEN_395
    & ~ldq_6_bits_addr_is_virtual & _GEN_396[0] & dword_addr_matches_6_0
    & (|_mask_overlap_T_12);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_398 =
    do_ld_search_0 & ldq_6_valid & ldq_6_bits_addr_valid & ~ldq_6_bits_addr_is_virtual
    & dword_addr_matches_6_0 & (|_mask_overlap_T_12);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_6 =
    lcam_ldq_idx_0 < 5'h6 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h6;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_399 = lcam_ldq_idx_0 != 5'h6;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_6;	// lsu.scala:1128:57
  wire              _GEN_400 = ~_GEN_394 | nacking_loads_6 | older_nacked_REG_6;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_401 = _GEN_393 | _GEN_397;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_6;	// lsu.scala:1131:58
  wire              _GEN_402 =
    _GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_107 = 15'h1 << ldq_7_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_111 =
    15'h3 << {12'h0, ldq_7_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_403 =
    {{8'hFF},
     {ldq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_111[7:0]},
     {_l_mask_mask_T_107[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_7_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h7;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_7_0 =
    lcam_addr_0[39:6] == ldq_7_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_7_0 =
    block_addr_matches_7_0 & lcam_addr_0[5:3] == ldq_7_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_14 = _GEN_403[ldq_7_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_404 =
    fired_release_0 & ldq_7_valid & ldq_7_bits_addr_valid & block_addr_matches_7_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_405 = ldq_7_bits_executed | ldq_7_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_406 = _GEN_405 | l_forwarders_7_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_407 = ldq_7_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_408 =
    do_st_search_0 & ldq_7_valid & ldq_7_bits_addr_valid & _GEN_406
    & ~ldq_7_bits_addr_is_virtual & _GEN_407[0] & dword_addr_matches_7_0
    & (|_mask_overlap_T_14);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_409 =
    do_ld_search_0 & ldq_7_valid & ldq_7_bits_addr_valid & ~ldq_7_bits_addr_is_virtual
    & dword_addr_matches_7_0 & (|_mask_overlap_T_14);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_7 =
    lcam_ldq_idx_0 < 5'h7 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[4:3]));	// lsu.scala:215:29, :305:44, :1036:26, util.scala:351:72, :363:{52,64,72,78}
  wire              _GEN_410 = lcam_ldq_idx_0 != 5'h7;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_7;	// lsu.scala:1128:57
  wire              _GEN_411 = ~_GEN_405 | nacking_loads_7 | older_nacked_REG_7;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_412 = _GEN_404 | _GEN_408;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_7;	// lsu.scala:1131:58
  wire              _GEN_413 =
    _GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_122 = 15'h1 << ldq_8_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_126 =
    15'h3 << {12'h0, ldq_8_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_414 =
    {{8'hFF},
     {ldq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_126[7:0]},
     {_l_mask_mask_T_122[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_8_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h8;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_8_0 =
    lcam_addr_0[39:6] == ldq_8_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_8_0 =
    block_addr_matches_8_0 & lcam_addr_0[5:3] == ldq_8_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_16 = _GEN_414[ldq_8_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_415 =
    fired_release_0 & ldq_8_valid & ldq_8_bits_addr_valid & block_addr_matches_8_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_416 = ldq_8_bits_executed | ldq_8_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_417 = _GEN_416 | l_forwarders_8_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_418 = ldq_8_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_419 =
    do_st_search_0 & ldq_8_valid & ldq_8_bits_addr_valid & _GEN_417
    & ~ldq_8_bits_addr_is_virtual & _GEN_418[0] & dword_addr_matches_8_0
    & (|_mask_overlap_T_16);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_420 =
    do_ld_search_0 & ldq_8_valid & ldq_8_bits_addr_valid & ~ldq_8_bits_addr_is_virtual
    & dword_addr_matches_8_0 & (|_mask_overlap_T_16);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_8 =
    lcam_ldq_idx_0 < 5'h8 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h8;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_421 = lcam_ldq_idx_0 != 5'h8;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_8;	// lsu.scala:1128:57
  wire              _GEN_422 = ~_GEN_416 | nacking_loads_8 | older_nacked_REG_8;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_423 = _GEN_415 | _GEN_419;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_8;	// lsu.scala:1131:58
  wire              _GEN_424 =
    _GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_137 = 15'h1 << ldq_9_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_141 =
    15'h3 << {12'h0, ldq_9_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_425 =
    {{8'hFF},
     {ldq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_141[7:0]},
     {_l_mask_mask_T_137[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_9_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h9;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_9_0 =
    lcam_addr_0[39:6] == ldq_9_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_9_0 =
    block_addr_matches_9_0 & lcam_addr_0[5:3] == ldq_9_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_18 = _GEN_425[ldq_9_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_426 =
    fired_release_0 & ldq_9_valid & ldq_9_bits_addr_valid & block_addr_matches_9_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_427 = ldq_9_bits_executed | ldq_9_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_428 = _GEN_427 | l_forwarders_9_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_429 = ldq_9_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_430 =
    do_st_search_0 & ldq_9_valid & ldq_9_bits_addr_valid & _GEN_428
    & ~ldq_9_bits_addr_is_virtual & _GEN_429[0] & dword_addr_matches_9_0
    & (|_mask_overlap_T_18);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_431 =
    do_ld_search_0 & ldq_9_valid & ldq_9_bits_addr_valid & ~ldq_9_bits_addr_is_virtual
    & dword_addr_matches_9_0 & (|_mask_overlap_T_18);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_9 =
    lcam_ldq_idx_0 < 5'h9 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h9;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_432 = lcam_ldq_idx_0 != 5'h9;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_9;	// lsu.scala:1128:57
  wire              _GEN_433 = ~_GEN_427 | nacking_loads_9 | older_nacked_REG_9;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_434 = _GEN_426 | _GEN_430;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_9;	// lsu.scala:1131:58
  wire              _GEN_435 =
    _GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_152 = 15'h1 << ldq_10_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_156 =
    15'h3 << {12'h0, ldq_10_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_436 =
    {{8'hFF},
     {ldq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_156[7:0]},
     {_l_mask_mask_T_152[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_10_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hA;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_10_0 =
    lcam_addr_0[39:6] == ldq_10_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_10_0 =
    block_addr_matches_10_0 & lcam_addr_0[5:3] == ldq_10_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_20 = _GEN_436[ldq_10_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_437 =
    fired_release_0 & ldq_10_valid & ldq_10_bits_addr_valid & block_addr_matches_10_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_438 = ldq_10_bits_executed | ldq_10_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_439 = _GEN_438 | l_forwarders_10_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_440 = ldq_10_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_441 =
    do_st_search_0 & ldq_10_valid & ldq_10_bits_addr_valid & _GEN_439
    & ~ldq_10_bits_addr_is_virtual & _GEN_440[0] & dword_addr_matches_10_0
    & (|_mask_overlap_T_20);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_442 =
    do_ld_search_0 & ldq_10_valid & ldq_10_bits_addr_valid & ~ldq_10_bits_addr_is_virtual
    & dword_addr_matches_10_0 & (|_mask_overlap_T_20);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_10 =
    lcam_ldq_idx_0 < 5'hA ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hA;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_443 = lcam_ldq_idx_0 != 5'hA;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_10;	// lsu.scala:1128:57
  wire              _GEN_444 = ~_GEN_438 | nacking_loads_10 | older_nacked_REG_10;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_445 = _GEN_437 | _GEN_441;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_10;	// lsu.scala:1131:58
  wire              _GEN_446 =
    _GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_167 = 15'h1 << ldq_11_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_171 =
    15'h3 << {12'h0, ldq_11_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_447 =
    {{8'hFF},
     {ldq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_171[7:0]},
     {_l_mask_mask_T_167[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_11_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hB;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_11_0 =
    lcam_addr_0[39:6] == ldq_11_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_11_0 =
    block_addr_matches_11_0 & lcam_addr_0[5:3] == ldq_11_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_22 = _GEN_447[ldq_11_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_448 =
    fired_release_0 & ldq_11_valid & ldq_11_bits_addr_valid & block_addr_matches_11_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_449 = ldq_11_bits_executed | ldq_11_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_450 = _GEN_449 | l_forwarders_11_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_451 = ldq_11_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_452 =
    do_st_search_0 & ldq_11_valid & ldq_11_bits_addr_valid & _GEN_450
    & ~ldq_11_bits_addr_is_virtual & _GEN_451[0] & dword_addr_matches_11_0
    & (|_mask_overlap_T_22);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_453 =
    do_ld_search_0 & ldq_11_valid & ldq_11_bits_addr_valid & ~ldq_11_bits_addr_is_virtual
    & dword_addr_matches_11_0 & (|_mask_overlap_T_22);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_11 =
    lcam_ldq_idx_0 < 5'hB ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hB;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_454 = lcam_ldq_idx_0 != 5'hB;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_11;	// lsu.scala:1128:57
  wire              _GEN_455 = ~_GEN_449 | nacking_loads_11 | older_nacked_REG_11;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_456 = _GEN_448 | _GEN_452;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_11;	// lsu.scala:1131:58
  wire              _GEN_457 =
    _GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_182 = 15'h1 << ldq_12_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_186 =
    15'h3 << {12'h0, ldq_12_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_458 =
    {{8'hFF},
     {ldq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_186[7:0]},
     {_l_mask_mask_T_182[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_12_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hC;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_12_0 =
    lcam_addr_0[39:6] == ldq_12_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_12_0 =
    block_addr_matches_12_0 & lcam_addr_0[5:3] == ldq_12_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_24 = _GEN_458[ldq_12_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_459 =
    fired_release_0 & ldq_12_valid & ldq_12_bits_addr_valid & block_addr_matches_12_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_460 = ldq_12_bits_executed | ldq_12_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_461 = _GEN_460 | l_forwarders_12_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_462 = ldq_12_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_463 =
    do_st_search_0 & ldq_12_valid & ldq_12_bits_addr_valid & _GEN_461
    & ~ldq_12_bits_addr_is_virtual & _GEN_462[0] & dword_addr_matches_12_0
    & (|_mask_overlap_T_24);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_464 =
    do_ld_search_0 & ldq_12_valid & ldq_12_bits_addr_valid & ~ldq_12_bits_addr_is_virtual
    & dword_addr_matches_12_0 & (|_mask_overlap_T_24);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_12 =
    lcam_ldq_idx_0 < 5'hC ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hC;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_465 = lcam_ldq_idx_0 != 5'hC;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_12;	// lsu.scala:1128:57
  wire              _GEN_466 = ~_GEN_460 | nacking_loads_12 | older_nacked_REG_12;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_467 = _GEN_459 | _GEN_463;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_12;	// lsu.scala:1131:58
  wire              _GEN_468 =
    _GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_197 = 15'h1 << ldq_13_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_201 =
    15'h3 << {12'h0, ldq_13_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_469 =
    {{8'hFF},
     {ldq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_201[7:0]},
     {_l_mask_mask_T_197[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_13_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hD;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_13_0 =
    lcam_addr_0[39:6] == ldq_13_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_13_0 =
    block_addr_matches_13_0 & lcam_addr_0[5:3] == ldq_13_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_26 = _GEN_469[ldq_13_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_470 =
    fired_release_0 & ldq_13_valid & ldq_13_bits_addr_valid & block_addr_matches_13_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_471 = ldq_13_bits_executed | ldq_13_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_472 = _GEN_471 | l_forwarders_13_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_473 = ldq_13_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_474 =
    do_st_search_0 & ldq_13_valid & ldq_13_bits_addr_valid & _GEN_472
    & ~ldq_13_bits_addr_is_virtual & _GEN_473[0] & dword_addr_matches_13_0
    & (|_mask_overlap_T_26);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_475 =
    do_ld_search_0 & ldq_13_valid & ldq_13_bits_addr_valid & ~ldq_13_bits_addr_is_virtual
    & dword_addr_matches_13_0 & (|_mask_overlap_T_26);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_13 =
    lcam_ldq_idx_0 < 5'hD ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hD;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_476 = lcam_ldq_idx_0 != 5'hD;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_13;	// lsu.scala:1128:57
  wire              _GEN_477 = ~_GEN_471 | nacking_loads_13 | older_nacked_REG_13;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_478 = _GEN_470 | _GEN_474;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_13;	// lsu.scala:1131:58
  wire              _GEN_479 =
    _GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_212 = 15'h1 << ldq_14_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_216 =
    15'h3 << {12'h0, ldq_14_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_480 =
    {{8'hFF},
     {ldq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_216[7:0]},
     {_l_mask_mask_T_212[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_14_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hE;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_14_0 =
    lcam_addr_0[39:6] == ldq_14_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_14_0 =
    block_addr_matches_14_0 & lcam_addr_0[5:3] == ldq_14_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_28 = _GEN_480[ldq_14_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_481 =
    fired_release_0 & ldq_14_valid & ldq_14_bits_addr_valid & block_addr_matches_14_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_482 = ldq_14_bits_executed | ldq_14_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_483 = _GEN_482 | l_forwarders_14_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_484 = ldq_14_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_485 =
    do_st_search_0 & ldq_14_valid & ldq_14_bits_addr_valid & _GEN_483
    & ~ldq_14_bits_addr_is_virtual & _GEN_484[0] & dword_addr_matches_14_0
    & (|_mask_overlap_T_28);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_486 =
    do_ld_search_0 & ldq_14_valid & ldq_14_bits_addr_valid & ~ldq_14_bits_addr_is_virtual
    & dword_addr_matches_14_0 & (|_mask_overlap_T_28);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_14 =
    lcam_ldq_idx_0 < 5'hE ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hE;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_487 = lcam_ldq_idx_0 != 5'hE;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_14;	// lsu.scala:1128:57
  wire              _GEN_488 = ~_GEN_482 | nacking_loads_14 | older_nacked_REG_14;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_489 = _GEN_481 | _GEN_485;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_14;	// lsu.scala:1131:58
  wire              _GEN_490 =
    _GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_227 = 15'h1 << ldq_15_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_231 =
    15'h3 << {12'h0, ldq_15_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_491 =
    {{8'hFF},
     {ldq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_231[7:0]},
     {_l_mask_mask_T_227[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_15_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hF;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_15_0 =
    lcam_addr_0[39:6] == ldq_15_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_15_0 =
    block_addr_matches_15_0 & lcam_addr_0[5:3] == ldq_15_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_30 = _GEN_491[ldq_15_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_492 =
    fired_release_0 & ldq_15_valid & ldq_15_bits_addr_valid & block_addr_matches_15_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_493 = ldq_15_bits_executed | ldq_15_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_494 = _GEN_493 | l_forwarders_15_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_495 = ldq_15_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_496 =
    do_st_search_0 & ldq_15_valid & ldq_15_bits_addr_valid & _GEN_494
    & ~ldq_15_bits_addr_is_virtual & _GEN_495[0] & dword_addr_matches_15_0
    & (|_mask_overlap_T_30);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_497 =
    do_ld_search_0 & ldq_15_valid & ldq_15_bits_addr_valid & ~ldq_15_bits_addr_is_virtual
    & dword_addr_matches_15_0 & (|_mask_overlap_T_30);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_15 =
    lcam_ldq_idx_0 < 5'hF ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head[4];	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_498 = lcam_ldq_idx_0 != 5'hF;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_15;	// lsu.scala:1128:57
  wire              _GEN_499 = ~_GEN_493 | nacking_loads_15 | older_nacked_REG_15;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_500 = _GEN_492 | _GEN_496;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_15;	// lsu.scala:1131:58
  wire              _GEN_501 =
    _GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_242 = 15'h1 << ldq_16_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_246 =
    15'h3 << {12'h0, ldq_16_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_502 =
    {{8'hFF},
     {ldq_16_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_246[7:0]},
     {_l_mask_mask_T_242[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_16_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h10;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_16_0 =
    lcam_addr_0[39:6] == ldq_16_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_16_0 =
    block_addr_matches_16_0 & lcam_addr_0[5:3] == ldq_16_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_32 = _GEN_502[ldq_16_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_503 =
    fired_release_0 & ldq_16_valid & ldq_16_bits_addr_valid & block_addr_matches_16_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_504 = ldq_16_bits_executed | ldq_16_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_505 = _GEN_504 | l_forwarders_16_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_506 = ldq_16_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_507 =
    do_st_search_0 & ldq_16_valid & ldq_16_bits_addr_valid & _GEN_505
    & ~ldq_16_bits_addr_is_virtual & _GEN_506[0] & dword_addr_matches_16_0
    & (|_mask_overlap_T_32);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_508 =
    do_ld_search_0 & ldq_16_valid & ldq_16_bits_addr_valid & ~ldq_16_bits_addr_is_virtual
    & dword_addr_matches_16_0 & (|_mask_overlap_T_32);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_16 =
    lcam_ldq_idx_0[4] ^ lcam_ldq_idx_0 >= ldq_head ^ ldq_head > 5'h10;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_509 = lcam_ldq_idx_0 != 5'h10;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_16;	// lsu.scala:1128:57
  wire              _GEN_510 = ~_GEN_504 | nacking_loads_16 | older_nacked_REG_16;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_511 = _GEN_503 | _GEN_507;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_16;	// lsu.scala:1131:58
  wire              _GEN_512 =
    _GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_257 = 15'h1 << ldq_17_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_261 =
    15'h3 << {12'h0, ldq_17_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_513 =
    {{8'hFF},
     {ldq_17_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_261[7:0]},
     {_l_mask_mask_T_257[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_17_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h11;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_17_0 =
    lcam_addr_0[39:6] == ldq_17_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_17_0 =
    block_addr_matches_17_0 & lcam_addr_0[5:3] == ldq_17_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_34 = _GEN_513[ldq_17_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_514 =
    fired_release_0 & ldq_17_valid & ldq_17_bits_addr_valid & block_addr_matches_17_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_515 = ldq_17_bits_executed | ldq_17_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_516 = _GEN_515 | l_forwarders_17_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_517 = ldq_17_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_518 =
    do_st_search_0 & ldq_17_valid & ldq_17_bits_addr_valid & _GEN_516
    & ~ldq_17_bits_addr_is_virtual & _GEN_517[0] & dword_addr_matches_17_0
    & (|_mask_overlap_T_34);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_519 =
    do_ld_search_0 & ldq_17_valid & ldq_17_bits_addr_valid & ~ldq_17_bits_addr_is_virtual
    & dword_addr_matches_17_0 & (|_mask_overlap_T_34);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_17 =
    lcam_ldq_idx_0 < 5'h11 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h11;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_520 = lcam_ldq_idx_0 != 5'h11;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_17;	// lsu.scala:1128:57
  wire              _GEN_521 = ~_GEN_515 | nacking_loads_17 | older_nacked_REG_17;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_522 = _GEN_514 | _GEN_518;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_17;	// lsu.scala:1131:58
  wire              _GEN_523 =
    _GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_272 = 15'h1 << ldq_18_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_276 =
    15'h3 << {12'h0, ldq_18_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_524 =
    {{8'hFF},
     {ldq_18_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_276[7:0]},
     {_l_mask_mask_T_272[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_18_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h12;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_18_0 =
    lcam_addr_0[39:6] == ldq_18_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_18_0 =
    block_addr_matches_18_0 & lcam_addr_0[5:3] == ldq_18_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_36 = _GEN_524[ldq_18_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_525 =
    fired_release_0 & ldq_18_valid & ldq_18_bits_addr_valid & block_addr_matches_18_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_526 = ldq_18_bits_executed | ldq_18_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_527 = _GEN_526 | l_forwarders_18_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_528 = ldq_18_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_529 =
    do_st_search_0 & ldq_18_valid & ldq_18_bits_addr_valid & _GEN_527
    & ~ldq_18_bits_addr_is_virtual & _GEN_528[0] & dword_addr_matches_18_0
    & (|_mask_overlap_T_36);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_530 =
    do_ld_search_0 & ldq_18_valid & ldq_18_bits_addr_valid & ~ldq_18_bits_addr_is_virtual
    & dword_addr_matches_18_0 & (|_mask_overlap_T_36);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_18 =
    lcam_ldq_idx_0 < 5'h12 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h12;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_531 = lcam_ldq_idx_0 != 5'h12;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_18;	// lsu.scala:1128:57
  wire              _GEN_532 = ~_GEN_526 | nacking_loads_18 | older_nacked_REG_18;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_533 = _GEN_525 | _GEN_529;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_18;	// lsu.scala:1131:58
  wire              _GEN_534 =
    _GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_287 = 15'h1 << ldq_19_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_291 =
    15'h3 << {12'h0, ldq_19_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_535 =
    {{8'hFF},
     {ldq_19_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_291[7:0]},
     {_l_mask_mask_T_287[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_19_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h13;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_19_0 =
    lcam_addr_0[39:6] == ldq_19_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_19_0 =
    block_addr_matches_19_0 & lcam_addr_0[5:3] == ldq_19_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_38 = _GEN_535[ldq_19_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_536 =
    fired_release_0 & ldq_19_valid & ldq_19_bits_addr_valid & block_addr_matches_19_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_537 = ldq_19_bits_executed | ldq_19_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_538 = _GEN_537 | l_forwarders_19_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_539 = ldq_19_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_540 =
    do_st_search_0 & ldq_19_valid & ldq_19_bits_addr_valid & _GEN_538
    & ~ldq_19_bits_addr_is_virtual & _GEN_539[0] & dword_addr_matches_19_0
    & (|_mask_overlap_T_38);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_541 =
    do_ld_search_0 & ldq_19_valid & ldq_19_bits_addr_valid & ~ldq_19_bits_addr_is_virtual
    & dword_addr_matches_19_0 & (|_mask_overlap_T_38);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_19 =
    lcam_ldq_idx_0 < 5'h13 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h13;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_542 = lcam_ldq_idx_0 != 5'h13;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_19;	// lsu.scala:1128:57
  wire              _GEN_543 = ~_GEN_537 | nacking_loads_19 | older_nacked_REG_19;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_544 = _GEN_536 | _GEN_540;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_19;	// lsu.scala:1131:58
  wire              _GEN_545 =
    _GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_302 = 15'h1 << ldq_20_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_306 =
    15'h3 << {12'h0, ldq_20_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_546 =
    {{8'hFF},
     {ldq_20_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_306[7:0]},
     {_l_mask_mask_T_302[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_20_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h14;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_20_0 =
    lcam_addr_0[39:6] == ldq_20_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_20_0 =
    block_addr_matches_20_0 & lcam_addr_0[5:3] == ldq_20_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_40 = _GEN_546[ldq_20_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_547 =
    fired_release_0 & ldq_20_valid & ldq_20_bits_addr_valid & block_addr_matches_20_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_548 = ldq_20_bits_executed | ldq_20_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_549 = _GEN_548 | l_forwarders_20_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_550 = ldq_20_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_551 =
    do_st_search_0 & ldq_20_valid & ldq_20_bits_addr_valid & _GEN_549
    & ~ldq_20_bits_addr_is_virtual & _GEN_550[0] & dword_addr_matches_20_0
    & (|_mask_overlap_T_40);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_552 =
    do_ld_search_0 & ldq_20_valid & ldq_20_bits_addr_valid & ~ldq_20_bits_addr_is_virtual
    & dword_addr_matches_20_0 & (|_mask_overlap_T_40);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_20 =
    lcam_ldq_idx_0 < 5'h14 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h14;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_553 = lcam_ldq_idx_0 != 5'h14;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_20;	// lsu.scala:1128:57
  wire              _GEN_554 = ~_GEN_548 | nacking_loads_20 | older_nacked_REG_20;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_555 = _GEN_547 | _GEN_551;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_20;	// lsu.scala:1131:58
  wire              _GEN_556 =
    _GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_317 = 15'h1 << ldq_21_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_321 =
    15'h3 << {12'h0, ldq_21_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_557 =
    {{8'hFF},
     {ldq_21_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_321[7:0]},
     {_l_mask_mask_T_317[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_21_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h15;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_21_0 =
    lcam_addr_0[39:6] == ldq_21_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_21_0 =
    block_addr_matches_21_0 & lcam_addr_0[5:3] == ldq_21_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_42 = _GEN_557[ldq_21_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_558 =
    fired_release_0 & ldq_21_valid & ldq_21_bits_addr_valid & block_addr_matches_21_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_559 = ldq_21_bits_executed | ldq_21_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_560 = _GEN_559 | l_forwarders_21_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_561 = ldq_21_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_562 =
    do_st_search_0 & ldq_21_valid & ldq_21_bits_addr_valid & _GEN_560
    & ~ldq_21_bits_addr_is_virtual & _GEN_561[0] & dword_addr_matches_21_0
    & (|_mask_overlap_T_42);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_563 =
    do_ld_search_0 & ldq_21_valid & ldq_21_bits_addr_valid & ~ldq_21_bits_addr_is_virtual
    & dword_addr_matches_21_0 & (|_mask_overlap_T_42);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_21 =
    lcam_ldq_idx_0 < 5'h15 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h15;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_564 = lcam_ldq_idx_0 != 5'h15;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_21;	// lsu.scala:1128:57
  wire              _GEN_565 = ~_GEN_559 | nacking_loads_21 | older_nacked_REG_21;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_566 = _GEN_558 | _GEN_562;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_21;	// lsu.scala:1131:58
  wire              _GEN_567 =
    _GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_332 = 15'h1 << ldq_22_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_336 =
    15'h3 << {12'h0, ldq_22_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_568 =
    {{8'hFF},
     {ldq_22_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_336[7:0]},
     {_l_mask_mask_T_332[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_22_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h16;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_22_0 =
    lcam_addr_0[39:6] == ldq_22_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_22_0 =
    block_addr_matches_22_0 & lcam_addr_0[5:3] == ldq_22_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_44 = _GEN_568[ldq_22_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_569 =
    fired_release_0 & ldq_22_valid & ldq_22_bits_addr_valid & block_addr_matches_22_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_570 = ldq_22_bits_executed | ldq_22_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_571 = _GEN_570 | l_forwarders_22_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_572 = ldq_22_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_573 =
    do_st_search_0 & ldq_22_valid & ldq_22_bits_addr_valid & _GEN_571
    & ~ldq_22_bits_addr_is_virtual & _GEN_572[0] & dword_addr_matches_22_0
    & (|_mask_overlap_T_44);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_574 =
    do_ld_search_0 & ldq_22_valid & ldq_22_bits_addr_valid & ~ldq_22_bits_addr_is_virtual
    & dword_addr_matches_22_0 & (|_mask_overlap_T_44);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_22 =
    lcam_ldq_idx_0 < 5'h16 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h16;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_575 = lcam_ldq_idx_0 != 5'h16;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_22;	// lsu.scala:1128:57
  wire              _GEN_576 = ~_GEN_570 | nacking_loads_22 | older_nacked_REG_22;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_577 = _GEN_569 | _GEN_573;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_22;	// lsu.scala:1131:58
  wire              _GEN_578 =
    _GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_347 = 15'h1 << ldq_23_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_351 =
    15'h3 << {12'h0, ldq_23_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_579 =
    {{8'hFF},
     {ldq_23_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_351[7:0]},
     {_l_mask_mask_T_347[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_23_0 =
    wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h17;	// lsu.scala:1064:36, :1065:36, :1075:{63,88}, util.scala:205:25
  wire              block_addr_matches_23_0 =
    lcam_addr_0[39:6] == ldq_23_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_23_0 =
    block_addr_matches_23_0 & lcam_addr_0[5:3] == ldq_23_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_46 = _GEN_579[ldq_23_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_580 =
    fired_release_0 & ldq_23_valid & ldq_23_bits_addr_valid & block_addr_matches_23_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_581 = ldq_23_bits_executed | ldq_23_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_582 = _GEN_581 | l_forwarders_23_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [23:0]       _GEN_583 = ldq_23_bits_st_dep_mask >> _GEN_330;	// lsu.scala:210:16, :1100:38
  wire              _GEN_584 =
    do_st_search_0 & ldq_23_valid & ldq_23_bits_addr_valid & _GEN_582
    & ~ldq_23_bits_addr_is_virtual & _GEN_583[0] & dword_addr_matches_23_0
    & (|_mask_overlap_T_46);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_585 =
    do_ld_search_0 & ldq_23_valid & ldq_23_bits_addr_valid & ~ldq_23_bits_addr_is_virtual
    & dword_addr_matches_23_0 & (|_mask_overlap_T_46);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_23 =
    lcam_ldq_idx_0 < 5'h17 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h17;	// lsu.scala:215:29, :1036:26, util.scala:205:25, :363:{52,64,72,78}
  wire              _GEN_586 = lcam_ldq_idx_0 != 5'h17;	// lsu.scala:1036:26, :1125:38, util.scala:205:25
  reg               older_nacked_REG_23;	// lsu.scala:1128:57
  wire              _GEN_587 = ~_GEN_581 | nacking_loads_23 | older_nacked_REG_23;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_588 = _GEN_580 | _GEN_584;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_23;	// lsu.scala:1131:58
  wire              _GEN_589 =
    _GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire              _GEN_590 =
    _GEN_589
      ? (_GEN_578
           ? (_GEN_567
                ? (_GEN_556
                     ? (_GEN_545
                          ? (_GEN_534
                               ? (_GEN_523
                                    ? (_GEN_512
                                         ? (_GEN_501
                                              ? (_GEN_490
                                                   ? (_GEN_479
                                                        ? (_GEN_468
                                                             ? (_GEN_457
                                                                  ? (_GEN_446
                                                                       ? (_GEN_435
                                                                            ? (_GEN_424
                                                                                 ? (_GEN_413
                                                                                      ? (_GEN_402
                                                                                           ? (_GEN_391
                                                                                                ? (_GEN_380
                                                                                                     ? (_GEN_369
                                                                                                          ? (_GEN_358
                                                                                                               ? (_GEN_347
                                                                                                                    ? ~_GEN_335
                                                                                                                      & _GEN_333
                                                                                                                      & ~searcher_is_older
                                                                                                                      & _GEN_336
                                                                                                                      & io_dmem_s1_kill_0_REG
                                                                                                                    : io_dmem_s1_kill_0_REG_1)
                                                                                                               : io_dmem_s1_kill_0_REG_2)
                                                                                                          : io_dmem_s1_kill_0_REG_3)
                                                                                                     : io_dmem_s1_kill_0_REG_4)
                                                                                                : io_dmem_s1_kill_0_REG_5)
                                                                                           : io_dmem_s1_kill_0_REG_6)
                                                                                      : io_dmem_s1_kill_0_REG_7)
                                                                                 : io_dmem_s1_kill_0_REG_8)
                                                                            : io_dmem_s1_kill_0_REG_9)
                                                                       : io_dmem_s1_kill_0_REG_10)
                                                                  : io_dmem_s1_kill_0_REG_11)
                                                             : io_dmem_s1_kill_0_REG_12)
                                                        : io_dmem_s1_kill_0_REG_13)
                                                   : io_dmem_s1_kill_0_REG_14)
                                              : io_dmem_s1_kill_0_REG_15)
                                         : io_dmem_s1_kill_0_REG_16)
                                    : io_dmem_s1_kill_0_REG_17)
                               : io_dmem_s1_kill_0_REG_18)
                          : io_dmem_s1_kill_0_REG_19)
                     : io_dmem_s1_kill_0_REG_20)
                : io_dmem_s1_kill_0_REG_21)
           : io_dmem_s1_kill_0_REG_22)
      : io_dmem_s1_kill_0_REG_23;	// lsu.scala:764:24, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:47, :1129:73, :1131:{48,58}, util.scala:363:72
  wire              can_forward_0 =
    _GEN_589 & _GEN_578 & _GEN_567 & _GEN_556 & _GEN_545 & _GEN_534 & _GEN_523 & _GEN_512
    & _GEN_501 & _GEN_490 & _GEN_479 & _GEN_468 & _GEN_457 & _GEN_446 & _GEN_435
    & _GEN_424 & _GEN_413 & _GEN_402 & _GEN_391 & _GEN_380 & _GEN_369 & _GEN_358
    & _GEN_347 & (_GEN_335 | ~_GEN_333 | searcher_is_older | ~_GEN_336)
    & (_can_forward_T ? ~mem_tlb_uncacheable_0 : ~_GEN_212[lcam_ldq_idx_0]);	// lsu.scala:502:88, :764:24, :926:41, :1016:61, :1036:26, :1045:{8,56}, :1046:7, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:47, :1129:73, :1131:48, :1132:48, util.scala:363:72
  wire              dword_addr_matches_24_0 =
    stq_0_bits_addr_valid & ~stq_0_bits_addr_is_virtual
    & stq_0_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_2 = 15'h1 << stq_0_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_6 =
    15'h3 << {12'h0, stq_0_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_591 =
    {{8'hFF},
     {stq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_6[7:0]},
     {_write_mask_mask_T_2[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_592 = do_ld_search_0 & stq_0_valid & lcam_st_dep_mask_0[0];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_593 = lcam_mask_0 & _GEN_591[stq_0_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_594 =
    _GEN_593 == lcam_mask_0 & ~stq_0_bits_uop_is_fence & dword_addr_matches_24_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_24;	// lsu.scala:1153:56
  wire              _GEN_595 = (|_GEN_593) & dword_addr_matches_24_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_25;	// lsu.scala:1159:56
  wire              _GEN_596 = stq_0_bits_uop_is_fence | stq_0_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_0 = _GEN_592 & (_GEN_594 | _GEN_595 | _GEN_596);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_26;	// lsu.scala:1165:56
  wire              _GEN_597 =
    _GEN_592
      ? (_GEN_594
           ? io_dmem_s1_kill_0_REG_24
           : _GEN_595
               ? io_dmem_s1_kill_0_REG_25
               : _GEN_596 ? io_dmem_s1_kill_0_REG_26 : _GEN_590)
      : _GEN_590;	// lsu.scala:1091:36, :1102:37, :1116:37, :1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_25_0 =
    stq_1_bits_addr_valid & ~stq_1_bits_addr_is_virtual
    & stq_1_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_17 = 15'h1 << stq_1_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_21 =
    15'h3 << {12'h0, stq_1_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_598 =
    {{8'hFF},
     {stq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_21[7:0]},
     {_write_mask_mask_T_17[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_599 = do_ld_search_0 & stq_1_valid & lcam_st_dep_mask_0[1];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_600 = lcam_mask_0 & _GEN_598[stq_1_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_601 =
    _GEN_600 == lcam_mask_0 & ~stq_1_bits_uop_is_fence & dword_addr_matches_25_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_27;	// lsu.scala:1153:56
  wire              _GEN_602 = (|_GEN_600) & dword_addr_matches_25_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_28;	// lsu.scala:1159:56
  wire              _GEN_603 = stq_1_bits_uop_is_fence | stq_1_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_1 = _GEN_599 & (_GEN_601 | _GEN_602 | _GEN_603);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_29;	// lsu.scala:1165:56
  wire              _GEN_604 =
    _GEN_599
      ? (_GEN_601
           ? io_dmem_s1_kill_0_REG_27
           : _GEN_602
               ? io_dmem_s1_kill_0_REG_28
               : _GEN_603 ? io_dmem_s1_kill_0_REG_29 : _GEN_597)
      : _GEN_597;	// lsu.scala:1091:36, :1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_26_0 =
    stq_2_bits_addr_valid & ~stq_2_bits_addr_is_virtual
    & stq_2_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_32 = 15'h1 << stq_2_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_36 =
    15'h3 << {12'h0, stq_2_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_605 =
    {{8'hFF},
     {stq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_36[7:0]},
     {_write_mask_mask_T_32[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_606 = do_ld_search_0 & stq_2_valid & lcam_st_dep_mask_0[2];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_607 = lcam_mask_0 & _GEN_605[stq_2_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_608 =
    _GEN_607 == lcam_mask_0 & ~stq_2_bits_uop_is_fence & dword_addr_matches_26_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_30;	// lsu.scala:1153:56
  wire              _GEN_609 = (|_GEN_607) & dword_addr_matches_26_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_31;	// lsu.scala:1159:56
  wire              _GEN_610 = stq_2_bits_uop_is_fence | stq_2_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_2 = _GEN_606 & (_GEN_608 | _GEN_609 | _GEN_610);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_32;	// lsu.scala:1165:56
  wire              _GEN_611 =
    _GEN_606
      ? (_GEN_608
           ? io_dmem_s1_kill_0_REG_30
           : _GEN_609
               ? io_dmem_s1_kill_0_REG_31
               : _GEN_610 ? io_dmem_s1_kill_0_REG_32 : _GEN_604)
      : _GEN_604;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_27_0 =
    stq_3_bits_addr_valid & ~stq_3_bits_addr_is_virtual
    & stq_3_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_47 = 15'h1 << stq_3_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_51 =
    15'h3 << {12'h0, stq_3_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_612 =
    {{8'hFF},
     {stq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_51[7:0]},
     {_write_mask_mask_T_47[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_613 = do_ld_search_0 & stq_3_valid & lcam_st_dep_mask_0[3];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_614 = lcam_mask_0 & _GEN_612[stq_3_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_615 =
    _GEN_614 == lcam_mask_0 & ~stq_3_bits_uop_is_fence & dword_addr_matches_27_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_33;	// lsu.scala:1153:56
  wire              _GEN_616 = (|_GEN_614) & dword_addr_matches_27_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_34;	// lsu.scala:1159:56
  wire              _GEN_617 = stq_3_bits_uop_is_fence | stq_3_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_3 = _GEN_613 & (_GEN_615 | _GEN_616 | _GEN_617);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_35;	// lsu.scala:1165:56
  wire              _GEN_618 =
    _GEN_613
      ? (_GEN_615
           ? io_dmem_s1_kill_0_REG_33
           : _GEN_616
               ? io_dmem_s1_kill_0_REG_34
               : _GEN_617 ? io_dmem_s1_kill_0_REG_35 : _GEN_611)
      : _GEN_611;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_28_0 =
    stq_4_bits_addr_valid & ~stq_4_bits_addr_is_virtual
    & stq_4_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_62 = 15'h1 << stq_4_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_66 =
    15'h3 << {12'h0, stq_4_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_619 =
    {{8'hFF},
     {stq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_66[7:0]},
     {_write_mask_mask_T_62[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_620 = do_ld_search_0 & stq_4_valid & lcam_st_dep_mask_0[4];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_621 = lcam_mask_0 & _GEN_619[stq_4_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_622 =
    _GEN_621 == lcam_mask_0 & ~stq_4_bits_uop_is_fence & dword_addr_matches_28_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_36;	// lsu.scala:1153:56
  wire              _GEN_623 = (|_GEN_621) & dword_addr_matches_28_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_37;	// lsu.scala:1159:56
  wire              _GEN_624 = stq_4_bits_uop_is_fence | stq_4_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_4 = _GEN_620 & (_GEN_622 | _GEN_623 | _GEN_624);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_38;	// lsu.scala:1165:56
  wire              _GEN_625 =
    _GEN_620
      ? (_GEN_622
           ? io_dmem_s1_kill_0_REG_36
           : _GEN_623
               ? io_dmem_s1_kill_0_REG_37
               : _GEN_624 ? io_dmem_s1_kill_0_REG_38 : _GEN_618)
      : _GEN_618;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_29_0 =
    stq_5_bits_addr_valid & ~stq_5_bits_addr_is_virtual
    & stq_5_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_77 = 15'h1 << stq_5_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_81 =
    15'h3 << {12'h0, stq_5_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_626 =
    {{8'hFF},
     {stq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_81[7:0]},
     {_write_mask_mask_T_77[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_627 = do_ld_search_0 & stq_5_valid & lcam_st_dep_mask_0[5];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_628 = lcam_mask_0 & _GEN_626[stq_5_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_629 =
    _GEN_628 == lcam_mask_0 & ~stq_5_bits_uop_is_fence & dword_addr_matches_29_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_39;	// lsu.scala:1153:56
  wire              _GEN_630 = (|_GEN_628) & dword_addr_matches_29_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_40;	// lsu.scala:1159:56
  wire              _GEN_631 = stq_5_bits_uop_is_fence | stq_5_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_5 = _GEN_627 & (_GEN_629 | _GEN_630 | _GEN_631);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_41;	// lsu.scala:1165:56
  wire              _GEN_632 =
    _GEN_627
      ? (_GEN_629
           ? io_dmem_s1_kill_0_REG_39
           : _GEN_630
               ? io_dmem_s1_kill_0_REG_40
               : _GEN_631 ? io_dmem_s1_kill_0_REG_41 : _GEN_625)
      : _GEN_625;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_30_0 =
    stq_6_bits_addr_valid & ~stq_6_bits_addr_is_virtual
    & stq_6_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_92 = 15'h1 << stq_6_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_96 =
    15'h3 << {12'h0, stq_6_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_633 =
    {{8'hFF},
     {stq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_96[7:0]},
     {_write_mask_mask_T_92[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_634 = do_ld_search_0 & stq_6_valid & lcam_st_dep_mask_0[6];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_635 = lcam_mask_0 & _GEN_633[stq_6_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_636 =
    _GEN_635 == lcam_mask_0 & ~stq_6_bits_uop_is_fence & dword_addr_matches_30_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_42;	// lsu.scala:1153:56
  wire              _GEN_637 = (|_GEN_635) & dword_addr_matches_30_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_43;	// lsu.scala:1159:56
  wire              _GEN_638 = stq_6_bits_uop_is_fence | stq_6_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_6 = _GEN_634 & (_GEN_636 | _GEN_637 | _GEN_638);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_44;	// lsu.scala:1165:56
  wire              _GEN_639 =
    _GEN_634
      ? (_GEN_636
           ? io_dmem_s1_kill_0_REG_42
           : _GEN_637
               ? io_dmem_s1_kill_0_REG_43
               : _GEN_638 ? io_dmem_s1_kill_0_REG_44 : _GEN_632)
      : _GEN_632;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_31_0 =
    stq_7_bits_addr_valid & ~stq_7_bits_addr_is_virtual
    & stq_7_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_107 = 15'h1 << stq_7_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_111 =
    15'h3 << {12'h0, stq_7_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_640 =
    {{8'hFF},
     {stq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_111[7:0]},
     {_write_mask_mask_T_107[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_641 = do_ld_search_0 & stq_7_valid & lcam_st_dep_mask_0[7];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_642 = lcam_mask_0 & _GEN_640[stq_7_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_643 =
    _GEN_642 == lcam_mask_0 & ~stq_7_bits_uop_is_fence & dword_addr_matches_31_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_45;	// lsu.scala:1153:56
  wire              _GEN_644 = (|_GEN_642) & dword_addr_matches_31_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_46;	// lsu.scala:1159:56
  wire              _GEN_645 = stq_7_bits_uop_is_fence | stq_7_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_7 = _GEN_641 & (_GEN_643 | _GEN_644 | _GEN_645);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_47;	// lsu.scala:1165:56
  wire              _GEN_646 =
    _GEN_641
      ? (_GEN_643
           ? io_dmem_s1_kill_0_REG_45
           : _GEN_644
               ? io_dmem_s1_kill_0_REG_46
               : _GEN_645 ? io_dmem_s1_kill_0_REG_47 : _GEN_639)
      : _GEN_639;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_32_0 =
    stq_8_bits_addr_valid & ~stq_8_bits_addr_is_virtual
    & stq_8_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_122 = 15'h1 << stq_8_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_126 =
    15'h3 << {12'h0, stq_8_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_647 =
    {{8'hFF},
     {stq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_126[7:0]},
     {_write_mask_mask_T_122[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_648 = do_ld_search_0 & stq_8_valid & lcam_st_dep_mask_0[8];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_649 = lcam_mask_0 & _GEN_647[stq_8_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_650 =
    _GEN_649 == lcam_mask_0 & ~stq_8_bits_uop_is_fence & dword_addr_matches_32_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_48;	// lsu.scala:1153:56
  wire              _GEN_651 = (|_GEN_649) & dword_addr_matches_32_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_49;	// lsu.scala:1159:56
  wire              _GEN_652 = stq_8_bits_uop_is_fence | stq_8_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_8 = _GEN_648 & (_GEN_650 | _GEN_651 | _GEN_652);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_50;	// lsu.scala:1165:56
  wire              _GEN_653 =
    _GEN_648
      ? (_GEN_650
           ? io_dmem_s1_kill_0_REG_48
           : _GEN_651
               ? io_dmem_s1_kill_0_REG_49
               : _GEN_652 ? io_dmem_s1_kill_0_REG_50 : _GEN_646)
      : _GEN_646;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_33_0 =
    stq_9_bits_addr_valid & ~stq_9_bits_addr_is_virtual
    & stq_9_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_137 = 15'h1 << stq_9_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_141 =
    15'h3 << {12'h0, stq_9_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_654 =
    {{8'hFF},
     {stq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_141[7:0]},
     {_write_mask_mask_T_137[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_655 = do_ld_search_0 & stq_9_valid & lcam_st_dep_mask_0[9];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_656 = lcam_mask_0 & _GEN_654[stq_9_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_657 =
    _GEN_656 == lcam_mask_0 & ~stq_9_bits_uop_is_fence & dword_addr_matches_33_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_51;	// lsu.scala:1153:56
  wire              _GEN_658 = (|_GEN_656) & dword_addr_matches_33_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_52;	// lsu.scala:1159:56
  wire              _GEN_659 = stq_9_bits_uop_is_fence | stq_9_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_9 = _GEN_655 & (_GEN_657 | _GEN_658 | _GEN_659);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_53;	// lsu.scala:1165:56
  wire              _GEN_660 =
    _GEN_655
      ? (_GEN_657
           ? io_dmem_s1_kill_0_REG_51
           : _GEN_658
               ? io_dmem_s1_kill_0_REG_52
               : _GEN_659 ? io_dmem_s1_kill_0_REG_53 : _GEN_653)
      : _GEN_653;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_34_0 =
    stq_10_bits_addr_valid & ~stq_10_bits_addr_is_virtual
    & stq_10_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_152 = 15'h1 << stq_10_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_156 =
    15'h3 << {12'h0, stq_10_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_661 =
    {{8'hFF},
     {stq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_156[7:0]},
     {_write_mask_mask_T_152[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_662 = do_ld_search_0 & stq_10_valid & lcam_st_dep_mask_0[10];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_663 = lcam_mask_0 & _GEN_661[stq_10_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_664 =
    _GEN_663 == lcam_mask_0 & ~stq_10_bits_uop_is_fence & dword_addr_matches_34_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_54;	// lsu.scala:1153:56
  wire              _GEN_665 = (|_GEN_663) & dword_addr_matches_34_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_55;	// lsu.scala:1159:56
  wire              _GEN_666 = stq_10_bits_uop_is_fence | stq_10_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_10 = _GEN_662 & (_GEN_664 | _GEN_665 | _GEN_666);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_56;	// lsu.scala:1165:56
  wire              _GEN_667 =
    _GEN_662
      ? (_GEN_664
           ? io_dmem_s1_kill_0_REG_54
           : _GEN_665
               ? io_dmem_s1_kill_0_REG_55
               : _GEN_666 ? io_dmem_s1_kill_0_REG_56 : _GEN_660)
      : _GEN_660;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_35_0 =
    stq_11_bits_addr_valid & ~stq_11_bits_addr_is_virtual
    & stq_11_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_167 = 15'h1 << stq_11_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_171 =
    15'h3 << {12'h0, stq_11_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_668 =
    {{8'hFF},
     {stq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_171[7:0]},
     {_write_mask_mask_T_167[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_669 = do_ld_search_0 & stq_11_valid & lcam_st_dep_mask_0[11];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_670 = lcam_mask_0 & _GEN_668[stq_11_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_671 =
    _GEN_670 == lcam_mask_0 & ~stq_11_bits_uop_is_fence & dword_addr_matches_35_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_57;	// lsu.scala:1153:56
  wire              _GEN_672 = (|_GEN_670) & dword_addr_matches_35_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_58;	// lsu.scala:1159:56
  wire              _GEN_673 = stq_11_bits_uop_is_fence | stq_11_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_11 = _GEN_669 & (_GEN_671 | _GEN_672 | _GEN_673);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_59;	// lsu.scala:1165:56
  wire              _GEN_674 =
    _GEN_669
      ? (_GEN_671
           ? io_dmem_s1_kill_0_REG_57
           : _GEN_672
               ? io_dmem_s1_kill_0_REG_58
               : _GEN_673 ? io_dmem_s1_kill_0_REG_59 : _GEN_667)
      : _GEN_667;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_36_0 =
    stq_12_bits_addr_valid & ~stq_12_bits_addr_is_virtual
    & stq_12_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_182 = 15'h1 << stq_12_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_186 =
    15'h3 << {12'h0, stq_12_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_675 =
    {{8'hFF},
     {stq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_186[7:0]},
     {_write_mask_mask_T_182[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_676 = do_ld_search_0 & stq_12_valid & lcam_st_dep_mask_0[12];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_677 = lcam_mask_0 & _GEN_675[stq_12_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_678 =
    _GEN_677 == lcam_mask_0 & ~stq_12_bits_uop_is_fence & dword_addr_matches_36_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_60;	// lsu.scala:1153:56
  wire              _GEN_679 = (|_GEN_677) & dword_addr_matches_36_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_61;	// lsu.scala:1159:56
  wire              _GEN_680 = stq_12_bits_uop_is_fence | stq_12_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_12 = _GEN_676 & (_GEN_678 | _GEN_679 | _GEN_680);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_62;	// lsu.scala:1165:56
  wire              _GEN_681 =
    _GEN_676
      ? (_GEN_678
           ? io_dmem_s1_kill_0_REG_60
           : _GEN_679
               ? io_dmem_s1_kill_0_REG_61
               : _GEN_680 ? io_dmem_s1_kill_0_REG_62 : _GEN_674)
      : _GEN_674;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_37_0 =
    stq_13_bits_addr_valid & ~stq_13_bits_addr_is_virtual
    & stq_13_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_197 = 15'h1 << stq_13_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_201 =
    15'h3 << {12'h0, stq_13_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_682 =
    {{8'hFF},
     {stq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_201[7:0]},
     {_write_mask_mask_T_197[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_683 = do_ld_search_0 & stq_13_valid & lcam_st_dep_mask_0[13];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_684 = lcam_mask_0 & _GEN_682[stq_13_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_685 =
    _GEN_684 == lcam_mask_0 & ~stq_13_bits_uop_is_fence & dword_addr_matches_37_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_63;	// lsu.scala:1153:56
  wire              _GEN_686 = (|_GEN_684) & dword_addr_matches_37_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_64;	// lsu.scala:1159:56
  wire              _GEN_687 = stq_13_bits_uop_is_fence | stq_13_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_13 = _GEN_683 & (_GEN_685 | _GEN_686 | _GEN_687);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_65;	// lsu.scala:1165:56
  wire              _GEN_688 =
    _GEN_683
      ? (_GEN_685
           ? io_dmem_s1_kill_0_REG_63
           : _GEN_686
               ? io_dmem_s1_kill_0_REG_64
               : _GEN_687 ? io_dmem_s1_kill_0_REG_65 : _GEN_681)
      : _GEN_681;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_38_0 =
    stq_14_bits_addr_valid & ~stq_14_bits_addr_is_virtual
    & stq_14_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_212 = 15'h1 << stq_14_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_216 =
    15'h3 << {12'h0, stq_14_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_689 =
    {{8'hFF},
     {stq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_216[7:0]},
     {_write_mask_mask_T_212[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_690 = do_ld_search_0 & stq_14_valid & lcam_st_dep_mask_0[14];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_691 = lcam_mask_0 & _GEN_689[stq_14_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_692 =
    _GEN_691 == lcam_mask_0 & ~stq_14_bits_uop_is_fence & dword_addr_matches_38_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_66;	// lsu.scala:1153:56
  wire              _GEN_693 = (|_GEN_691) & dword_addr_matches_38_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_67;	// lsu.scala:1159:56
  wire              _GEN_694 = stq_14_bits_uop_is_fence | stq_14_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_14 = _GEN_690 & (_GEN_692 | _GEN_693 | _GEN_694);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_68;	// lsu.scala:1165:56
  wire              _GEN_695 =
    _GEN_690
      ? (_GEN_692
           ? io_dmem_s1_kill_0_REG_66
           : _GEN_693
               ? io_dmem_s1_kill_0_REG_67
               : _GEN_694 ? io_dmem_s1_kill_0_REG_68 : _GEN_688)
      : _GEN_688;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_39_0 =
    stq_15_bits_addr_valid & ~stq_15_bits_addr_is_virtual
    & stq_15_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_227 = 15'h1 << stq_15_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_231 =
    15'h3 << {12'h0, stq_15_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_696 =
    {{8'hFF},
     {stq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_231[7:0]},
     {_write_mask_mask_T_227[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_697 = do_ld_search_0 & stq_15_valid & lcam_st_dep_mask_0[15];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_698 = lcam_mask_0 & _GEN_696[stq_15_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_699 =
    _GEN_698 == lcam_mask_0 & ~stq_15_bits_uop_is_fence & dword_addr_matches_39_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_69;	// lsu.scala:1153:56
  wire              _GEN_700 = (|_GEN_698) & dword_addr_matches_39_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_70;	// lsu.scala:1159:56
  wire              _GEN_701 = stq_15_bits_uop_is_fence | stq_15_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_15 = _GEN_697 & (_GEN_699 | _GEN_700 | _GEN_701);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_71;	// lsu.scala:1165:56
  wire              _GEN_702 =
    _GEN_697
      ? (_GEN_699
           ? io_dmem_s1_kill_0_REG_69
           : _GEN_700
               ? io_dmem_s1_kill_0_REG_70
               : _GEN_701 ? io_dmem_s1_kill_0_REG_71 : _GEN_695)
      : _GEN_695;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_40_0 =
    stq_16_bits_addr_valid & ~stq_16_bits_addr_is_virtual
    & stq_16_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_242 = 15'h1 << stq_16_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_246 =
    15'h3 << {12'h0, stq_16_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_703 =
    {{8'hFF},
     {stq_16_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_246[7:0]},
     {_write_mask_mask_T_242[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_704 = do_ld_search_0 & stq_16_valid & lcam_st_dep_mask_0[16];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_705 = lcam_mask_0 & _GEN_703[stq_16_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_706 =
    _GEN_705 == lcam_mask_0 & ~stq_16_bits_uop_is_fence & dword_addr_matches_40_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_72;	// lsu.scala:1153:56
  wire              _GEN_707 = (|_GEN_705) & dword_addr_matches_40_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_73;	// lsu.scala:1159:56
  wire              _GEN_708 = stq_16_bits_uop_is_fence | stq_16_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_16 = _GEN_704 & (_GEN_706 | _GEN_707 | _GEN_708);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_74;	// lsu.scala:1165:56
  wire              _GEN_709 =
    _GEN_704
      ? (_GEN_706
           ? io_dmem_s1_kill_0_REG_72
           : _GEN_707
               ? io_dmem_s1_kill_0_REG_73
               : _GEN_708 ? io_dmem_s1_kill_0_REG_74 : _GEN_702)
      : _GEN_702;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_41_0 =
    stq_17_bits_addr_valid & ~stq_17_bits_addr_is_virtual
    & stq_17_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_257 = 15'h1 << stq_17_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_261 =
    15'h3 << {12'h0, stq_17_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_710 =
    {{8'hFF},
     {stq_17_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_261[7:0]},
     {_write_mask_mask_T_257[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_711 = do_ld_search_0 & stq_17_valid & lcam_st_dep_mask_0[17];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_712 = lcam_mask_0 & _GEN_710[stq_17_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_713 =
    _GEN_712 == lcam_mask_0 & ~stq_17_bits_uop_is_fence & dword_addr_matches_41_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_75;	// lsu.scala:1153:56
  wire              _GEN_714 = (|_GEN_712) & dword_addr_matches_41_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_76;	// lsu.scala:1159:56
  wire              _GEN_715 = stq_17_bits_uop_is_fence | stq_17_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_17 = _GEN_711 & (_GEN_713 | _GEN_714 | _GEN_715);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_77;	// lsu.scala:1165:56
  wire              _GEN_716 =
    _GEN_711
      ? (_GEN_713
           ? io_dmem_s1_kill_0_REG_75
           : _GEN_714
               ? io_dmem_s1_kill_0_REG_76
               : _GEN_715 ? io_dmem_s1_kill_0_REG_77 : _GEN_709)
      : _GEN_709;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_42_0 =
    stq_18_bits_addr_valid & ~stq_18_bits_addr_is_virtual
    & stq_18_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_272 = 15'h1 << stq_18_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_276 =
    15'h3 << {12'h0, stq_18_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_717 =
    {{8'hFF},
     {stq_18_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_276[7:0]},
     {_write_mask_mask_T_272[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_718 = do_ld_search_0 & stq_18_valid & lcam_st_dep_mask_0[18];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_719 = lcam_mask_0 & _GEN_717[stq_18_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_720 =
    _GEN_719 == lcam_mask_0 & ~stq_18_bits_uop_is_fence & dword_addr_matches_42_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_78;	// lsu.scala:1153:56
  wire              _GEN_721 = (|_GEN_719) & dword_addr_matches_42_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_79;	// lsu.scala:1159:56
  wire              _GEN_722 = stq_18_bits_uop_is_fence | stq_18_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_18 = _GEN_718 & (_GEN_720 | _GEN_721 | _GEN_722);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_80;	// lsu.scala:1165:56
  wire              _GEN_723 =
    _GEN_718
      ? (_GEN_720
           ? io_dmem_s1_kill_0_REG_78
           : _GEN_721
               ? io_dmem_s1_kill_0_REG_79
               : _GEN_722 ? io_dmem_s1_kill_0_REG_80 : _GEN_716)
      : _GEN_716;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_43_0 =
    stq_19_bits_addr_valid & ~stq_19_bits_addr_is_virtual
    & stq_19_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_287 = 15'h1 << stq_19_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_291 =
    15'h3 << {12'h0, stq_19_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_724 =
    {{8'hFF},
     {stq_19_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_291[7:0]},
     {_write_mask_mask_T_287[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_725 = do_ld_search_0 & stq_19_valid & lcam_st_dep_mask_0[19];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_726 = lcam_mask_0 & _GEN_724[stq_19_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_727 =
    _GEN_726 == lcam_mask_0 & ~stq_19_bits_uop_is_fence & dword_addr_matches_43_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_81;	// lsu.scala:1153:56
  wire              _GEN_728 = (|_GEN_726) & dword_addr_matches_43_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_82;	// lsu.scala:1159:56
  wire              _GEN_729 = stq_19_bits_uop_is_fence | stq_19_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_19 = _GEN_725 & (_GEN_727 | _GEN_728 | _GEN_729);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_83;	// lsu.scala:1165:56
  wire              _GEN_730 =
    _GEN_725
      ? (_GEN_727
           ? io_dmem_s1_kill_0_REG_81
           : _GEN_728
               ? io_dmem_s1_kill_0_REG_82
               : _GEN_729 ? io_dmem_s1_kill_0_REG_83 : _GEN_723)
      : _GEN_723;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_44_0 =
    stq_20_bits_addr_valid & ~stq_20_bits_addr_is_virtual
    & stq_20_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_302 = 15'h1 << stq_20_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_306 =
    15'h3 << {12'h0, stq_20_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_731 =
    {{8'hFF},
     {stq_20_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_306[7:0]},
     {_write_mask_mask_T_302[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_732 = do_ld_search_0 & stq_20_valid & lcam_st_dep_mask_0[20];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_733 = lcam_mask_0 & _GEN_731[stq_20_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_734 =
    _GEN_733 == lcam_mask_0 & ~stq_20_bits_uop_is_fence & dword_addr_matches_44_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_84;	// lsu.scala:1153:56
  wire              _GEN_735 = (|_GEN_733) & dword_addr_matches_44_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_85;	// lsu.scala:1159:56
  wire              _GEN_736 = stq_20_bits_uop_is_fence | stq_20_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_20 = _GEN_732 & (_GEN_734 | _GEN_735 | _GEN_736);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_86;	// lsu.scala:1165:56
  wire              _GEN_737 =
    _GEN_732
      ? (_GEN_734
           ? io_dmem_s1_kill_0_REG_84
           : _GEN_735
               ? io_dmem_s1_kill_0_REG_85
               : _GEN_736 ? io_dmem_s1_kill_0_REG_86 : _GEN_730)
      : _GEN_730;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_45_0 =
    stq_21_bits_addr_valid & ~stq_21_bits_addr_is_virtual
    & stq_21_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_317 = 15'h1 << stq_21_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_321 =
    15'h3 << {12'h0, stq_21_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_738 =
    {{8'hFF},
     {stq_21_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_321[7:0]},
     {_write_mask_mask_T_317[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_739 = do_ld_search_0 & stq_21_valid & lcam_st_dep_mask_0[21];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_740 = lcam_mask_0 & _GEN_738[stq_21_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_741 =
    _GEN_740 == lcam_mask_0 & ~stq_21_bits_uop_is_fence & dword_addr_matches_45_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_87;	// lsu.scala:1153:56
  wire              _GEN_742 = (|_GEN_740) & dword_addr_matches_45_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_88;	// lsu.scala:1159:56
  wire              _GEN_743 = stq_21_bits_uop_is_fence | stq_21_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_21 = _GEN_739 & (_GEN_741 | _GEN_742 | _GEN_743);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_89;	// lsu.scala:1165:56
  wire              _GEN_744 =
    _GEN_739
      ? (_GEN_741
           ? io_dmem_s1_kill_0_REG_87
           : _GEN_742
               ? io_dmem_s1_kill_0_REG_88
               : _GEN_743 ? io_dmem_s1_kill_0_REG_89 : _GEN_737)
      : _GEN_737;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_46_0 =
    stq_22_bits_addr_valid & ~stq_22_bits_addr_is_virtual
    & stq_22_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_332 = 15'h1 << stq_22_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_336 =
    15'h3 << {12'h0, stq_22_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_745 =
    {{8'hFF},
     {stq_22_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_336[7:0]},
     {_write_mask_mask_T_332[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_746 = do_ld_search_0 & stq_22_valid & lcam_st_dep_mask_0[22];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_747 = lcam_mask_0 & _GEN_745[stq_22_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_748 =
    _GEN_747 == lcam_mask_0 & ~stq_22_bits_uop_is_fence & dword_addr_matches_46_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_90;	// lsu.scala:1153:56
  wire              _GEN_749 = (|_GEN_747) & dword_addr_matches_46_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_91;	// lsu.scala:1159:56
  wire              _GEN_750 = stq_22_bits_uop_is_fence | stq_22_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_22 = _GEN_746 & (_GEN_748 | _GEN_749 | _GEN_750);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_92;	// lsu.scala:1165:56
  wire              _GEN_751 =
    _GEN_746
      ? (_GEN_748
           ? io_dmem_s1_kill_0_REG_90
           : _GEN_749
               ? io_dmem_s1_kill_0_REG_91
               : _GEN_750 ? io_dmem_s1_kill_0_REG_92 : _GEN_744)
      : _GEN_744;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_47_0 =
    stq_23_bits_addr_valid & ~stq_23_bits_addr_is_virtual
    & stq_23_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_347 = 15'h1 << stq_23_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_351 =
    15'h3 << {12'h0, stq_23_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_752 =
    {{8'hFF},
     {stq_23_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_351[7:0]},
     {_write_mask_mask_T_347[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_753 = do_ld_search_0 & stq_23_valid & lcam_st_dep_mask_0[23];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_754 = lcam_mask_0 & _GEN_752[stq_23_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_755 =
    _GEN_754 == lcam_mask_0 & ~stq_23_bits_uop_is_fence & dword_addr_matches_47_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_93;	// lsu.scala:1153:56
  wire              _GEN_756 = (|_GEN_754) & dword_addr_matches_47_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_94;	// lsu.scala:1159:56
  wire              _GEN_757 = stq_23_bits_uop_is_fence | stq_23_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_23 = _GEN_753 & (_GEN_755 | _GEN_756 | _GEN_757);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_95;	// lsu.scala:1165:56
  reg               REG_1;	// lsu.scala:1189:64
  reg               REG_2;	// lsu.scala:1199:18
  reg  [3:0]        store_blocked_counter;	// lsu.scala:1204:36
  assign block_load_wakeup = (&store_blocked_counter) | REG_2;	// lsu.scala:1199:{18,80}, :1204:36, :1210:{33,43}, :1211:25
  reg               r_xcpt_valid;	// lsu.scala:1235:29
  reg  [15:0]       r_xcpt_uop_br_mask;	// lsu.scala:1236:25
  reg  [6:0]        r_xcpt_uop_rob_idx;	// lsu.scala:1236:25
  reg  [4:0]        r_xcpt_cause;	// lsu.scala:1236:25
  reg  [39:0]       r_xcpt_badvaddr;	// lsu.scala:1236:25
  wire              _io_core_spec_ld_wakeup_0_valid_output =
    fired_load_incoming_REG & ~mem_incoming_uop_0_fp_val & (|mem_incoming_uop_0_pdst);	// lsu.scala:894:51, :908:37, :1260:{40,69}, :1261:65
  wire              _GEN_758 = io_dmem_nack_0_valid & io_dmem_nack_0_bits_is_hella;	// lsu.scala:1287:7
  wire              _GEN_759 = hella_state == 3'h4;	// lsu.scala:242:38, :1288:28, util.scala:351:72
  wire              _GEN_760 = hella_state == 3'h6;	// lsu.scala:242:38, :1288:54, util.scala:351:72
  wire              _GEN_761 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h0;	// lsu.scala:1293:62
  wire              _GEN_762 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1;	// lsu.scala:305:44, :1293:62
  wire              _GEN_763 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h2;	// lsu.scala:305:44, :1293:62
  wire              _GEN_764 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h3;	// lsu.scala:305:44, :1293:62
  wire              _GEN_765 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h4;	// lsu.scala:305:44, :1293:62
  wire              _GEN_766 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h5;	// lsu.scala:305:44, :1293:62
  wire              _GEN_767 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h6;	// lsu.scala:305:44, :1293:62
  wire              _GEN_768 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h7;	// lsu.scala:305:44, :1293:62
  wire              _GEN_769 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h8;	// lsu.scala:305:44, :1293:62
  wire              _GEN_770 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h9;	// lsu.scala:305:44, :1293:62
  wire              _GEN_771 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hA;	// lsu.scala:305:44, :1293:62
  wire              _GEN_772 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hB;	// lsu.scala:305:44, :1293:62
  wire              _GEN_773 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hC;	// lsu.scala:305:44, :1293:62
  wire              _GEN_774 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hD;	// lsu.scala:305:44, :1293:62
  wire              _GEN_775 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hE;	// lsu.scala:305:44, :1293:62
  wire              _GEN_776 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hF;	// lsu.scala:305:44, :1293:62
  wire              _GEN_777 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h10;	// lsu.scala:305:44, :1293:62
  wire              _GEN_778 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h11;	// lsu.scala:305:44, :1293:62
  wire              _GEN_779 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h12;	// lsu.scala:305:44, :1293:62
  wire              _GEN_780 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h13;	// lsu.scala:305:44, :1293:62
  wire              _GEN_781 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h14;	// lsu.scala:305:44, :1293:62
  wire              _GEN_782 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h15;	// lsu.scala:305:44, :1293:62
  wire              _GEN_783 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h16;	// lsu.scala:305:44, :1293:62
  wire              _GEN_784 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h17;	// lsu.scala:1293:62, util.scala:205:25
  assign nacking_loads_0 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_761;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_1 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_762;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_2 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_763;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_3 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_764;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_4 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_765;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_5 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_766;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_6 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_767;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_7 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_768;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_8 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_769;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_9 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_770;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_10 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_771;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_11 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_772;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_12 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_773;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_13 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_774;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_14 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_775;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_15 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_776;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_16 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_777;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_17 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_778;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_18 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_779;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_19 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_780;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_20 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_781;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_21 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_782;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_22 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_783;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_23 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_784;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  wire              _GEN_785 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq;	// lsu.scala:1308:7
  wire              send_iresp = _GEN_185[io_dmem_resp_0_bits_uop_ldq_idx] == 2'h0;	// lsu.scala:465:79, :1311:58
  wire              send_fresp = _GEN_185[io_dmem_resp_0_bits_uop_ldq_idx] == 2'h1;	// lsu.scala:465:79, :1311:58, :1312:58
  wire              _GEN_786 =
    io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_is_amo;	// lsu.scala:1328:7, :1331:48
  wire              dmem_resp_fired_0 =
    io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq | _GEN_786);	// lsu.scala:1306:5, :1308:7, :1322:28, :1328:7, :1331:48
  wire              _GEN_787 = dmem_resp_fired_0 & wb_forward_valid_0;	// lsu.scala:1064:36, :1306:5, :1308:7, :1343:30
  wire              _GEN_788 = ~dmem_resp_fired_0 & wb_forward_valid_0;	// lsu.scala:1064:36, :1306:5, :1308:7, :1347:{18,38}
  wire [15:0]       _GEN_789 = _GEN_110[wb_forward_ldq_idx_0];	// lsu.scala:264:49, :1065:36, util.scala:118:51
  wire [6:0]        _GEN_790 = _GEN_148[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire [6:0]        _GEN_791 = _GEN_153[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire [1:0]        _GEN_792 = _GEN_112[wb_forward_ldq_idx_0];	// lsu.scala:264:49, :1065:36, util.scala:118:51
  wire              _GEN_793 = _GEN_168[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire              _GEN_794 = _GEN_171[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire              _GEN_795 = _GEN_174[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire [1:0]        _GEN_796 = _GEN_185[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire              live = (io_core_brupdate_b1_mispredict_mask & _GEN_789) == 16'h0;	// util.scala:118:{51,59}
  wire              _GEN_797 = _GEN_91[wb_forward_stq_idx_0];	// AMOALU.scala:10:17, lsu.scala:224:42, :1067:36
  wire [63:0]       _GEN_798 = _GEN_92[wb_forward_stq_idx_0];	// AMOALU.scala:10:17, lsu.scala:224:42, :1067:36
  wire [3:0][63:0]  _GEN_799 =
    {{_GEN_798},
     {{2{_GEN_798[31:0]}}},
     {{2{{2{_GEN_798[15:0]}}}}},
     {{2{{2{{2{_GEN_798[7:0]}}}}}}}};	// AMOALU.scala:10:17, :26:{13,19,66}, Cat.scala:30:58
  wire [63:0]       _GEN_800 = _GEN_799[_GEN_55[wb_forward_stq_idx_0]];	// AMOALU.scala:10:17, :26:{13,19}, lsu.scala:224:42, :1067:36
  wire              _GEN_801 = _GEN_787 | ~_GEN_788;	// lsu.scala:1306:5, :1343:30, :1344:5, :1347:38, :1348:5
  wire              _io_core_exe_0_iresp_valid_output =
    _GEN_801
      ? io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq ? send_iresp : _GEN_786)
      : _GEN_796 == 2'h0 & _GEN_797 & live;	// AMOALU.scala:10:17, lsu.scala:1275:32, :1306:5, :1308:7, :1311:58, :1316:40, :1328:7, :1331:48, :1344:5, :1348:5, :1362:{60,86}, util.scala:118:{51,59}
  wire              _io_core_exe_0_fresp_valid_output =
    _GEN_801 ? _GEN_785 & send_fresp : _GEN_796 == 2'h1 & _GEN_797 & live;	// AMOALU.scala:10:17, lsu.scala:1276:32, :1306:5, :1308:7, :1312:58, :1318:40, :1344:5, :1348:5, :1363:{60,86}, util.scala:118:{51,59}
  wire [31:0]       io_core_exe_0_iresp_bits_data_lo =
    wb_forward_ld_addr_0[2] ? _GEN_800[63:32] : _GEN_800[31:0];	// AMOALU.scala:26:13, :39:{24,29,37,55}, lsu.scala:1066:36
  wire              _ldq_bits_debug_wb_data_T_1 = _GEN_792 == 2'h2;	// AMOALU.scala:42:26, util.scala:118:51, :351:72
  wire [15:0]       io_core_exe_0_iresp_bits_data_lo_1 =
    wb_forward_ld_addr_0[1]
      ? io_core_exe_0_iresp_bits_data_lo[31:16]
      : io_core_exe_0_iresp_bits_data_lo[15:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  wire              _ldq_bits_debug_wb_data_T_9 = _GEN_792 == 2'h1;	// AMOALU.scala:42:26, lsu.scala:1312:58, util.scala:118:51
  wire [7:0]        io_core_exe_0_iresp_bits_data_lo_2 =
    wb_forward_ld_addr_0[0]
      ? io_core_exe_0_iresp_bits_data_lo_1[15:8]
      : io_core_exe_0_iresp_bits_data_lo_1[7:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  wire              _ldq_bits_debug_wb_data_T_17 = _GEN_792 == 2'h0;	// AMOALU.scala:42:26, util.scala:118:51
  wire [31:0]       io_core_exe_0_fresp_bits_data_lo =
    wb_forward_ld_addr_0[2] ? _GEN_800[63:32] : _GEN_800[31:0];	// AMOALU.scala:26:13, :39:{24,29,37,55}, lsu.scala:1066:36
  wire [15:0]       io_core_exe_0_fresp_bits_data_lo_1 =
    wb_forward_ld_addr_0[1]
      ? io_core_exe_0_fresp_bits_data_lo[31:16]
      : io_core_exe_0_fresp_bits_data_lo[15:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  wire [7:0]        io_core_exe_0_fresp_bits_data_lo_2 =
    wb_forward_ld_addr_0[0]
      ? io_core_exe_0_fresp_bits_data_lo_1[15:8]
      : io_core_exe_0_fresp_bits_data_lo_1[7:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  reg               io_core_ld_miss_REG;	// lsu.scala:1380:37
  reg               spec_ld_succeed_REG;	// lsu.scala:1382:13
  reg  [4:0]        spec_ld_succeed_REG_1;	// lsu.scala:1384:56
  wire [15:0]       _GEN_802 =
    io_core_brupdate_b1_mispredict_mask & stq_0_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_803 =
    io_core_brupdate_b1_mispredict_mask & stq_1_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_804 =
    io_core_brupdate_b1_mispredict_mask & stq_2_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_805 =
    io_core_brupdate_b1_mispredict_mask & stq_3_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_806 =
    io_core_brupdate_b1_mispredict_mask & stq_4_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_807 =
    io_core_brupdate_b1_mispredict_mask & stq_5_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_808 =
    io_core_brupdate_b1_mispredict_mask & stq_6_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_809 =
    io_core_brupdate_b1_mispredict_mask & stq_7_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_810 =
    io_core_brupdate_b1_mispredict_mask & stq_8_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_811 =
    io_core_brupdate_b1_mispredict_mask & stq_9_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_812 =
    io_core_brupdate_b1_mispredict_mask & stq_10_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_813 =
    io_core_brupdate_b1_mispredict_mask & stq_11_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_814 =
    io_core_brupdate_b1_mispredict_mask & stq_12_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_815 =
    io_core_brupdate_b1_mispredict_mask & stq_13_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_816 =
    io_core_brupdate_b1_mispredict_mask & stq_14_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_817 =
    io_core_brupdate_b1_mispredict_mask & stq_15_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_818 =
    io_core_brupdate_b1_mispredict_mask & stq_16_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_819 =
    io_core_brupdate_b1_mispredict_mask & stq_17_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_820 =
    io_core_brupdate_b1_mispredict_mask & stq_18_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_821 =
    io_core_brupdate_b1_mispredict_mask & stq_19_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_822 =
    io_core_brupdate_b1_mispredict_mask & stq_20_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_823 =
    io_core_brupdate_b1_mispredict_mask & stq_21_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_824 =
    io_core_brupdate_b1_mispredict_mask & stq_22_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [15:0]       _GEN_825 =
    io_core_brupdate_b1_mispredict_mask & stq_23_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire              commit_store =
    io_core_commit_valids_0 & io_core_commit_uops_0_uses_stq;	// lsu.scala:1451:49
  wire              commit_load =
    io_core_commit_valids_0 & io_core_commit_uops_0_uses_ldq;	// lsu.scala:1452:49
  wire [4:0]        idx = commit_store ? stq_commit_head : ldq_head;	// lsu.scala:215:29, :219:29, :1451:49, :1453:18
  wire              wrap_12 = stq_commit_head == 5'h17;	// lsu.scala:219:29, util.scala:205:25
  wire [4:0]        _GEN_826 = stq_commit_head + 5'h1;	// lsu.scala:219:29, :305:44, util.scala:206:28
  wire [4:0]        _GEN_827 =
    commit_store ? (wrap_12 ? 5'h0 : _GEN_826) : stq_commit_head;	// lsu.scala:219:29, :1451:49, :1482:31, util.scala:205:25, :206:{10,28}
  wire              wrap_13 = ldq_head == 5'h17;	// lsu.scala:215:29, util.scala:205:25
  wire [4:0]        _GEN_828 = ldq_head + 5'h1;	// lsu.scala:215:29, :305:44, util.scala:206:28
  wire [4:0]        _GEN_829 = commit_load ? (wrap_13 ? 5'h0 : _GEN_828) : ldq_head;	// lsu.scala:215:29, :1452:49, :1486:31, util.scala:205:25, :206:{10,28}
  wire              commit_store_1 =
    io_core_commit_valids_1 & io_core_commit_uops_1_uses_stq;	// lsu.scala:1451:49
  wire              commit_load_1 =
    io_core_commit_valids_1 & io_core_commit_uops_1_uses_ldq;	// lsu.scala:1452:49
  wire [4:0]        idx_1 = commit_store_1 ? _GEN_827 : _GEN_829;	// lsu.scala:1451:49, :1453:18, :1482:31, :1486:31
  wire              wrap_14 = _GEN_827 == 5'h17;	// lsu.scala:1482:31, util.scala:205:25
  wire [4:0]        _GEN_830 = _GEN_827 + 5'h1;	// lsu.scala:305:44, :1482:31, util.scala:206:28
  wire [4:0]        _GEN_831 = commit_store_1 ? (wrap_14 ? 5'h0 : _GEN_830) : _GEN_827;	// lsu.scala:1451:49, :1482:31, util.scala:205:25, :206:{10,28}
  wire              wrap_15 = _GEN_829 == 5'h17;	// lsu.scala:1486:31, util.scala:205:25
  wire [4:0]        _GEN_832 = _GEN_829 + 5'h1;	// lsu.scala:305:44, :1486:31, util.scala:206:28
  wire [4:0]        _GEN_833 = commit_load_1 ? (wrap_15 ? 5'h0 : _GEN_832) : _GEN_829;	// lsu.scala:1452:49, :1486:31, util.scala:205:25, :206:{10,28}
  wire              commit_store_2 =
    io_core_commit_valids_2 & io_core_commit_uops_2_uses_stq;	// lsu.scala:1451:49
  wire              commit_load_2 =
    io_core_commit_valids_2 & io_core_commit_uops_2_uses_ldq;	// lsu.scala:1452:49
  wire [4:0]        idx_2 = commit_store_2 ? _GEN_831 : _GEN_833;	// lsu.scala:1451:49, :1453:18, :1482:31, :1486:31
  `ifndef SYNTHESIS	// lsu.scala:224:10
    always @(posedge clock) begin	// lsu.scala:224:10
      automatic logic        _GEN_834 = ~dis_ld_val & dis_st_val;	// lsu.scala:301:85, :302:85, :304:5, :321:5
      automatic logic        _GEN_835 = ~dis_ld_val_1 & dis_st_val_1;	// lsu.scala:301:85, :302:85, :304:5, :321:5
      automatic logic        _GEN_836 = ~dis_ld_val_2 & dis_st_val_2;	// lsu.scala:301:85, :302:85, :304:5, :321:5
      automatic logic        _GEN_837 =
        ~can_fire_load_incoming_0 & ~will_fire_load_retry_0 & ~will_fire_store_commit_0;	// lsu.scala:441:63, :535:65, :584:6, :766:39, :773:43, :780:45
      automatic logic        _GEN_838 = _GEN_837 & ~will_fire_load_wakeup_0;	// lsu.scala:535:65, :780:45, :794:44
      automatic logic        _GEN_839 =
        io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella;	// lsu.scala:1287:7
      automatic logic        _GEN_840 = ~io_dmem_resp_0_bits_is_hella | reset;	// lsu.scala:1309:{15,16}
      automatic logic        _GEN_841 = ~commit_store & commit_load;	// lsu.scala:1451:49, :1452:49, :1455:5, :1457:31
      automatic logic [31:0] _GEN_842;	// lsu.scala:1458:14
      automatic logic        _GEN_843 = ~commit_store_1 & commit_load_1;	// lsu.scala:1451:49, :1452:49, :1455:5, :1457:31
      automatic logic        _GEN_844 = ~commit_store_2 & commit_load_2;	// lsu.scala:1451:49, :1452:49, :1455:5, :1457:31
      _GEN_842 =
        {{ldq_0_bits_forward_std_val},
         {ldq_0_bits_forward_std_val},
         {ldq_0_bits_forward_std_val},
         {ldq_0_bits_forward_std_val},
         {ldq_0_bits_forward_std_val},
         {ldq_0_bits_forward_std_val},
         {ldq_0_bits_forward_std_val},
         {ldq_0_bits_forward_std_val},
         {ldq_23_bits_forward_std_val},
         {ldq_22_bits_forward_std_val},
         {ldq_21_bits_forward_std_val},
         {ldq_20_bits_forward_std_val},
         {ldq_19_bits_forward_std_val},
         {ldq_18_bits_forward_std_val},
         {ldq_17_bits_forward_std_val},
         {ldq_16_bits_forward_std_val},
         {ldq_15_bits_forward_std_val},
         {ldq_14_bits_forward_std_val},
         {ldq_13_bits_forward_std_val},
         {ldq_12_bits_forward_std_val},
         {ldq_11_bits_forward_std_val},
         {ldq_10_bits_forward_std_val},
         {ldq_9_bits_forward_std_val},
         {ldq_8_bits_forward_std_val},
         {ldq_7_bits_forward_std_val},
         {ldq_6_bits_forward_std_val},
         {ldq_5_bits_forward_std_val},
         {ldq_4_bits_forward_std_val},
         {ldq_3_bits_forward_std_val},
         {ldq_2_bits_forward_std_val},
         {ldq_1_bits_forward_std_val},
         {ldq_0_bits_forward_std_val}};	// lsu.scala:210:16, :1458:14
      if (~(io_core_brupdate_b2_mispredict | _GEN_3 | stq_head == stq_execute_head
            | stq_tail == stq_execute_head | reset)) begin	// lsu.scala:217:29, :218:29, :220:29, :224:{10,42}, :226:20, :227:20
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:224:10
          $error("Assertion failed: stq_execute_head got off track.\n    at lsu.scala:224 assert (io.core.brupdate.b2.mispredict ||\n");	// lsu.scala:224:10
        if (`STOP_COND_)	// lsu.scala:224:10
          $fatal;	// lsu.scala:224:10
      end
      if (dis_ld_val & ~(ldq_tail == io_core_dis_uops_0_bits_ldq_idx | reset)) begin	// lsu.scala:216:29, :301:85, :317:{14,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:317:14
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:317 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");	// lsu.scala:317:14
        if (`STOP_COND_)	// lsu.scala:317:14
          $fatal;	// lsu.scala:317:14
      end
      if (dis_ld_val & ~(~_GEN_99[ldq_tail] | reset)) begin	// lsu.scala:216:29, :301:85, :305:44, :318:{14,15}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:318:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:318 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");	// lsu.scala:318:14
        if (`STOP_COND_)	// lsu.scala:318:14
          $fatal;	// lsu.scala:318:14
      end
      if (_GEN_834 & ~(stq_tail == io_core_dis_uops_0_bits_stq_idx | reset)) begin	// lsu.scala:218:29, :321:5, :329:{14,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:329:14
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:329 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");	// lsu.scala:329:14
        if (`STOP_COND_)	// lsu.scala:329:14
          $fatal;	// lsu.scala:329:14
      end
      if (_GEN_834 & ~(~_GEN_2[stq_tail] | reset)) begin	// lsu.scala:218:29, :224:42, :321:5, :322:39, :330:{14,15}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:330:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:330 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");	// lsu.scala:330:14
        if (`STOP_COND_)	// lsu.scala:330:14
          $fatal;	// lsu.scala:330:14
      end
      if (~(~(dis_ld_val & dis_st_val) | reset)) begin	// lsu.scala:301:85, :302:85, :341:{11,12,25}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:341:11
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:341 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");	// lsu.scala:341:11
        if (`STOP_COND_)	// lsu.scala:341:11
          $fatal;	// lsu.scala:341:11
      end
      if (dis_ld_val_1 & ~(_GEN_100 == io_core_dis_uops_1_bits_ldq_idx | reset)) begin	// lsu.scala:301:85, :317:{14,26}, :333:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:317:14
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:317 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");	// lsu.scala:317:14
        if (`STOP_COND_)	// lsu.scala:317:14
          $fatal;	// lsu.scala:317:14
      end
      if (dis_ld_val_1 & ~(~_GEN_99[_GEN_100] | reset)) begin	// lsu.scala:301:85, :305:44, :318:{14,15}, :333:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:318:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:318 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");	// lsu.scala:318:14
        if (`STOP_COND_)	// lsu.scala:318:14
          $fatal;	// lsu.scala:318:14
      end
      if (_GEN_835 & ~(_GEN_101 == io_core_dis_uops_1_bits_stq_idx | reset)) begin	// lsu.scala:321:5, :329:{14,26}, :338:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:329:14
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:329 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");	// lsu.scala:329:14
        if (`STOP_COND_)	// lsu.scala:329:14
          $fatal;	// lsu.scala:329:14
      end
      if (_GEN_835 & ~(~_GEN_2[_GEN_101] | reset)) begin	// lsu.scala:224:42, :321:5, :322:39, :330:{14,15}, :338:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:330:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:330 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");	// lsu.scala:330:14
        if (`STOP_COND_)	// lsu.scala:330:14
          $fatal;	// lsu.scala:330:14
      end
      if (~(~(dis_ld_val_1 & dis_st_val_1) | reset)) begin	// lsu.scala:301:85, :302:85, :341:{11,12,25}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:341:11
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:341 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");	// lsu.scala:341:11
        if (`STOP_COND_)	// lsu.scala:341:11
          $fatal;	// lsu.scala:341:11
      end
      if (dis_ld_val_2 & ~(_GEN_106 == io_core_dis_uops_2_bits_ldq_idx | reset)) begin	// lsu.scala:301:85, :317:{14,26}, :333:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:317:14
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:317 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");	// lsu.scala:317:14
        if (`STOP_COND_)	// lsu.scala:317:14
          $fatal;	// lsu.scala:317:14
      end
      if (dis_ld_val_2 & ~(~_GEN_99[_GEN_106] | reset)) begin	// lsu.scala:301:85, :305:44, :318:{14,15}, :333:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:318:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:318 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");	// lsu.scala:318:14
        if (`STOP_COND_)	// lsu.scala:318:14
          $fatal;	// lsu.scala:318:14
      end
      if (_GEN_836 & ~(_GEN_107 == io_core_dis_uops_2_bits_stq_idx | reset)) begin	// lsu.scala:321:5, :329:{14,26}, :338:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:329:14
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:329 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");	// lsu.scala:329:14
        if (`STOP_COND_)	// lsu.scala:329:14
          $fatal;	// lsu.scala:329:14
      end
      if (_GEN_836 & ~(~_GEN_2[_GEN_107] | reset)) begin	// lsu.scala:224:42, :321:5, :322:39, :330:{14,15}, :338:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:330:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:330 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");	// lsu.scala:330:14
        if (`STOP_COND_)	// lsu.scala:330:14
          $fatal;	// lsu.scala:330:14
      end
      if (~(~(dis_ld_val_2 & dis_st_val_2) | reset)) begin	// lsu.scala:301:85, :302:85, :341:{11,12,25}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:341:11
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:341 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");	// lsu.scala:341:11
        if (`STOP_COND_)	// lsu.scala:341:11
          $fatal;	// lsu.scala:341:11
      end
      if (~(~(io_core_exe_0_req_valid
              & ~(_GEN_215 | will_fire_std_incoming_0 | will_fire_sfence_0))
            | reset)) begin	// lsu.scala:536:61, :567:{11,12,31,34,93,151}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:567:11
          $error("Assertion failed\n    at lsu.scala:567 assert(!(exe_req(w).valid && !(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) || will_fire_std_incoming(w) || will_fire_sfence(w))))\n");	// lsu.scala:567:11
        if (`STOP_COND_)	// lsu.scala:567:11
          $fatal;	// lsu.scala:567:11
      end
      if (~(~((|hella_state) & hella_req_cmd == 5'h14) | reset)) begin	// lsu.scala:242:38, :243:34, :305:44, :593:{9,10,24,36,53}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:593:9
          $error("Assertion failed: SFENCE through hella interface not supported\n    at lsu.scala:593 assert(!(hella_state =/= h_ready && hella_req.cmd === rocket.M_SFENCE),\n");	// lsu.scala:593:9
        if (`STOP_COND_)	// lsu.scala:593:9
          $fatal;	// lsu.scala:593:9
      end
      if (~(~(~_will_fire_store_commit_0_T_2 & exe_tlb_uop_0_is_fence) | reset)) begin	// lsu.scala:538:31, :576:25, :597:24, :682:{12,13,36}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:682:12
          $error("Assertion failed: Fence is pretending to talk to the TLB\n    at lsu.scala:682 assert (!(dtlb.io.req(w).valid && exe_tlb_uop(w).is_fence), \"Fence is pretending to talk to the TLB\")\n");	// lsu.scala:682:12
        if (`STOP_COND_)	// lsu.scala:682:12
          $fatal;	// lsu.scala:682:12
      end
      if (~(~((can_fire_load_incoming_0 | will_fire_sta_incoming_0
               | will_fire_stad_incoming_0) & io_core_exe_0_req_bits_mxcpt_valid
              & ~_will_fire_store_commit_0_T_2
              & ~(exe_tlb_uop_0_ctrl_is_load | exe_tlb_uop_0_ctrl_is_sta)) | reset)) begin	// lsu.scala:441:63, :534:63, :536:61, :538:31, :576:25, :597:24, :683:{12,13,72}, :684:59, :685:{5,35}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:683:12
          $error("Assertion failed: A uop that's not a load or store-address is throwing a memory exception.\n    at lsu.scala:683 assert (!((will_fire_load_incoming(w) || will_fire_sta_incoming(w) || will_fire_stad_incoming(w)) &&\n");	// lsu.scala:683:12
        if (`STOP_COND_)	// lsu.scala:683:12
          $fatal;	// lsu.scala:683:12
      end
      if (~(exe_tlb_paddr_0 == _dtlb_io_resp_0_paddr | io_core_exe_0_req_bits_sfence_valid
            | reset)) begin	// Cat.scala:30:58, lsu.scala:249:20, :714:{12,30}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:714:12
          $error("Assertion failed: [lsu] paddrs should match.\n    at lsu.scala:714 assert (exe_tlb_paddr(w) === dtlb.io.resp(w).paddr || exe_req(w).bits.sfence.valid, \"[lsu] paddrs should match.\")\n");	// lsu.scala:714:12
        if (`STOP_COND_)	// lsu.scala:714:12
          $fatal;	// lsu.scala:714:12
      end
      if (mem_xcpt_valids_0 & ~(REG | reset)) begin	// lsu.scala:667:32, :718:{13,21}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:718:13
          $error("Assertion failed\n    at lsu.scala:718 assert(RegNext(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) ||\n");	// lsu.scala:718:13
        if (`STOP_COND_)	// lsu.scala:718:13
          $fatal;	// lsu.scala:718:13
      end
      if (mem_xcpt_valids_0
          & ~(mem_xcpt_uops_0_uses_ldq ^ mem_xcpt_uops_0_uses_stq | reset)) begin	// lsu.scala:667:32, :671:32, :721:{13,40}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:721:13
          $error("Assertion failed\n    at lsu.scala:721 assert(mem_xcpt_uops(w).uses_ldq ^ mem_xcpt_uops(w).uses_stq)\n");	// lsu.scala:721:13
        if (`STOP_COND_)	// lsu.scala:721:13
          $fatal;	// lsu.scala:721:13
      end
      if (can_fire_load_incoming_0
          & ~(~_GEN_114[io_core_exe_0_req_bits_uop_ldq_idx] | reset)) begin	// lsu.scala:264:49, :441:63, :772:{13,14}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:772:13
          $error("Assertion failed\n    at lsu.scala:772 assert(!ldq_incoming_e(w).bits.executed)\n");	// lsu.scala:772:13
        if (`STOP_COND_)	// lsu.scala:772:13
          $fatal;	// lsu.scala:772:13
      end
      if (~can_fire_load_incoming_0 & will_fire_load_retry_0
          & ~(~_GEN_114[ldq_retry_idx] | reset)) begin	// lsu.scala:264:49, :415:30, :441:63, :465:79, :535:65, :766:39, :779:{13,14}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:779:13
          $error("Assertion failed\n    at lsu.scala:779 assert(!ldq_retry_e.bits.executed)\n");	// lsu.scala:779:13
        if (`STOP_COND_)	// lsu.scala:779:13
          $fatal;	// lsu.scala:779:13
      end
      if (_GEN_837 & will_fire_load_wakeup_0 & ~(~_GEN_213 & ~_GEN_211 | reset)) begin	// lsu.scala:502:88, :505:31, :506:31, :535:65, :780:45, :801:{13,42}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:801:13
          $error("Assertion failed\n    at lsu.scala:801 assert(!ldq_wakeup_e.bits.executed && !ldq_wakeup_e.bits.addr_is_virtual)\n");	// lsu.scala:801:13
        if (`STOP_COND_)	// lsu.scala:801:13
          $fatal;	// lsu.scala:801:13
      end
      if (_GEN_838 & will_fire_hella_incoming_0 & ~(_GEN_1 | reset)) begin	// lsu.scala:535:65, :794:44, :803:{13,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:803:13
          $error("Assertion failed\n    at lsu.scala:803 assert(hella_state === h_s1)\n");	// lsu.scala:803:13
        if (`STOP_COND_)	// lsu.scala:803:13
          $fatal;	// lsu.scala:803:13
      end
      if (_GEN_838 & ~will_fire_hella_incoming_0 & will_fire_hella_wakeup_0
          & ~(_GEN_0 | reset)) begin	// lsu.scala:535:65, :794:44, :802:47, :820:{13,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:820:13
          $error("Assertion failed\n    at lsu.scala:820 assert(hella_state === h_replay)\n");	// lsu.scala:820:13
        if (`STOP_COND_)	// lsu.scala:820:13
          $fatal;	// lsu.scala:820:13
      end
      if (_GEN_315
          & ~(~(can_fire_load_incoming_0 & _GEN_113[io_core_exe_0_req_bits_uop_ldq_idx])
              | reset)) begin	// lsu.scala:220:29, :264:49, :441:63, :766:39, :773:43, :780:45, :844:{13,14,43}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:844:13
          $error("Assertion failed: [lsu] Incoming load is overwriting a valid address\n    at lsu.scala:844 assert(!(will_fire_load_incoming(w) && ldq_incoming_e(w).bits.addr.valid),\n");	// lsu.scala:844:13
        if (`STOP_COND_)	// lsu.scala:844:13
          $fatal;	// lsu.scala:844:13
      end
      if (_GEN_321
          & ~(~(will_fire_sta_incoming_0 & _GEN_87[io_core_exe_0_req_bits_uop_stq_idx])
              | reset)) begin	// lsu.scala:224:42, :264:49, :536:61, :848:67, :858:{13,14,42}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:858:13
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid address\n    at lsu.scala:858 assert(!(will_fire_sta_incoming(w) && stq_incoming_e(w).bits.addr.valid),\n");	// lsu.scala:858:13
        if (`STOP_COND_)	// lsu.scala:858:13
          $fatal;	// lsu.scala:858:13
      end
      if (_GEN_322 & ~(~_GEN_91[sidx] | reset)) begin	// lsu.scala:224:42, :868:67, :870:21, :873:33, :877:{13,14}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:877:13
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid data entry\n    at lsu.scala:877 assert(!(stq(sidx).bits.data.valid),\n");	// lsu.scala:877:13
        if (`STOP_COND_)	// lsu.scala:877:13
          $fatal;	// lsu.scala:877:13
      end
      if (_GEN_758 & ~(_GEN_759 | _GEN_760 | reset)) begin	// lsu.scala:1287:7, :1288:{15,28,54}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1288:15
          $error("Assertion failed\n    at lsu.scala:1288 assert(hella_state === h_wait || hella_state === h_dead)\n");	// lsu.scala:1288:15
        if (`STOP_COND_)	// lsu.scala:1288:15
          $fatal;	// lsu.scala:1288:15
      end
      if (_GEN_839 & io_dmem_nack_0_bits_uop_uses_ldq
          & ~(_GEN_114[io_dmem_nack_0_bits_uop_ldq_idx] | reset)) begin	// lsu.scala:264:49, :1287:7, :1292:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1292:15
          $error("Assertion failed\n    at lsu.scala:1292 assert(ldq(io.dmem.nack(w).bits.uop.ldq_idx).bits.executed)\n");	// lsu.scala:1292:15
        if (`STOP_COND_)	// lsu.scala:1292:15
          $fatal;	// lsu.scala:1292:15
      end
      if (_GEN_839 & ~io_dmem_nack_0_bits_uop_uses_ldq
          & ~(io_dmem_nack_0_bits_uop_uses_stq | reset)) begin	// lsu.scala:1287:7, :1291:7, :1298:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1298:15
          $error("Assertion failed\n    at lsu.scala:1298 assert(io.dmem.nack(w).bits.uop.uses_stq)\n");	// lsu.scala:1298:15
        if (`STOP_COND_)	// lsu.scala:1298:15
          $fatal;	// lsu.scala:1298:15
      end
      if (_GEN_785 & ~_GEN_840) begin	// lsu.scala:1308:7, :1309:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1309:15
          $error("Assertion failed\n    at lsu.scala:1309 assert(!io.dmem.resp(w).bits.is_hella)\n");	// lsu.scala:1309:15
        if (`STOP_COND_)	// lsu.scala:1309:15
          $fatal;	// lsu.scala:1309:15
      end
      if (_GEN_785 & ~(send_iresp ^ send_fresp | reset)) begin	// lsu.scala:1308:7, :1311:58, :1312:58, :1321:{15,27}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1321:15
          $error("Assertion failed\n    at lsu.scala:1321 assert(send_iresp ^ send_fresp)\n");	// lsu.scala:1321:15
        if (`STOP_COND_)	// lsu.scala:1321:15
          $fatal;	// lsu.scala:1321:15
      end
      if (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
          & io_dmem_resp_0_bits_uop_uses_stq & ~_GEN_840) begin	// lsu.scala:1308:7, :1309:15, :1329:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1329:15
          $error("Assertion failed\n    at lsu.scala:1329 assert(!io.dmem.resp(w).bits.is_hella)\n");	// lsu.scala:1329:15
        if (`STOP_COND_)	// lsu.scala:1329:15
          $fatal;	// lsu.scala:1329:15
      end
      if (~(~((|_GEN_802) & stq_0_valid & stq_0_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_803) & stq_1_valid & stq_1_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_804) & stq_2_valid & stq_2_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_805) & stq_3_valid & stq_3_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_806) & stq_4_valid & stq_4_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_807) & stq_5_valid & stq_5_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_808) & stq_6_valid & stq_6_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_809) & stq_7_valid & stq_7_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_810) & stq_8_valid & stq_8_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_811) & stq_9_valid & stq_9_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_812) & stq_10_valid & stq_10_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_813) & stq_11_valid & stq_11_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_814) & stq_12_valid & stq_12_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_815) & stq_13_valid & stq_13_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_816) & stq_14_valid & stq_14_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_817) & stq_15_valid & stq_15_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_818) & stq_16_valid & stq_16_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_819) & stq_17_valid & stq_17_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_820) & stq_18_valid & stq_18_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_821) & stq_19_valid & stq_19_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_822) & stq_20_valid & stq_20_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_823) & stq_21_valid & stq_21_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_824) & stq_22_valid & stq_22_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_825) & stq_23_valid & stq_23_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (_GEN_841 & ~(_GEN_99[idx] | reset)) begin	// lsu.scala:305:44, :1453:18, :1457:31, :1458:14
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1458:14
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1458 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");	// lsu.scala:1458:14
        if (`STOP_COND_)	// lsu.scala:1458:14
          $fatal;	// lsu.scala:1458:14
      end
      if (_GEN_841 & ~((_GEN_114[idx] | _GEN_842[idx]) & _GEN_214[idx] | reset)) begin	// lsu.scala:264:49, :502:88, :1453:18, :1457:31, :1458:14, :1459:{14,39,73}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1459:14
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1459 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");	// lsu.scala:1459:14
        if (`STOP_COND_)	// lsu.scala:1459:14
          $fatal;	// lsu.scala:1459:14
      end
      if (_GEN_843 & ~(_GEN_99[idx_1] | reset)) begin	// lsu.scala:305:44, :1453:18, :1457:31, :1458:14
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1458:14
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1458 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");	// lsu.scala:1458:14
        if (`STOP_COND_)	// lsu.scala:1458:14
          $fatal;	// lsu.scala:1458:14
      end
      if (_GEN_843
          & ~((_GEN_114[idx_1] | _GEN_842[idx_1]) & _GEN_214[idx_1] | reset)) begin	// lsu.scala:264:49, :502:88, :1453:18, :1457:31, :1458:14, :1459:{14,39,73}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1459:14
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1459 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");	// lsu.scala:1459:14
        if (`STOP_COND_)	// lsu.scala:1459:14
          $fatal;	// lsu.scala:1459:14
      end
      if (_GEN_844 & ~(_GEN_99[idx_2] | reset)) begin	// lsu.scala:305:44, :1453:18, :1457:31, :1458:14
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1458:14
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1458 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");	// lsu.scala:1458:14
        if (`STOP_COND_)	// lsu.scala:1458:14
          $fatal;	// lsu.scala:1458:14
      end
      if (_GEN_844
          & ~((_GEN_114[idx_2] | _GEN_842[idx_2]) & _GEN_214[idx_2] | reset)) begin	// lsu.scala:264:49, :502:88, :1453:18, :1457:31, :1458:14, :1459:{14,39,73}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1459:14
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1459 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");	// lsu.scala:1459:14
        if (`STOP_COND_)	// lsu.scala:1459:14
          $fatal;	// lsu.scala:1459:14
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire              _GEN_845 = _GEN_58[stq_head];	// lsu.scala:217:29, :224:42, :1494:29
  wire [31:0]       _GEN_846 =
    {{stq_0_bits_succeeded},
     {stq_0_bits_succeeded},
     {stq_0_bits_succeeded},
     {stq_0_bits_succeeded},
     {stq_0_bits_succeeded},
     {stq_0_bits_succeeded},
     {stq_0_bits_succeeded},
     {stq_0_bits_succeeded},
     {stq_23_bits_succeeded},
     {stq_22_bits_succeeded},
     {stq_21_bits_succeeded},
     {stq_20_bits_succeeded},
     {stq_19_bits_succeeded},
     {stq_18_bits_succeeded},
     {stq_17_bits_succeeded},
     {stq_16_bits_succeeded},
     {stq_15_bits_succeeded},
     {stq_14_bits_succeeded},
     {stq_13_bits_succeeded},
     {stq_12_bits_succeeded},
     {stq_11_bits_succeeded},
     {stq_10_bits_succeeded},
     {stq_9_bits_succeeded},
     {stq_8_bits_succeeded},
     {stq_7_bits_succeeded},
     {stq_6_bits_succeeded},
     {stq_5_bits_succeeded},
     {stq_4_bits_succeeded},
     {stq_3_bits_succeeded},
     {stq_2_bits_succeeded},
     {stq_1_bits_succeeded},
     {stq_0_bits_succeeded}};	// lsu.scala:211:16, :1494:29
  wire              _GEN_847 = _GEN_2[stq_head] & _GEN_94[stq_head];	// lsu.scala:217:29, :224:42, :1494:29
  wire              _GEN_848 = _GEN_845 & ~io_dmem_ordered;	// lsu.scala:1494:29, :1496:{43,46}
  assign store_needs_order = _GEN_847 & _GEN_848;	// lsu.scala:1494:29, :1495:3, :1496:{43,64}
  wire              clear_store =
    _GEN_847 & (_GEN_845 ? io_dmem_ordered : _GEN_846[stq_head]);	// lsu.scala:217:29, :1494:29, :1495:3, :1500:{17,23}
  wire              _GEN_849 = hella_state == 3'h3;	// lsu.scala:242:38, :1548:19, :1550:28
  wire              _GEN_850 = ~(|hella_state) | _GEN_1;	// lsu.scala:242:38, :593:24, :803:26, :1524:27, :1527:{21,34}, :1533:38, :1550:43
  wire              _GEN_851 = hella_state == 3'h2;	// lsu.scala:242:38, :1546:19, :1553:28
  wire              _GEN_852 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_is_hella;	// lsu.scala:1562:35
  assign _GEN = ~(~(|hella_state) | _GEN_1 | _GEN_849 | _GEN_851 | _GEN_759);	// lsu.scala:242:38, :593:24, :803:26, :1288:28, :1527:{21,34}, :1533:38, :1550:{28,43}, :1553:{28,38}, :1560:40, :1576:42
  always @(posedge clock) begin
    automatic logic [31:0] _ldq_23_bits_st_dep_mask_T;	// lsu.scala:260:71
    automatic logic [23:0] _GEN_853;	// lsu.scala:260:33
    automatic logic [23:0] _GEN_854;	// lsu.scala:260:33
    automatic logic        _GEN_855;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_856;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_857;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_858;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_859;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_860;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_861;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_862;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_863;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_864;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_865;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_866;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_867;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_868;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_869;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_870;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_871;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_872;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_873;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_874;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_875;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_876;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_877;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_878;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_879;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_880;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_881;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_882;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_883;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_884;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_885;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_886;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_887;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_888;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_889;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_890;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_891;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_892;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_893;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_894;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_895;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_896;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_897;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_898;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_899;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_900;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_901;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_902;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_903;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_904;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_905;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_906;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_907;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_908;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_909;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_910;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_911;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_912;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_913;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_914;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_915;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_916;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_917;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_918;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_919;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_920;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_921;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_922;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_923;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_924;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_925;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_926;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic [31:0] _GEN_927;	// lsu.scala:336:72
    automatic logic [23:0] _GEN_928;	// lsu.scala:336:31
    automatic logic        _GEN_929 = _GEN_100 == 5'h0;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_930;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_931 = _GEN_100 == 5'h1;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_932;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_933 = _GEN_100 == 5'h2;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_934;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_935 = _GEN_100 == 5'h3;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_936;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_937 = _GEN_100 == 5'h4;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_938;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_939 = _GEN_100 == 5'h5;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_940;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_941 = _GEN_100 == 5'h6;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_942;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_943 = _GEN_100 == 5'h7;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_944;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_945 = _GEN_100 == 5'h8;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_946;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_947 = _GEN_100 == 5'h9;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_948;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_949 = _GEN_100 == 5'hA;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_950;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_951 = _GEN_100 == 5'hB;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_952;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_953 = _GEN_100 == 5'hC;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_954;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_955 = _GEN_100 == 5'hD;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_956;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_957 = _GEN_100 == 5'hE;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_958;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_959 = _GEN_100 == 5'hF;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_960;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_961 = _GEN_100 == 5'h10;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_962;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_963 = _GEN_100 == 5'h11;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_964;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_965 = _GEN_100 == 5'h12;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_966;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_967 = _GEN_100 == 5'h13;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_968;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_969 = _GEN_100 == 5'h14;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_970;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_971 = _GEN_100 == 5'h15;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_972;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_973 = _GEN_100 == 5'h16;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_974;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_975 = _GEN_100 == 5'h17;	// lsu.scala:305:44, :333:21, util.scala:205:25
    automatic logic        _GEN_976;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_977;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_978;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_979;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_980;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_981;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_982;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_983;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_984;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_985;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_986;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_987;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_988;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_989;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_990;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_991;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_992;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_993;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_994;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_995;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_996;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_997;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_998;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_999;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_1000;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_1001;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1002;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1003;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1004;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1005;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1006;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1007;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1008;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1009;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1010;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1011;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1012;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1013;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1014;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1015;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1016;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1017;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1018;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1019;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1020;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1021;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1022;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1023;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1024;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_1025;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1026;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1027;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1028;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1029;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1030;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1031;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1032;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1033;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1034;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1035;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1036;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1037;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1038;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1039;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1040;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1041;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1042;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1043;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1044;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1045;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1046;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1047;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1048;	// lsu.scala:304:5, :321:5
    automatic logic [31:0] _GEN_1049 = 32'h1 << _GEN_101;	// lsu.scala:260:71, :336:72, :338:21
    automatic logic [23:0] _GEN_1050;	// lsu.scala:336:31
    automatic logic        _GEN_1051;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1052;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1053;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1054;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1055;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1056;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1057;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1058;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1059;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1060;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1061;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1062;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1063;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1064;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1065;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1066;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1067;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1068;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1069;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1070;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1071;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1072;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1073;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1074;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1075;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1076;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1077;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1078;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1079;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1080;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1081;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1082;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1083;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1084;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1085;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1086;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1087;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1088;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1089;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1090;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1091;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1092;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1093;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1094;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1095;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1096;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1097;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1098;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_1099;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1100;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1101;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1102;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1103;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1104;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1105;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1106;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1107;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1108;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1109;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1110;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1111;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1112;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1113;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1114;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1115;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1116;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1117;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1118;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1119;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1120;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1121;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1122;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_1123;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1124;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1125;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1126;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1127;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1128;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1129;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1130;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1131;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1132;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1133;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1134;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1135;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1136;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1137;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1138;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1139;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1140;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1141;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1142;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1143;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1144;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1145;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1146;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_1147 = dis_st_val_2 & _GEN_107 == 5'h0;	// lsu.scala:302:85, :304:5, :321:5, :322:39, :338:21
    automatic logic        _GEN_1148;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1149 = dis_st_val_2 & _GEN_107 == 5'h1;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1150;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1151 = dis_st_val_2 & _GEN_107 == 5'h2;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1152;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1153 = dis_st_val_2 & _GEN_107 == 5'h3;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1154;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1155 = dis_st_val_2 & _GEN_107 == 5'h4;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1156;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1157 = dis_st_val_2 & _GEN_107 == 5'h5;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1158;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1159 = dis_st_val_2 & _GEN_107 == 5'h6;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1160;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1161 = dis_st_val_2 & _GEN_107 == 5'h7;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1162;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1163 = dis_st_val_2 & _GEN_107 == 5'h8;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1164;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1165 = dis_st_val_2 & _GEN_107 == 5'h9;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1166;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1167 = dis_st_val_2 & _GEN_107 == 5'hA;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1168;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1169 = dis_st_val_2 & _GEN_107 == 5'hB;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1170;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1171 = dis_st_val_2 & _GEN_107 == 5'hC;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1172;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1173 = dis_st_val_2 & _GEN_107 == 5'hD;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1174;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1175 = dis_st_val_2 & _GEN_107 == 5'hE;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1176;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1177 = dis_st_val_2 & _GEN_107 == 5'hF;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1178;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1179 = dis_st_val_2 & _GEN_107 == 5'h10;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1180;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1181 = dis_st_val_2 & _GEN_107 == 5'h11;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1182;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1183 = dis_st_val_2 & _GEN_107 == 5'h12;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1184;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1185 = dis_st_val_2 & _GEN_107 == 5'h13;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1186;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1187 = dis_st_val_2 & _GEN_107 == 5'h14;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1188;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1189 = dis_st_val_2 & _GEN_107 == 5'h15;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1190;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1191 = dis_st_val_2 & _GEN_107 == 5'h16;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    automatic logic        _GEN_1192;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1193 = dis_st_val_2 & _GEN_107 == 5'h17;	// lsu.scala:302:85, :304:5, :321:5, :322:39, :338:21, util.scala:205:25
    automatic logic        _GEN_1194;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1195;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1196;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1197;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1198;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1199;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1200;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1201;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1202;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1203;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1204;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1205;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1206;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1207;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1208;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1209;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1210;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1211;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1212;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1213;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1214;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1215;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1216;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1217;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1218;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1219;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1220;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1221;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1222;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1223;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1224;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1225;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1226;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1227;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1228;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1229;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1230;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1231;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1232;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1233;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1234;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1235;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1236;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1237;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1238;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1239;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1240;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1241;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_1242;	// lsu.scala:304:5, :321:5
    automatic logic        ldq_retry_idx_block;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_2;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_1;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_5;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_2;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_8;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_3;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_11;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_4;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_14;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_5;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_17;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_6;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_20;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_7;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_23;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_8;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_26;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_9;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_29;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_10;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_32;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_11;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_35;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_12;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_38;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_13;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_41;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_14;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_44;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_15;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_47;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_16;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_50;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_17;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_53;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_18;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_56;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_19;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_59;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_20;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_62;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_21;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_65;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_22;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_68;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_23;	// lsu.scala:417:36
    automatic logic        _temp_bits_T;	// util.scala:351:72
    automatic logic        _temp_bits_T_2;	// util.scala:351:72
    automatic logic        _temp_bits_T_4;	// util.scala:351:72
    automatic logic        _temp_bits_T_6;	// util.scala:351:72
    automatic logic        _temp_bits_T_8;	// util.scala:351:72
    automatic logic        _temp_bits_T_10;	// util.scala:351:72
    automatic logic        _temp_bits_T_12;	// util.scala:351:72
    automatic logic        _temp_bits_T_14;	// util.scala:351:72
    automatic logic        _temp_bits_T_16;	// util.scala:351:72
    automatic logic        _temp_bits_T_18;	// util.scala:351:72
    automatic logic        _temp_bits_T_20;	// util.scala:351:72
    automatic logic        _temp_bits_T_22;	// util.scala:351:72
    automatic logic        _temp_bits_T_24;	// util.scala:351:72
    automatic logic        _temp_bits_T_26;	// util.scala:351:72
    automatic logic        _temp_bits_T_28;	// util.scala:351:72
    automatic logic        _temp_bits_T_32;	// util.scala:351:72
    automatic logic        _temp_bits_T_34;	// util.scala:351:72
    automatic logic        _temp_bits_T_36;	// util.scala:351:72
    automatic logic        _temp_bits_T_38;	// util.scala:351:72
    automatic logic        _temp_bits_T_40;	// util.scala:351:72
    automatic logic        _temp_bits_T_42;	// util.scala:351:72
    automatic logic        _temp_bits_T_44;	// util.scala:351:72
    automatic logic        _temp_bits_T_46;	// util.scala:351:72
    automatic logic        _stq_retry_idx_T;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_1;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_2;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_3;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_4;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_5;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_6;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_7;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_8;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_9;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_10;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_11;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_12;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_13;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_14;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_15;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_16;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_17;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_18;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_19;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_20;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_21;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_22;	// lsu.scala:424:18
    automatic logic        _ldq_wakeup_idx_T_7;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_15;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_23;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_31;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_39;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_47;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_55;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_63;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_71;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_79;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_87;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_95;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_103;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_111;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_119;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_127;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_135;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_143;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_151;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_159;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_167;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_175;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_183;	// lsu.scala:433:71
    automatic logic        ma_ld_0 =
      can_fire_load_incoming_0 & io_core_exe_0_req_bits_mxcpt_valid;	// lsu.scala:441:63, :659:56
    automatic logic        ma_st_0;	// lsu.scala:660:87
    automatic logic        pf_ld_0;	// lsu.scala:661:75
    automatic logic        pf_st_0;	// lsu.scala:662:75
    automatic logic        ae_ld_0;	// lsu.scala:663:75
    automatic logic        dmem_req_fire_0;	// lsu.scala:752:55
    automatic logic [4:0]  ldq_idx;	// lsu.scala:837:24
    automatic logic        _GEN_1243;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1244;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1245;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1246;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1247;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1248;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1249;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1250;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1251;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1252;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1253;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1254;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1255;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1256;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1257;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1258;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1259;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1260;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1261;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1262;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1263;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1264;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1265;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1266;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1267;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1268;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1269;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1270;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1271;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1272;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1273;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1274;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1275;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1276;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1277;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1278;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1279;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1280;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1281;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1282;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1283;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1284;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1285;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1286;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1287;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1288;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1289;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_1290;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:842:71
    automatic logic [4:0]  stq_idx;	// lsu.scala:850:24
    automatic logic        _GEN_1291;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1292;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1293;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1294;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1295;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1296;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1297;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1298;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1299;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1300;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1301;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1302;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1303;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1304;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1305;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1306;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1307;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1308;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1309;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1310;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1311;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1312;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1313;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1314;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1315;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1316;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1317;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1318;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1319;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1320;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1321;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1322;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1323;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1324;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1325;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1326;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1327;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1328;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1329;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1330;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1331;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1332;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1333;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1334;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1335;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1336;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1337;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1338;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_1339 = _GEN_322 & sidx == 5'h0;	// lsu.scala:304:5, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1340;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1341 = _GEN_322 & sidx == 5'h1;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1342;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1343 = _GEN_322 & sidx == 5'h2;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1344;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1345 = _GEN_322 & sidx == 5'h3;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1346;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1347 = _GEN_322 & sidx == 5'h4;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1348;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1349 = _GEN_322 & sidx == 5'h5;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1350;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1351 = _GEN_322 & sidx == 5'h6;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1352;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1353 = _GEN_322 & sidx == 5'h7;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1354;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1355 = _GEN_322 & sidx == 5'h8;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1356;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1357 = _GEN_322 & sidx == 5'h9;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1358;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1359 = _GEN_322 & sidx == 5'hA;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1360;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1361 = _GEN_322 & sidx == 5'hB;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1362;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1363 = _GEN_322 & sidx == 5'hC;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1364;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1365 = _GEN_322 & sidx == 5'hD;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1366;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1367 = _GEN_322 & sidx == 5'hE;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1368;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1369 = _GEN_322 & sidx == 5'hF;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1370;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1371 = _GEN_322 & sidx == 5'h10;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1372;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1373 = _GEN_322 & sidx == 5'h11;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1374;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1375 = _GEN_322 & sidx == 5'h12;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1376;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1377 = _GEN_322 & sidx == 5'h13;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1378;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1379 = _GEN_322 & sidx == 5'h14;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1380;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1381 = _GEN_322 & sidx == 5'h15;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1382;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1383 = _GEN_322 & sidx == 5'h16;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_1384;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_1385 = _GEN_322 & sidx == 5'h17;	// lsu.scala:304:5, :868:67, :869:5, :870:21, :873:33, util.scala:205:25
    automatic logic        _GEN_1386;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _fired_std_incoming_T =
      (io_core_brupdate_b1_mispredict_mask & io_core_exe_0_req_bits_uop_br_mask) == 16'h0;	// util.scala:118:{51,59}
    automatic logic [15:0] _mem_stq_retry_e_out_valid_T =
      io_core_brupdate_b1_mispredict_mask & _GEN_205;	// lsu.scala:478:79, util.scala:118:51
    automatic logic [4:0]  l_forward_stq_idx;	// lsu.scala:1077:32
    automatic logic        _GEN_1387;	// lsu.scala:1106:39
    automatic logic        _GEN_1388;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_24;	// lsu.scala:1091:36, :1102:37
    automatic logic        _GEN_1389 = lcam_ldq_idx_0 == 5'h1;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1390 = lcam_ldq_idx_0 == 5'h2;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1391 = lcam_ldq_idx_0 == 5'h3;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1392 = lcam_ldq_idx_0 == 5'h4;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1393 = lcam_ldq_idx_0 == 5'h5;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1394 = lcam_ldq_idx_0 == 5'h6;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1395 = lcam_ldq_idx_0 == 5'h7;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1396 = lcam_ldq_idx_0 == 5'h8;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1397 = lcam_ldq_idx_0 == 5'h9;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1398 = lcam_ldq_idx_0 == 5'hA;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1399 = lcam_ldq_idx_0 == 5'hB;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1400 = lcam_ldq_idx_0 == 5'hC;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1401 = lcam_ldq_idx_0 == 5'hD;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1402 = lcam_ldq_idx_0 == 5'hE;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1403 = lcam_ldq_idx_0 == 5'hF;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1404 = lcam_ldq_idx_0 == 5'h10;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1405 = lcam_ldq_idx_0 == 5'h11;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1406 = lcam_ldq_idx_0 == 5'h12;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1407 = lcam_ldq_idx_0 == 5'h13;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1408 = lcam_ldq_idx_0 == 5'h14;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1409 = lcam_ldq_idx_0 == 5'h15;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1410 = lcam_ldq_idx_0 == 5'h16;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_1411 = lcam_ldq_idx_0 == 5'h17;	// lsu.scala:1036:26, :1130:48, util.scala:205:25
    automatic logic [4:0]  l_forward_stq_idx_1;	// lsu.scala:1077:32
    automatic logic        _GEN_1412;	// lsu.scala:1106:39
    automatic logic        _GEN_1413;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_25;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_2;	// lsu.scala:1077:32
    automatic logic        _GEN_1414;	// lsu.scala:1106:39
    automatic logic        _GEN_1415;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_26;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_3;	// lsu.scala:1077:32
    automatic logic        _GEN_1416;	// lsu.scala:1106:39
    automatic logic        _GEN_1417;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_27;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_4;	// lsu.scala:1077:32
    automatic logic        _GEN_1418;	// lsu.scala:1106:39
    automatic logic        _GEN_1419;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_28;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_5;	// lsu.scala:1077:32
    automatic logic        _GEN_1420;	// lsu.scala:1106:39
    automatic logic        _GEN_1421;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_29;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_6;	// lsu.scala:1077:32
    automatic logic        _GEN_1422;	// lsu.scala:1106:39
    automatic logic        _GEN_1423;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_30;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_7;	// lsu.scala:1077:32
    automatic logic        _GEN_1424;	// lsu.scala:1106:39
    automatic logic        _GEN_1425;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_31;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_8;	// lsu.scala:1077:32
    automatic logic        _GEN_1426;	// lsu.scala:1106:39
    automatic logic        _GEN_1427;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_32;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_9;	// lsu.scala:1077:32
    automatic logic        _GEN_1428;	// lsu.scala:1106:39
    automatic logic        _GEN_1429;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_33;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_10;	// lsu.scala:1077:32
    automatic logic        _GEN_1430;	// lsu.scala:1106:39
    automatic logic        _GEN_1431;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_34;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_11;	// lsu.scala:1077:32
    automatic logic        _GEN_1432;	// lsu.scala:1106:39
    automatic logic        _GEN_1433;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_35;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_12;	// lsu.scala:1077:32
    automatic logic        _GEN_1434;	// lsu.scala:1106:39
    automatic logic        _GEN_1435;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_36;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_13;	// lsu.scala:1077:32
    automatic logic        _GEN_1436;	// lsu.scala:1106:39
    automatic logic        _GEN_1437;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_37;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_14;	// lsu.scala:1077:32
    automatic logic        _GEN_1438;	// lsu.scala:1106:39
    automatic logic        _GEN_1439;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_38;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_15;	// lsu.scala:1077:32
    automatic logic        _GEN_1440;	// lsu.scala:1106:39
    automatic logic        _GEN_1441;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_39;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_16;	// lsu.scala:1077:32
    automatic logic        _GEN_1442;	// lsu.scala:1106:39
    automatic logic        _GEN_1443;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_40;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_17;	// lsu.scala:1077:32
    automatic logic        _GEN_1444;	// lsu.scala:1106:39
    automatic logic        _GEN_1445;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_41;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_18;	// lsu.scala:1077:32
    automatic logic        _GEN_1446;	// lsu.scala:1106:39
    automatic logic        _GEN_1447;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_42;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_19;	// lsu.scala:1077:32
    automatic logic        _GEN_1448;	// lsu.scala:1106:39
    automatic logic        _GEN_1449;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_43;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_20;	// lsu.scala:1077:32
    automatic logic        _GEN_1450;	// lsu.scala:1106:39
    automatic logic        _GEN_1451;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_44;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_21;	// lsu.scala:1077:32
    automatic logic        _GEN_1452;	// lsu.scala:1106:39
    automatic logic        _GEN_1453;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_45;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_22;	// lsu.scala:1077:32
    automatic logic        _GEN_1454;	// lsu.scala:1106:39
    automatic logic        _GEN_1455;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_46;	// lsu.scala:1091:36, :1102:37
    automatic logic [4:0]  l_forward_stq_idx_23;	// lsu.scala:1077:32
    automatic logic        _GEN_1456;	// lsu.scala:1106:39
    automatic logic        _GEN_1457;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_47;	// lsu.scala:1091:36, :1102:37
    automatic logic        _GEN_1458;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1459;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1460;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1461;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1462;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1463;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1464;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1465;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1466;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1467;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1468;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1469;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1470;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1471;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1472;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1473;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1474;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1475;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1476;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1477;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1478;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1479;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1480;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1481;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        ldst_forward_matches_0_0 = _GEN_592 & _GEN_594;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9
    automatic logic        _GEN_1482 = _GEN_594 | _GEN_595;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1483;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1484;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1485;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1486;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1487;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1488;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1489;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1490;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1491;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1492;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1493;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1494;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1495;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1496;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1497;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1498;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1499;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1500;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1501;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1502;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1503;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1504;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1505;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1506;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1507 = _GEN_601 | _GEN_602;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1508;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1509;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1510;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1511;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1512;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1513;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1514;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1515;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1516;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1517;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1518;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1519;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1520;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1521;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1522;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1523;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1524;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1525;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1526;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1527;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1528;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1529;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1530;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1531;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1532 = _GEN_608 | _GEN_609;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1533;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1534;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1535;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1536;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1537;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1538;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1539;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1540;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1541;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1542;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1543;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1544;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1545;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1546;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1547;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1548;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1549;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1550;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1551;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1552;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1553;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1554;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1555;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1556;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1557 = _GEN_615 | _GEN_616;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1558;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1559;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1560;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1561;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1562;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1563;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1564;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1565;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1566;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1567;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1568;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1569;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1570;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1571;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1572;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1573;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1574;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1575;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1576;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1577;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1578;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1579;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1580;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1581;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1582 = _GEN_622 | _GEN_623;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1583;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1584;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1585;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1586;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1587;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1588;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1589;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1590;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1591;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1592;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1593;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1594;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1595;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1596;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1597;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1598;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1599;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1600;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1601;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1602;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1603;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1604;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1605;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1606;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1607 = _GEN_629 | _GEN_630;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1608;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1609;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1610;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1611;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1612;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1613;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1614;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1615;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1616;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1617;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1618;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1619;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1620;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1621;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1622;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1623;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1624;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1625;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1626;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1627;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1628;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1629;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1630;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1631;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1632 = _GEN_636 | _GEN_637;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1633;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1634;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1635;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1636;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1637;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1638;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1639;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1640;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1641;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1642;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1643;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1644;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1645;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1646;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1647;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1648;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1649;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1650;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1651;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1652;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1653;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1654;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1655;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1656;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1657 = _GEN_643 | _GEN_644;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1658;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1659;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1660;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1661;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1662;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1663;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1664;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1665;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1666;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1667;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1668;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1669;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1670;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1671;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1672;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1673;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1674;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1675;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1676;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1677;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1678;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1679;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1680;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1681;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1682 = _GEN_650 | _GEN_651;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1683;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1684;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1685;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1686;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1687;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1688;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1689;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1690;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1691;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1692;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1693;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1694;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1695;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1696;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1697;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1698;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1699;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1700;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1701;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1702;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1703;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1704;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1705;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1706;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1707 = _GEN_657 | _GEN_658;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1708;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1709;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1710;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1711;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1712;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1713;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1714;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1715;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1716;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1717;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1718;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1719;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1720;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1721;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1722;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1723;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1724;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1725;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1726;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1727;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1728;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1729;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1730;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1731;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1732 = _GEN_664 | _GEN_665;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1733;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1734;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1735;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1736;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1737;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1738;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1739;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1740;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1741;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1742;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1743;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1744;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1745;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1746;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1747;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1748;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1749;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1750;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1751;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1752;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1753;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1754;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1755;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1756;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1757 = _GEN_671 | _GEN_672;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1758;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1759;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1760;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1761;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1762;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1763;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1764;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1765;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1766;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1767;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1768;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1769;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1770;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1771;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1772;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1773;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1774;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1775;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1776;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1777;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1778;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1779;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1780;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1781;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1782 = _GEN_678 | _GEN_679;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1783;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1784;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1785;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1786;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1787;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1788;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1789;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1790;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1791;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1792;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1793;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1794;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1795;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1796;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1797;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1798;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1799;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1800;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1801;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1802;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1803;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1804;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1805;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1806;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1807 = _GEN_685 | _GEN_686;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1808;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1809;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1810;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1811;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1812;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1813;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1814;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1815;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1816;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1817;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1818;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1819;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1820;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1821;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1822;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1823;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1824;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1825;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1826;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1827;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1828;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1829;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1830;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1831;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1832 = _GEN_692 | _GEN_693;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1833;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1834;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1835;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1836;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1837;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1838;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1839;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1840;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1841;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1842;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1843;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1844;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1845;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1846;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1847;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1848;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1849;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1850;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1851;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1852;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1853;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1854;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1855;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1856;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1857 = _GEN_699 | _GEN_700;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1858;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1859;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1860;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1861;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1862;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1863;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1864;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1865;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1866;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1867;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1868;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1869;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1870;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1871;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1872;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1873;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1874;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1875;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1876;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1877;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1878;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1879;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1880;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1881;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1882 = _GEN_706 | _GEN_707;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1883;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1884;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1885;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1886;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1887;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1888;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1889;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1890;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1891;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1892;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1893;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1894;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1895;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1896;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1897;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1898;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1899;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1900;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1901;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1902;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1903;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1904;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1905;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1906;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1907 = _GEN_713 | _GEN_714;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1908;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1909;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1910;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1911;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1912;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1913;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1914;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1915;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1916;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1917;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1918;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1919;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1920;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1921;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1922;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1923;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1924;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1925;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1926;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1927;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1928;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1929;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1930;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1931;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1932 = _GEN_720 | _GEN_721;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1933;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1934;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1935;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1936;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1937;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1938;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1939;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1940;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1941;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1942;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1943;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1944;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1945;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1946;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1947;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1948;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1949;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1950;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1951;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1952;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1953;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1954;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1955;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1956;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1957 = _GEN_727 | _GEN_728;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1958;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1959;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1960;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1961;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1962;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1963;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1964;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1965;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1966;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1967;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1968;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1969;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1970;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1971;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1972;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1973;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1974;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1975;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1976;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1977;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1978;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1979;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1980;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1981;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1982 = _GEN_734 | _GEN_735;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1983;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1984;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1985;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1986;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1987;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1988;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1989;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1990;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1991;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1992;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1993;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1994;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1995;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1996;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1997;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1998;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1999;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2000;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2001;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2002;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2003;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2004;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2005;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2006;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2007 = _GEN_741 | _GEN_742;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_2008;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2009;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2010;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2011;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2012;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2013;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2014;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2015;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2016;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2017;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2018;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2019;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2020;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2021;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2022;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2023;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2024;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2025;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2026;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2027;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2028;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2029;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2030;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2031;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2032 = _GEN_748 | _GEN_749;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_2033;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2034;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2035;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2036;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2037;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2038;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2039;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2040;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2041;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2042;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2043;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2044;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2045;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2046;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2047;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2048;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2049;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2050;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2051;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2052;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2053;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2054;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2055;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2056;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_2057 = _GEN_755 | _GEN_756;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic [31:0] _GEN_2058 =
      {{ldst_forward_matches_0_0},
       {ldst_forward_matches_0_0},
       {ldst_forward_matches_0_0},
       {ldst_forward_matches_0_0},
       {ldst_forward_matches_0_0},
       {ldst_forward_matches_0_0},
       {ldst_forward_matches_0_0},
       {ldst_forward_matches_0_0},
       {_GEN_753 & _GEN_755},
       {_GEN_746 & _GEN_748},
       {_GEN_739 & _GEN_741},
       {_GEN_732 & _GEN_734},
       {_GEN_725 & _GEN_727},
       {_GEN_718 & _GEN_720},
       {_GEN_711 & _GEN_713},
       {_GEN_704 & _GEN_706},
       {_GEN_697 & _GEN_699},
       {_GEN_690 & _GEN_692},
       {_GEN_683 & _GEN_685},
       {_GEN_676 & _GEN_678},
       {_GEN_669 & _GEN_671},
       {_GEN_662 & _GEN_664},
       {_GEN_655 & _GEN_657},
       {_GEN_648 & _GEN_650},
       {_GEN_641 & _GEN_643},
       {_GEN_634 & _GEN_636},
       {_GEN_627 & _GEN_629},
       {_GEN_620 & _GEN_622},
       {_GEN_613 & _GEN_615},
       {_GEN_606 & _GEN_608},
       {_GEN_599 & _GEN_601},
       {ldst_forward_matches_0_0}};	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1187:86
    automatic logic        mem_forward_valid_0;	// lsu.scala:1189:53
    automatic logic [5:0]  l_idx;	// Mux.scala:47:69
    automatic logic        ld_xcpt_valid;	// lsu.scala:1238:44
    automatic logic [4:0]  _ld_xcpt_uop_T_3;	// lsu.scala:1239:30
    automatic logic        use_mem_xcpt;	// lsu.scala:1241:115
    automatic logic [15:0] xcpt_uop_br_mask;	// lsu.scala:1243:21
    automatic logic        _ldq_bits_succeeded_T =
      _io_core_exe_0_iresp_valid_output | _io_core_exe_0_fresp_valid_output;	// lsu.scala:1306:5, :1324:72, :1344:5, :1348:5
    automatic logic        _GEN_2059 = _GEN_797 & live;	// AMOALU.scala:10:17, lsu.scala:1369:24, util.scala:118:59
    automatic logic        _GEN_2060;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2061;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2062;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2063;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2064;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2065;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2066;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2067;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2068;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2069;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2070;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2071;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2072;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2073;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2074;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2075;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2076;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2077;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2078;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2079;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2080;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2081;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2082;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2083;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2084;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2085;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2086;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2087;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2088;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2089;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2090;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2091;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2092;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2093;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2094;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2095;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2096;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2097;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2098;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2099;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2100;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2101;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2102;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2103;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2104;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2105;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2106;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_2107;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_2108;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2109;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2110;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2111;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2112;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2113;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2114;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2115;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2116;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2117;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2118;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2119;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2120;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2121;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2122;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2123;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2124;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2125;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2126;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2127;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2128;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2129;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2130;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2131;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_2132;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2133;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2134;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2135;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2136;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2137;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2138;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2139;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2140;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2141;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2142;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2143;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2144;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2145;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2146;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2147;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2148;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2149;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2150;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2151;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2152;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2153;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2154;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2155;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_2156 = idx == 5'h0;	// lsu.scala:1453:18, :1456:31
    automatic logic        _GEN_2157 = commit_store & _GEN_2156;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2158 = idx == 5'h1;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2159 = commit_store & _GEN_2158;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2160 = idx == 5'h2;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2161 = commit_store & _GEN_2160;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2162 = idx == 5'h3;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2163 = commit_store & _GEN_2162;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2164 = idx == 5'h4;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2165 = commit_store & _GEN_2164;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2166 = idx == 5'h5;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2167 = commit_store & _GEN_2166;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2168 = idx == 5'h6;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2169 = commit_store & _GEN_2168;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2170 = idx == 5'h7;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2171 = commit_store & _GEN_2170;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2172 = idx == 5'h8;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2173 = commit_store & _GEN_2172;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2174 = idx == 5'h9;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2175 = commit_store & _GEN_2174;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2176 = idx == 5'hA;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2177 = commit_store & _GEN_2176;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2178 = idx == 5'hB;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2179 = commit_store & _GEN_2178;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2180 = idx == 5'hC;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2181 = commit_store & _GEN_2180;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2182 = idx == 5'hD;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2183 = commit_store & _GEN_2182;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2184 = idx == 5'hE;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2185 = commit_store & _GEN_2184;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2186 = idx == 5'hF;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2187 = commit_store & _GEN_2186;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2188 = idx == 5'h10;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2189 = commit_store & _GEN_2188;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2190 = idx == 5'h11;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2191 = commit_store & _GEN_2190;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2192 = idx == 5'h12;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2193 = commit_store & _GEN_2192;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2194 = idx == 5'h13;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2195 = commit_store & _GEN_2194;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2196 = idx == 5'h14;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2197 = commit_store & _GEN_2196;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2198 = idx == 5'h15;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2199 = commit_store & _GEN_2198;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2200 = idx == 5'h16;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2201 = commit_store & _GEN_2200;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2202 = idx == 5'h17;	// lsu.scala:1453:18, :1456:31, util.scala:205:25
    automatic logic        _GEN_2203 = commit_store & _GEN_2202;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_2204;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2205 = commit_store | ~commit_load;	// lsu.scala:1424:5, :1451:49, :1452:49, :1455:5, :1457:31
    automatic logic        _GEN_2206;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2207;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2208;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2209;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2210;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2211;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2212;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2213;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2214;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2215;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2216;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2217;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2218;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2219;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2220;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2221;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2222;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2223;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2224;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2225;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2226;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2227;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2228;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_2229 = commit_store | ~(commit_load & _GEN_2156);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2230 = commit_store | ~(commit_load & _GEN_2158);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2231 = commit_store | ~(commit_load & _GEN_2160);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2232 = commit_store | ~(commit_load & _GEN_2162);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2233 = commit_store | ~(commit_load & _GEN_2164);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2234 = commit_store | ~(commit_load & _GEN_2166);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2235 = commit_store | ~(commit_load & _GEN_2168);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2236 = commit_store | ~(commit_load & _GEN_2170);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2237 = commit_store | ~(commit_load & _GEN_2172);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2238 = commit_store | ~(commit_load & _GEN_2174);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2239 = commit_store | ~(commit_load & _GEN_2176);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2240 = commit_store | ~(commit_load & _GEN_2178);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2241 = commit_store | ~(commit_load & _GEN_2180);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2242 = commit_store | ~(commit_load & _GEN_2182);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2243 = commit_store | ~(commit_load & _GEN_2184);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2244 = commit_store | ~(commit_load & _GEN_2186);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2245 = commit_store | ~(commit_load & _GEN_2188);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2246 = commit_store | ~(commit_load & _GEN_2190);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2247 = commit_store | ~(commit_load & _GEN_2192);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2248 = commit_store | ~(commit_load & _GEN_2194);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2249 = commit_store | ~(commit_load & _GEN_2196);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2250 = commit_store | ~(commit_load & _GEN_2198);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2251 = commit_store | ~(commit_load & _GEN_2200);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2252 = commit_store | ~(commit_load & _GEN_2202);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_2253 = idx_1 == 5'h0;	// lsu.scala:1453:18, :1456:31
    automatic logic        _GEN_2254 = idx_1 == 5'h1;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2255 = idx_1 == 5'h2;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2256 = idx_1 == 5'h3;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2257 = idx_1 == 5'h4;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2258 = idx_1 == 5'h5;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2259 = idx_1 == 5'h6;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2260 = idx_1 == 5'h7;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2261 = idx_1 == 5'h8;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2262 = idx_1 == 5'h9;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2263 = idx_1 == 5'hA;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2264 = idx_1 == 5'hB;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2265 = idx_1 == 5'hC;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2266 = idx_1 == 5'hD;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2267 = idx_1 == 5'hE;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2268 = idx_1 == 5'hF;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2269 = idx_1 == 5'h10;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2270 = idx_1 == 5'h11;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2271 = idx_1 == 5'h12;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2272 = idx_1 == 5'h13;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2273 = idx_1 == 5'h14;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2274 = idx_1 == 5'h15;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2275 = idx_1 == 5'h16;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2276 = idx_1 == 5'h17;	// lsu.scala:1453:18, :1456:31, util.scala:205:25
    automatic logic        _GEN_2277 = commit_store_1 | ~(commit_load_1 & _GEN_2253);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2278 = commit_store_1 | ~(commit_load_1 & _GEN_2254);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2279 = commit_store_1 | ~(commit_load_1 & _GEN_2255);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2280 = commit_store_1 | ~(commit_load_1 & _GEN_2256);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2281 = commit_store_1 | ~(commit_load_1 & _GEN_2257);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2282 = commit_store_1 | ~(commit_load_1 & _GEN_2258);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2283 = commit_store_1 | ~(commit_load_1 & _GEN_2259);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2284 = commit_store_1 | ~(commit_load_1 & _GEN_2260);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2285 = commit_store_1 | ~(commit_load_1 & _GEN_2261);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2286 = commit_store_1 | ~(commit_load_1 & _GEN_2262);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2287 = commit_store_1 | ~(commit_load_1 & _GEN_2263);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2288 = commit_store_1 | ~(commit_load_1 & _GEN_2264);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2289 = commit_store_1 | ~(commit_load_1 & _GEN_2265);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2290 = commit_store_1 | ~(commit_load_1 & _GEN_2266);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2291 = commit_store_1 | ~(commit_load_1 & _GEN_2267);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2292 = commit_store_1 | ~(commit_load_1 & _GEN_2268);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2293 = commit_store_1 | ~(commit_load_1 & _GEN_2269);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2294 = commit_store_1 | ~(commit_load_1 & _GEN_2270);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2295 = commit_store_1 | ~(commit_load_1 & _GEN_2271);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2296 = commit_store_1 | ~(commit_load_1 & _GEN_2272);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2297 = commit_store_1 | ~(commit_load_1 & _GEN_2273);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2298 = commit_store_1 | ~(commit_load_1 & _GEN_2274);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2299 = commit_store_1 | ~(commit_load_1 & _GEN_2275);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2300 = commit_store_1 | ~(commit_load_1 & _GEN_2276);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2301 = idx_2 == 5'h0;	// lsu.scala:1453:18, :1456:31
    automatic logic        _GEN_2302 = idx_2 == 5'h1;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2303 = idx_2 == 5'h2;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2304 = idx_2 == 5'h3;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2305 = idx_2 == 5'h4;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2306 = idx_2 == 5'h5;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2307 = idx_2 == 5'h6;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2308 = idx_2 == 5'h7;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2309 = idx_2 == 5'h8;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2310 = idx_2 == 5'h9;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2311 = idx_2 == 5'hA;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2312 = idx_2 == 5'hB;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2313 = idx_2 == 5'hC;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2314 = idx_2 == 5'hD;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2315 = idx_2 == 5'hE;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2316 = idx_2 == 5'hF;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2317 = idx_2 == 5'h10;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2318 = idx_2 == 5'h11;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2319 = idx_2 == 5'h12;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2320 = idx_2 == 5'h13;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2321 = idx_2 == 5'h14;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2322 = idx_2 == 5'h15;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2323 = idx_2 == 5'h16;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_2324 = idx_2 == 5'h17;	// lsu.scala:1453:18, :1456:31, util.scala:205:25
    automatic logic        _GEN_2325 = commit_store_2 | ~(commit_load_2 & _GEN_2301);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2326 = commit_store_2 | ~(commit_load_2 & _GEN_2302);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2327 = commit_store_2 | ~(commit_load_2 & _GEN_2303);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2328 = commit_store_2 | ~(commit_load_2 & _GEN_2304);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2329 = commit_store_2 | ~(commit_load_2 & _GEN_2305);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2330 = commit_store_2 | ~(commit_load_2 & _GEN_2306);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2331 = commit_store_2 | ~(commit_load_2 & _GEN_2307);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2332 = commit_store_2 | ~(commit_load_2 & _GEN_2308);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2333 = commit_store_2 | ~(commit_load_2 & _GEN_2309);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2334 = commit_store_2 | ~(commit_load_2 & _GEN_2310);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2335 = commit_store_2 | ~(commit_load_2 & _GEN_2311);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2336 = commit_store_2 | ~(commit_load_2 & _GEN_2312);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2337 = commit_store_2 | ~(commit_load_2 & _GEN_2313);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2338 = commit_store_2 | ~(commit_load_2 & _GEN_2314);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2339 = commit_store_2 | ~(commit_load_2 & _GEN_2315);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2340 = commit_store_2 | ~(commit_load_2 & _GEN_2316);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2341 = commit_store_2 | ~(commit_load_2 & _GEN_2317);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2342 = commit_store_2 | ~(commit_load_2 & _GEN_2318);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2343 = commit_store_2 | ~(commit_load_2 & _GEN_2319);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2344 = commit_store_2 | ~(commit_load_2 & _GEN_2320);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2345 = commit_store_2 | ~(commit_load_2 & _GEN_2321);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2346 = commit_store_2 | ~(commit_load_2 & _GEN_2322);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2347 = commit_store_2 | ~(commit_load_2 & _GEN_2323);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2348 = commit_store_2 | ~(commit_load_2 & _GEN_2324);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_2349;	// lsu.scala:1506:35
    automatic logic        _GEN_2350;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2351;	// lsu.scala:1506:35
    automatic logic        _GEN_2352;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2353;	// lsu.scala:1506:35
    automatic logic        _GEN_2354;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2355;	// lsu.scala:1506:35
    automatic logic        _GEN_2356;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2357;	// lsu.scala:1506:35
    automatic logic        _GEN_2358;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2359;	// lsu.scala:1506:35
    automatic logic        _GEN_2360;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2361;	// lsu.scala:1506:35
    automatic logic        _GEN_2362;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2363;	// lsu.scala:1506:35
    automatic logic        _GEN_2364;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2365;	// lsu.scala:1506:35
    automatic logic        _GEN_2366;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2367;	// lsu.scala:1506:35
    automatic logic        _GEN_2368;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2369;	// lsu.scala:1506:35
    automatic logic        _GEN_2370;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2371;	// lsu.scala:1506:35
    automatic logic        _GEN_2372;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2373;	// lsu.scala:1506:35
    automatic logic        _GEN_2374;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2375;	// lsu.scala:1506:35
    automatic logic        _GEN_2376;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2377;	// lsu.scala:1506:35
    automatic logic        _GEN_2378;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2379;	// lsu.scala:1506:35
    automatic logic        _GEN_2380;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2381;	// lsu.scala:1506:35
    automatic logic        _GEN_2382;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2383;	// lsu.scala:1506:35
    automatic logic        _GEN_2384;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2385;	// lsu.scala:1506:35
    automatic logic        _GEN_2386;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2387;	// lsu.scala:1506:35
    automatic logic        _GEN_2388;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2389;	// lsu.scala:1506:35
    automatic logic        _GEN_2390;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2391;	// lsu.scala:1506:35
    automatic logic        _GEN_2392;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2393;	// lsu.scala:1506:35
    automatic logic        _GEN_2394;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2395;	// lsu.scala:1506:35
    automatic logic        _GEN_2396;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_2397;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2398;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2399;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2400;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2401;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2402;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2403;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2404;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2405;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2406;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2407;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2408;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2409;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2410;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2411;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2412;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2413;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2414;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2415;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2416;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2417;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2418;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2419;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2420;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_2421;	// Decoupled.scala:40:37
    automatic logic        _GEN_2422;	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
    automatic logic        _GEN_2423;	// lsu.scala:244:34, :1527:34, :1533:38
    automatic logic        _GEN_2424;	// lsu.scala:1596:22
    automatic logic        _GEN_2425;	// lsu.scala:1505:3, :1597:3, :1602:5, :1603:16
    automatic logic        _GEN_2426;	// lsu.scala:1622:38
    automatic logic        _GEN_2427;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2428;	// lsu.scala:1622:38
    automatic logic        _GEN_2429;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2430;	// lsu.scala:1622:38
    automatic logic        _GEN_2431;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2432;	// lsu.scala:1622:38
    automatic logic        _GEN_2433;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2434;	// lsu.scala:1622:38
    automatic logic        _GEN_2435;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2436;	// lsu.scala:1622:38
    automatic logic        _GEN_2437;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2438;	// lsu.scala:1622:38
    automatic logic        _GEN_2439;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2440;	// lsu.scala:1622:38
    automatic logic        _GEN_2441;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2442;	// lsu.scala:1622:38
    automatic logic        _GEN_2443;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2444;	// lsu.scala:1622:38
    automatic logic        _GEN_2445;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2446;	// lsu.scala:1622:38
    automatic logic        _GEN_2447;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2448;	// lsu.scala:1622:38
    automatic logic        _GEN_2449;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2450;	// lsu.scala:1622:38
    automatic logic        _GEN_2451;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2452;	// lsu.scala:1622:38
    automatic logic        _GEN_2453;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2454;	// lsu.scala:1622:38
    automatic logic        _GEN_2455;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2456;	// lsu.scala:1622:38
    automatic logic        _GEN_2457;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2458;	// lsu.scala:1622:38
    automatic logic        _GEN_2459;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2460;	// lsu.scala:1622:38
    automatic logic        _GEN_2461;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2462;	// lsu.scala:1622:38
    automatic logic        _GEN_2463;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2464;	// lsu.scala:1622:38
    automatic logic        _GEN_2465;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2466;	// lsu.scala:1622:38
    automatic logic        _GEN_2467;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2468;	// lsu.scala:1622:38
    automatic logic        _GEN_2469;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2470;	// lsu.scala:1622:38
    automatic logic        _GEN_2471;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_2472;	// lsu.scala:1622:38
    automatic logic        _GEN_2473;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic [5:0]  _ldq_retry_idx_idx_T_34;	// Mux.scala:47:69
    automatic logic [5:0]  _stq_retry_idx_idx_T_34;	// Mux.scala:47:69
    automatic logic [5:0]  _ldq_wakeup_idx_idx_T_34;	// Mux.scala:47:69
    _ldq_23_bits_st_dep_mask_T = 32'h1 << stq_head;	// lsu.scala:217:29, :260:71
    _GEN_853 = {24{~clear_store}};	// lsu.scala:260:33, :1495:3, :1500:17
    _GEN_854 = (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & live_store_mask;	// lsu.scala:259:32, :260:{33,65,71}
    _GEN_855 = dis_ld_val & ldq_tail == 5'h0;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_856 = dis_ld_val & ldq_tail == 5'h1;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_857 = dis_ld_val & ldq_tail == 5'h2;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_858 = dis_ld_val & ldq_tail == 5'h3;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_859 = dis_ld_val & ldq_tail == 5'h4;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_860 = dis_ld_val & ldq_tail == 5'h5;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_861 = dis_ld_val & ldq_tail == 5'h6;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_862 = dis_ld_val & ldq_tail == 5'h7;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_863 = dis_ld_val & ldq_tail == 5'h8;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_864 = dis_ld_val & ldq_tail == 5'h9;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_865 = dis_ld_val & ldq_tail == 5'hA;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_866 = dis_ld_val & ldq_tail == 5'hB;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_867 = dis_ld_val & ldq_tail == 5'hC;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_868 = dis_ld_val & ldq_tail == 5'hD;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_869 = dis_ld_val & ldq_tail == 5'hE;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_870 = dis_ld_val & ldq_tail == 5'hF;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_871 = dis_ld_val & ldq_tail == 5'h10;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_872 = dis_ld_val & ldq_tail == 5'h11;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_873 = dis_ld_val & ldq_tail == 5'h12;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_874 = dis_ld_val & ldq_tail == 5'h13;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_875 = dis_ld_val & ldq_tail == 5'h14;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_876 = dis_ld_val & ldq_tail == 5'h15;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_877 = dis_ld_val & ldq_tail == 5'h16;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_878 = dis_ld_val & ldq_tail == 5'h17;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44, util.scala:205:25
    _GEN_879 = dis_st_val & stq_tail == 5'h0;	// lsu.scala:211:16, :218:29, :302:85, :321:5, :322:39
    _GEN_880 = dis_st_val & stq_tail == 5'h1;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_881 = dis_st_val & stq_tail == 5'h2;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_882 = dis_st_val & stq_tail == 5'h3;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_883 = dis_st_val & stq_tail == 5'h4;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_884 = dis_st_val & stq_tail == 5'h5;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_885 = dis_st_val & stq_tail == 5'h6;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_886 = dis_st_val & stq_tail == 5'h7;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_887 = dis_st_val & stq_tail == 5'h8;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_888 = dis_st_val & stq_tail == 5'h9;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_889 = dis_st_val & stq_tail == 5'hA;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_890 = dis_st_val & stq_tail == 5'hB;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_891 = dis_st_val & stq_tail == 5'hC;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_892 = dis_st_val & stq_tail == 5'hD;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_893 = dis_st_val & stq_tail == 5'hE;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_894 = dis_st_val & stq_tail == 5'hF;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_895 = dis_st_val & stq_tail == 5'h10;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_896 = dis_st_val & stq_tail == 5'h11;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_897 = dis_st_val & stq_tail == 5'h12;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_898 = dis_st_val & stq_tail == 5'h13;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_899 = dis_st_val & stq_tail == 5'h14;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_900 = dis_st_val & stq_tail == 5'h15;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_901 = dis_st_val & stq_tail == 5'h16;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_902 = dis_st_val & stq_tail == 5'h17;	// lsu.scala:211:16, :218:29, :302:85, :321:5, :322:39, util.scala:205:25
    _GEN_903 = dis_ld_val | ~_GEN_879;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_904 = dis_ld_val | ~_GEN_880;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_905 = dis_ld_val | ~_GEN_881;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_906 = dis_ld_val | ~_GEN_882;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_907 = dis_ld_val | ~_GEN_883;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_908 = dis_ld_val | ~_GEN_884;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_909 = dis_ld_val | ~_GEN_885;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_910 = dis_ld_val | ~_GEN_886;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_911 = dis_ld_val | ~_GEN_887;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_912 = dis_ld_val | ~_GEN_888;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_913 = dis_ld_val | ~_GEN_889;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_914 = dis_ld_val | ~_GEN_890;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_915 = dis_ld_val | ~_GEN_891;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_916 = dis_ld_val | ~_GEN_892;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_917 = dis_ld_val | ~_GEN_893;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_918 = dis_ld_val | ~_GEN_894;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_919 = dis_ld_val | ~_GEN_895;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_920 = dis_ld_val | ~_GEN_896;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_921 = dis_ld_val | ~_GEN_897;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_922 = dis_ld_val | ~_GEN_898;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_923 = dis_ld_val | ~_GEN_899;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_924 = dis_ld_val | ~_GEN_900;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_925 = dis_ld_val | ~_GEN_901;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_926 = dis_ld_val | ~_GEN_902;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_927 = 32'h1 << stq_tail;	// lsu.scala:218:29, :260:71, :336:72
    _GEN_928 = {24{dis_st_val}} & _GEN_927[23:0] | _GEN_854;	// lsu.scala:260:33, :302:85, :336:{31,72}
    _GEN_930 = _GEN_929 | _GEN_855;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_932 = _GEN_931 | _GEN_856;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_934 = _GEN_933 | _GEN_857;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_936 = _GEN_935 | _GEN_858;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_938 = _GEN_937 | _GEN_859;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_940 = _GEN_939 | _GEN_860;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_942 = _GEN_941 | _GEN_861;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_944 = _GEN_943 | _GEN_862;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_946 = _GEN_945 | _GEN_863;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_948 = _GEN_947 | _GEN_864;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_950 = _GEN_949 | _GEN_865;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_952 = _GEN_951 | _GEN_866;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_954 = _GEN_953 | _GEN_867;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_956 = _GEN_955 | _GEN_868;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_958 = _GEN_957 | _GEN_869;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_960 = _GEN_959 | _GEN_870;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_962 = _GEN_961 | _GEN_871;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_964 = _GEN_963 | _GEN_872;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_966 = _GEN_965 | _GEN_873;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_968 = _GEN_967 | _GEN_874;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_970 = _GEN_969 | _GEN_875;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_972 = _GEN_971 | _GEN_876;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_974 = _GEN_973 | _GEN_877;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_976 = _GEN_975 | _GEN_878;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_977 = dis_ld_val_1 & _GEN_929;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_978 = dis_ld_val_1 & _GEN_931;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_979 = dis_ld_val_1 & _GEN_933;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_980 = dis_ld_val_1 & _GEN_935;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_981 = dis_ld_val_1 & _GEN_937;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_982 = dis_ld_val_1 & _GEN_939;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_983 = dis_ld_val_1 & _GEN_941;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_984 = dis_ld_val_1 & _GEN_943;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_985 = dis_ld_val_1 & _GEN_945;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_986 = dis_ld_val_1 & _GEN_947;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_987 = dis_ld_val_1 & _GEN_949;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_988 = dis_ld_val_1 & _GEN_951;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_989 = dis_ld_val_1 & _GEN_953;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_990 = dis_ld_val_1 & _GEN_955;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_991 = dis_ld_val_1 & _GEN_957;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_992 = dis_ld_val_1 & _GEN_959;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_993 = dis_ld_val_1 & _GEN_961;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_994 = dis_ld_val_1 & _GEN_963;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_995 = dis_ld_val_1 & _GEN_965;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_996 = dis_ld_val_1 & _GEN_967;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_997 = dis_ld_val_1 & _GEN_969;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_998 = dis_ld_val_1 & _GEN_971;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_999 = dis_ld_val_1 & _GEN_973;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_1000 = dis_ld_val_1 & _GEN_975;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_1001 = dis_st_val_1 & _GEN_101 == 5'h0;	// lsu.scala:302:85, :304:5, :321:5, :322:39, :338:21
    _GEN_1002 = dis_st_val_1 & _GEN_101 == 5'h1;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1003 = dis_st_val_1 & _GEN_101 == 5'h2;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1004 = dis_st_val_1 & _GEN_101 == 5'h3;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1005 = dis_st_val_1 & _GEN_101 == 5'h4;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1006 = dis_st_val_1 & _GEN_101 == 5'h5;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1007 = dis_st_val_1 & _GEN_101 == 5'h6;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1008 = dis_st_val_1 & _GEN_101 == 5'h7;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1009 = dis_st_val_1 & _GEN_101 == 5'h8;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1010 = dis_st_val_1 & _GEN_101 == 5'h9;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1011 = dis_st_val_1 & _GEN_101 == 5'hA;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1012 = dis_st_val_1 & _GEN_101 == 5'hB;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1013 = dis_st_val_1 & _GEN_101 == 5'hC;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1014 = dis_st_val_1 & _GEN_101 == 5'hD;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1015 = dis_st_val_1 & _GEN_101 == 5'hE;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1016 = dis_st_val_1 & _GEN_101 == 5'hF;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1017 = dis_st_val_1 & _GEN_101 == 5'h10;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1018 = dis_st_val_1 & _GEN_101 == 5'h11;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1019 = dis_st_val_1 & _GEN_101 == 5'h12;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1020 = dis_st_val_1 & _GEN_101 == 5'h13;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1021 = dis_st_val_1 & _GEN_101 == 5'h14;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1022 = dis_st_val_1 & _GEN_101 == 5'h15;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1023 = dis_st_val_1 & _GEN_101 == 5'h16;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_1024 = dis_st_val_1 & _GEN_101 == 5'h17;	// lsu.scala:302:85, :304:5, :321:5, :322:39, :338:21, util.scala:205:25
    _GEN_1025 = dis_ld_val_1 | ~_GEN_1001;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1026 = dis_ld_val_1 | ~_GEN_1002;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1027 = dis_ld_val_1 | ~_GEN_1003;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1028 = dis_ld_val_1 | ~_GEN_1004;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1029 = dis_ld_val_1 | ~_GEN_1005;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1030 = dis_ld_val_1 | ~_GEN_1006;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1031 = dis_ld_val_1 | ~_GEN_1007;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1032 = dis_ld_val_1 | ~_GEN_1008;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1033 = dis_ld_val_1 | ~_GEN_1009;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1034 = dis_ld_val_1 | ~_GEN_1010;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1035 = dis_ld_val_1 | ~_GEN_1011;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1036 = dis_ld_val_1 | ~_GEN_1012;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1037 = dis_ld_val_1 | ~_GEN_1013;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1038 = dis_ld_val_1 | ~_GEN_1014;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1039 = dis_ld_val_1 | ~_GEN_1015;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1040 = dis_ld_val_1 | ~_GEN_1016;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1041 = dis_ld_val_1 | ~_GEN_1017;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1042 = dis_ld_val_1 | ~_GEN_1018;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1043 = dis_ld_val_1 | ~_GEN_1019;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1044 = dis_ld_val_1 | ~_GEN_1020;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1045 = dis_ld_val_1 | ~_GEN_1021;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1046 = dis_ld_val_1 | ~_GEN_1022;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1047 = dis_ld_val_1 | ~_GEN_1023;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1048 = dis_ld_val_1 | ~_GEN_1024;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1050 = {24{dis_st_val_1}} & _GEN_1049[23:0] | _GEN_928;	// lsu.scala:302:85, :336:{31,72}
    _GEN_1051 = dis_ld_val_2 & _GEN_106 == 5'h0;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1052 =
      _GEN_1051 | (dis_ld_val_1 ? _GEN_930 | ldq_0_valid : _GEN_855 | ldq_0_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1053 = dis_ld_val_2 & _GEN_106 == 5'h1;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1054 =
      _GEN_1053 | (dis_ld_val_1 ? _GEN_932 | ldq_1_valid : _GEN_856 | ldq_1_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1055 = dis_ld_val_2 & _GEN_106 == 5'h2;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1056 =
      _GEN_1055 | (dis_ld_val_1 ? _GEN_934 | ldq_2_valid : _GEN_857 | ldq_2_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1057 = dis_ld_val_2 & _GEN_106 == 5'h3;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1058 =
      _GEN_1057 | (dis_ld_val_1 ? _GEN_936 | ldq_3_valid : _GEN_858 | ldq_3_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1059 = dis_ld_val_2 & _GEN_106 == 5'h4;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1060 =
      _GEN_1059 | (dis_ld_val_1 ? _GEN_938 | ldq_4_valid : _GEN_859 | ldq_4_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1061 = dis_ld_val_2 & _GEN_106 == 5'h5;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1062 =
      _GEN_1061 | (dis_ld_val_1 ? _GEN_940 | ldq_5_valid : _GEN_860 | ldq_5_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1063 = dis_ld_val_2 & _GEN_106 == 5'h6;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1064 =
      _GEN_1063 | (dis_ld_val_1 ? _GEN_942 | ldq_6_valid : _GEN_861 | ldq_6_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1065 = dis_ld_val_2 & _GEN_106 == 5'h7;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1066 =
      _GEN_1065 | (dis_ld_val_1 ? _GEN_944 | ldq_7_valid : _GEN_862 | ldq_7_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1067 = dis_ld_val_2 & _GEN_106 == 5'h8;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1068 =
      _GEN_1067 | (dis_ld_val_1 ? _GEN_946 | ldq_8_valid : _GEN_863 | ldq_8_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1069 = dis_ld_val_2 & _GEN_106 == 5'h9;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1070 =
      _GEN_1069 | (dis_ld_val_1 ? _GEN_948 | ldq_9_valid : _GEN_864 | ldq_9_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1071 = dis_ld_val_2 & _GEN_106 == 5'hA;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1072 =
      _GEN_1071 | (dis_ld_val_1 ? _GEN_950 | ldq_10_valid : _GEN_865 | ldq_10_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1073 = dis_ld_val_2 & _GEN_106 == 5'hB;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1074 =
      _GEN_1073 | (dis_ld_val_1 ? _GEN_952 | ldq_11_valid : _GEN_866 | ldq_11_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1075 = dis_ld_val_2 & _GEN_106 == 5'hC;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1076 =
      _GEN_1075 | (dis_ld_val_1 ? _GEN_954 | ldq_12_valid : _GEN_867 | ldq_12_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1077 = dis_ld_val_2 & _GEN_106 == 5'hD;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1078 =
      _GEN_1077 | (dis_ld_val_1 ? _GEN_956 | ldq_13_valid : _GEN_868 | ldq_13_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1079 = dis_ld_val_2 & _GEN_106 == 5'hE;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1080 =
      _GEN_1079 | (dis_ld_val_1 ? _GEN_958 | ldq_14_valid : _GEN_869 | ldq_14_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1081 = dis_ld_val_2 & _GEN_106 == 5'hF;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1082 =
      _GEN_1081 | (dis_ld_val_1 ? _GEN_960 | ldq_15_valid : _GEN_870 | ldq_15_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1083 = dis_ld_val_2 & _GEN_106 == 5'h10;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1084 =
      _GEN_1083 | (dis_ld_val_1 ? _GEN_962 | ldq_16_valid : _GEN_871 | ldq_16_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1085 = dis_ld_val_2 & _GEN_106 == 5'h11;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1086 =
      _GEN_1085 | (dis_ld_val_1 ? _GEN_964 | ldq_17_valid : _GEN_872 | ldq_17_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1087 = dis_ld_val_2 & _GEN_106 == 5'h12;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1088 =
      _GEN_1087 | (dis_ld_val_1 ? _GEN_966 | ldq_18_valid : _GEN_873 | ldq_18_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1089 = dis_ld_val_2 & _GEN_106 == 5'h13;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1090 =
      _GEN_1089 | (dis_ld_val_1 ? _GEN_968 | ldq_19_valid : _GEN_874 | ldq_19_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1091 = dis_ld_val_2 & _GEN_106 == 5'h14;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1092 =
      _GEN_1091 | (dis_ld_val_1 ? _GEN_970 | ldq_20_valid : _GEN_875 | ldq_20_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1093 = dis_ld_val_2 & _GEN_106 == 5'h15;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1094 =
      _GEN_1093 | (dis_ld_val_1 ? _GEN_972 | ldq_21_valid : _GEN_876 | ldq_21_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1095 = dis_ld_val_2 & _GEN_106 == 5'h16;	// lsu.scala:301:85, :304:5, :305:44, :333:21
    _GEN_1096 =
      _GEN_1095 | (dis_ld_val_1 ? _GEN_974 | ldq_22_valid : _GEN_877 | ldq_22_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1097 = dis_ld_val_2 & _GEN_106 == 5'h17;	// lsu.scala:301:85, :304:5, :305:44, :333:21, util.scala:205:25
    _GEN_1098 =
      _GEN_1097 | (dis_ld_val_1 ? _GEN_976 | ldq_23_valid : _GEN_878 | ldq_23_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_1099 = _GEN_1051 | _GEN_977 | _GEN_855;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1100 = _GEN_1053 | _GEN_978 | _GEN_856;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1101 = _GEN_1055 | _GEN_979 | _GEN_857;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1102 = _GEN_1057 | _GEN_980 | _GEN_858;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1103 = _GEN_1059 | _GEN_981 | _GEN_859;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1104 = _GEN_1061 | _GEN_982 | _GEN_860;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1105 = _GEN_1063 | _GEN_983 | _GEN_861;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1106 = _GEN_1065 | _GEN_984 | _GEN_862;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1107 = _GEN_1067 | _GEN_985 | _GEN_863;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1108 = _GEN_1069 | _GEN_986 | _GEN_864;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1109 = _GEN_1071 | _GEN_987 | _GEN_865;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1110 = _GEN_1073 | _GEN_988 | _GEN_866;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1111 = _GEN_1075 | _GEN_989 | _GEN_867;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1112 = _GEN_1077 | _GEN_990 | _GEN_868;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1113 = _GEN_1079 | _GEN_991 | _GEN_869;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1114 = _GEN_1081 | _GEN_992 | _GEN_870;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1115 = _GEN_1083 | _GEN_993 | _GEN_871;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1116 = _GEN_1085 | _GEN_994 | _GEN_872;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1117 = _GEN_1087 | _GEN_995 | _GEN_873;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1118 = _GEN_1089 | _GEN_996 | _GEN_874;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1119 = _GEN_1091 | _GEN_997 | _GEN_875;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1120 = _GEN_1093 | _GEN_998 | _GEN_876;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1121 = _GEN_1095 | _GEN_999 | _GEN_877;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1122 = _GEN_1097 | _GEN_1000 | _GEN_878;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_1123 =
      ~_GEN_1051
      & (dis_ld_val_1
           ? ~_GEN_930 & ldq_0_bits_order_fail
           : ~_GEN_855 & ldq_0_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1124 =
      ~_GEN_1053
      & (dis_ld_val_1
           ? ~_GEN_932 & ldq_1_bits_order_fail
           : ~_GEN_856 & ldq_1_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1125 =
      ~_GEN_1055
      & (dis_ld_val_1
           ? ~_GEN_934 & ldq_2_bits_order_fail
           : ~_GEN_857 & ldq_2_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1126 =
      ~_GEN_1057
      & (dis_ld_val_1
           ? ~_GEN_936 & ldq_3_bits_order_fail
           : ~_GEN_858 & ldq_3_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1127 =
      ~_GEN_1059
      & (dis_ld_val_1
           ? ~_GEN_938 & ldq_4_bits_order_fail
           : ~_GEN_859 & ldq_4_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1128 =
      ~_GEN_1061
      & (dis_ld_val_1
           ? ~_GEN_940 & ldq_5_bits_order_fail
           : ~_GEN_860 & ldq_5_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1129 =
      ~_GEN_1063
      & (dis_ld_val_1
           ? ~_GEN_942 & ldq_6_bits_order_fail
           : ~_GEN_861 & ldq_6_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1130 =
      ~_GEN_1065
      & (dis_ld_val_1
           ? ~_GEN_944 & ldq_7_bits_order_fail
           : ~_GEN_862 & ldq_7_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1131 =
      ~_GEN_1067
      & (dis_ld_val_1
           ? ~_GEN_946 & ldq_8_bits_order_fail
           : ~_GEN_863 & ldq_8_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1132 =
      ~_GEN_1069
      & (dis_ld_val_1
           ? ~_GEN_948 & ldq_9_bits_order_fail
           : ~_GEN_864 & ldq_9_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1133 =
      ~_GEN_1071
      & (dis_ld_val_1
           ? ~_GEN_950 & ldq_10_bits_order_fail
           : ~_GEN_865 & ldq_10_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1134 =
      ~_GEN_1073
      & (dis_ld_val_1
           ? ~_GEN_952 & ldq_11_bits_order_fail
           : ~_GEN_866 & ldq_11_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1135 =
      ~_GEN_1075
      & (dis_ld_val_1
           ? ~_GEN_954 & ldq_12_bits_order_fail
           : ~_GEN_867 & ldq_12_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1136 =
      ~_GEN_1077
      & (dis_ld_val_1
           ? ~_GEN_956 & ldq_13_bits_order_fail
           : ~_GEN_868 & ldq_13_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1137 =
      ~_GEN_1079
      & (dis_ld_val_1
           ? ~_GEN_958 & ldq_14_bits_order_fail
           : ~_GEN_869 & ldq_14_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1138 =
      ~_GEN_1081
      & (dis_ld_val_1
           ? ~_GEN_960 & ldq_15_bits_order_fail
           : ~_GEN_870 & ldq_15_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1139 =
      ~_GEN_1083
      & (dis_ld_val_1
           ? ~_GEN_962 & ldq_16_bits_order_fail
           : ~_GEN_871 & ldq_16_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1140 =
      ~_GEN_1085
      & (dis_ld_val_1
           ? ~_GEN_964 & ldq_17_bits_order_fail
           : ~_GEN_872 & ldq_17_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1141 =
      ~_GEN_1087
      & (dis_ld_val_1
           ? ~_GEN_966 & ldq_18_bits_order_fail
           : ~_GEN_873 & ldq_18_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1142 =
      ~_GEN_1089
      & (dis_ld_val_1
           ? ~_GEN_968 & ldq_19_bits_order_fail
           : ~_GEN_874 & ldq_19_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1143 =
      ~_GEN_1091
      & (dis_ld_val_1
           ? ~_GEN_970 & ldq_20_bits_order_fail
           : ~_GEN_875 & ldq_20_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1144 =
      ~_GEN_1093
      & (dis_ld_val_1
           ? ~_GEN_972 & ldq_21_bits_order_fail
           : ~_GEN_876 & ldq_21_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1145 =
      ~_GEN_1095
      & (dis_ld_val_1
           ? ~_GEN_974 & ldq_22_bits_order_fail
           : ~_GEN_877 & ldq_22_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1146 =
      ~_GEN_1097
      & (dis_ld_val_1
           ? ~_GEN_976 & ldq_23_bits_order_fail
           : ~_GEN_878 & ldq_23_bits_order_fail);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_1148 =
      ~dis_ld_val_2 & _GEN_1147 | ~dis_ld_val_1 & _GEN_1001 | ~dis_ld_val & _GEN_879
      | stq_0_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1150 =
      ~dis_ld_val_2 & _GEN_1149 | ~dis_ld_val_1 & _GEN_1002 | ~dis_ld_val & _GEN_880
      | stq_1_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1152 =
      ~dis_ld_val_2 & _GEN_1151 | ~dis_ld_val_1 & _GEN_1003 | ~dis_ld_val & _GEN_881
      | stq_2_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1154 =
      ~dis_ld_val_2 & _GEN_1153 | ~dis_ld_val_1 & _GEN_1004 | ~dis_ld_val & _GEN_882
      | stq_3_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1156 =
      ~dis_ld_val_2 & _GEN_1155 | ~dis_ld_val_1 & _GEN_1005 | ~dis_ld_val & _GEN_883
      | stq_4_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1158 =
      ~dis_ld_val_2 & _GEN_1157 | ~dis_ld_val_1 & _GEN_1006 | ~dis_ld_val & _GEN_884
      | stq_5_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1160 =
      ~dis_ld_val_2 & _GEN_1159 | ~dis_ld_val_1 & _GEN_1007 | ~dis_ld_val & _GEN_885
      | stq_6_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1162 =
      ~dis_ld_val_2 & _GEN_1161 | ~dis_ld_val_1 & _GEN_1008 | ~dis_ld_val & _GEN_886
      | stq_7_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1164 =
      ~dis_ld_val_2 & _GEN_1163 | ~dis_ld_val_1 & _GEN_1009 | ~dis_ld_val & _GEN_887
      | stq_8_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1166 =
      ~dis_ld_val_2 & _GEN_1165 | ~dis_ld_val_1 & _GEN_1010 | ~dis_ld_val & _GEN_888
      | stq_9_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1168 =
      ~dis_ld_val_2 & _GEN_1167 | ~dis_ld_val_1 & _GEN_1011 | ~dis_ld_val & _GEN_889
      | stq_10_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1170 =
      ~dis_ld_val_2 & _GEN_1169 | ~dis_ld_val_1 & _GEN_1012 | ~dis_ld_val & _GEN_890
      | stq_11_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1172 =
      ~dis_ld_val_2 & _GEN_1171 | ~dis_ld_val_1 & _GEN_1013 | ~dis_ld_val & _GEN_891
      | stq_12_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1174 =
      ~dis_ld_val_2 & _GEN_1173 | ~dis_ld_val_1 & _GEN_1014 | ~dis_ld_val & _GEN_892
      | stq_13_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1176 =
      ~dis_ld_val_2 & _GEN_1175 | ~dis_ld_val_1 & _GEN_1015 | ~dis_ld_val & _GEN_893
      | stq_14_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1178 =
      ~dis_ld_val_2 & _GEN_1177 | ~dis_ld_val_1 & _GEN_1016 | ~dis_ld_val & _GEN_894
      | stq_15_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1180 =
      ~dis_ld_val_2 & _GEN_1179 | ~dis_ld_val_1 & _GEN_1017 | ~dis_ld_val & _GEN_895
      | stq_16_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1182 =
      ~dis_ld_val_2 & _GEN_1181 | ~dis_ld_val_1 & _GEN_1018 | ~dis_ld_val & _GEN_896
      | stq_17_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1184 =
      ~dis_ld_val_2 & _GEN_1183 | ~dis_ld_val_1 & _GEN_1019 | ~dis_ld_val & _GEN_897
      | stq_18_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1186 =
      ~dis_ld_val_2 & _GEN_1185 | ~dis_ld_val_1 & _GEN_1020 | ~dis_ld_val & _GEN_898
      | stq_19_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1188 =
      ~dis_ld_val_2 & _GEN_1187 | ~dis_ld_val_1 & _GEN_1021 | ~dis_ld_val & _GEN_899
      | stq_20_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1190 =
      ~dis_ld_val_2 & _GEN_1189 | ~dis_ld_val_1 & _GEN_1022 | ~dis_ld_val & _GEN_900
      | stq_21_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1192 =
      ~dis_ld_val_2 & _GEN_1191 | ~dis_ld_val_1 & _GEN_1023 | ~dis_ld_val & _GEN_901
      | stq_22_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1194 =
      ~dis_ld_val_2 & _GEN_1193 | ~dis_ld_val_1 & _GEN_1024 | ~dis_ld_val & _GEN_902
      | stq_23_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_1195 = dis_ld_val_2 | ~_GEN_1147;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1196 = dis_ld_val_2 | ~_GEN_1149;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1197 = dis_ld_val_2 | ~_GEN_1151;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1198 = dis_ld_val_2 | ~_GEN_1153;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1199 = dis_ld_val_2 | ~_GEN_1155;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1200 = dis_ld_val_2 | ~_GEN_1157;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1201 = dis_ld_val_2 | ~_GEN_1159;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1202 = dis_ld_val_2 | ~_GEN_1161;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1203 = dis_ld_val_2 | ~_GEN_1163;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1204 = dis_ld_val_2 | ~_GEN_1165;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1205 = dis_ld_val_2 | ~_GEN_1167;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1206 = dis_ld_val_2 | ~_GEN_1169;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1207 = dis_ld_val_2 | ~_GEN_1171;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1208 = dis_ld_val_2 | ~_GEN_1173;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1209 = dis_ld_val_2 | ~_GEN_1175;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1210 = dis_ld_val_2 | ~_GEN_1177;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1211 = dis_ld_val_2 | ~_GEN_1179;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1212 = dis_ld_val_2 | ~_GEN_1181;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1213 = dis_ld_val_2 | ~_GEN_1183;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1214 = dis_ld_val_2 | ~_GEN_1185;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1215 = dis_ld_val_2 | ~_GEN_1187;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1216 = dis_ld_val_2 | ~_GEN_1189;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1217 = dis_ld_val_2 | ~_GEN_1191;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1218 = dis_ld_val_2 | ~_GEN_1193;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_1219 = _GEN_1195 & _GEN_1025 & _GEN_903 & stq_0_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1220 = _GEN_1196 & _GEN_1026 & _GEN_904 & stq_1_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1221 = _GEN_1197 & _GEN_1027 & _GEN_905 & stq_2_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1222 = _GEN_1198 & _GEN_1028 & _GEN_906 & stq_3_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1223 = _GEN_1199 & _GEN_1029 & _GEN_907 & stq_4_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1224 = _GEN_1200 & _GEN_1030 & _GEN_908 & stq_5_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1225 = _GEN_1201 & _GEN_1031 & _GEN_909 & stq_6_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1226 = _GEN_1202 & _GEN_1032 & _GEN_910 & stq_7_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1227 = _GEN_1203 & _GEN_1033 & _GEN_911 & stq_8_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1228 = _GEN_1204 & _GEN_1034 & _GEN_912 & stq_9_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1229 = _GEN_1205 & _GEN_1035 & _GEN_913 & stq_10_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1230 = _GEN_1206 & _GEN_1036 & _GEN_914 & stq_11_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1231 = _GEN_1207 & _GEN_1037 & _GEN_915 & stq_12_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1232 = _GEN_1208 & _GEN_1038 & _GEN_916 & stq_13_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1233 = _GEN_1209 & _GEN_1039 & _GEN_917 & stq_14_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1234 = _GEN_1210 & _GEN_1040 & _GEN_918 & stq_15_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1235 = _GEN_1211 & _GEN_1041 & _GEN_919 & stq_16_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1236 = _GEN_1212 & _GEN_1042 & _GEN_920 & stq_17_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1237 = _GEN_1213 & _GEN_1043 & _GEN_921 & stq_18_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1238 = _GEN_1214 & _GEN_1044 & _GEN_922 & stq_19_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1239 = _GEN_1215 & _GEN_1045 & _GEN_923 & stq_20_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1240 = _GEN_1216 & _GEN_1046 & _GEN_924 & stq_21_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1241 = _GEN_1217 & _GEN_1047 & _GEN_925 & stq_22_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_1242 = _GEN_1218 & _GEN_1048 & _GEN_926 & stq_23_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    ldq_retry_idx_block =
      (will_fire_load_wakeup_0
         ? _GEN_216
         : can_fire_load_incoming_0 ? _GEN_240 : _GEN_265) | p1_block_load_mask_0;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_2 =
      ldq_0_bits_addr_valid & ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_1 =
      (will_fire_load_wakeup_0
         ? _GEN_217
         : can_fire_load_incoming_0 ? _GEN_241 : _GEN_267) | p1_block_load_mask_1;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_5 =
      ldq_1_bits_addr_valid & ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_2 =
      (will_fire_load_wakeup_0
         ? _GEN_218
         : can_fire_load_incoming_0 ? _GEN_242 : _GEN_269) | p1_block_load_mask_2;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_8 =
      ldq_2_bits_addr_valid & ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_3 =
      (will_fire_load_wakeup_0
         ? _GEN_219
         : can_fire_load_incoming_0 ? _GEN_243 : _GEN_271) | p1_block_load_mask_3;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_11 =
      ldq_3_bits_addr_valid & ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_4 =
      (will_fire_load_wakeup_0
         ? _GEN_220
         : can_fire_load_incoming_0 ? _GEN_244 : _GEN_273) | p1_block_load_mask_4;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_14 =
      ldq_4_bits_addr_valid & ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_5 =
      (will_fire_load_wakeup_0
         ? _GEN_221
         : can_fire_load_incoming_0 ? _GEN_245 : _GEN_275) | p1_block_load_mask_5;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_17 =
      ldq_5_bits_addr_valid & ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_6 =
      (will_fire_load_wakeup_0
         ? _GEN_222
         : can_fire_load_incoming_0 ? _GEN_246 : _GEN_277) | p1_block_load_mask_6;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_20 =
      ldq_6_bits_addr_valid & ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_7 =
      (will_fire_load_wakeup_0
         ? _GEN_223
         : can_fire_load_incoming_0 ? _GEN_247 : _GEN_279) | p1_block_load_mask_7;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_23 =
      ldq_7_bits_addr_valid & ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_8 =
      (will_fire_load_wakeup_0
         ? _GEN_224
         : can_fire_load_incoming_0 ? _GEN_248 : _GEN_281) | p1_block_load_mask_8;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_26 =
      ldq_8_bits_addr_valid & ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_9 =
      (will_fire_load_wakeup_0
         ? _GEN_225
         : can_fire_load_incoming_0 ? _GEN_249 : _GEN_283) | p1_block_load_mask_9;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_29 =
      ldq_9_bits_addr_valid & ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_10 =
      (will_fire_load_wakeup_0
         ? _GEN_226
         : can_fire_load_incoming_0 ? _GEN_250 : _GEN_285) | p1_block_load_mask_10;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_32 =
      ldq_10_bits_addr_valid & ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_11 =
      (will_fire_load_wakeup_0
         ? _GEN_227
         : can_fire_load_incoming_0 ? _GEN_251 : _GEN_287) | p1_block_load_mask_11;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_35 =
      ldq_11_bits_addr_valid & ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_12 =
      (will_fire_load_wakeup_0
         ? _GEN_228
         : can_fire_load_incoming_0 ? _GEN_252 : _GEN_289) | p1_block_load_mask_12;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_38 =
      ldq_12_bits_addr_valid & ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_13 =
      (will_fire_load_wakeup_0
         ? _GEN_229
         : can_fire_load_incoming_0 ? _GEN_253 : _GEN_291) | p1_block_load_mask_13;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_41 =
      ldq_13_bits_addr_valid & ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_14 =
      (will_fire_load_wakeup_0
         ? _GEN_230
         : can_fire_load_incoming_0 ? _GEN_254 : _GEN_293) | p1_block_load_mask_14;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_44 =
      ldq_14_bits_addr_valid & ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_15 =
      (will_fire_load_wakeup_0
         ? _GEN_231
         : can_fire_load_incoming_0 ? _GEN_255 : _GEN_295) | p1_block_load_mask_15;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_47 =
      ldq_15_bits_addr_valid & ldq_15_bits_addr_is_virtual & ~ldq_retry_idx_block_15;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_16 =
      (will_fire_load_wakeup_0
         ? _GEN_232
         : can_fire_load_incoming_0 ? _GEN_256 : _GEN_297) | p1_block_load_mask_16;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_50 =
      ldq_16_bits_addr_valid & ldq_16_bits_addr_is_virtual & ~ldq_retry_idx_block_16;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_17 =
      (will_fire_load_wakeup_0
         ? _GEN_233
         : can_fire_load_incoming_0 ? _GEN_257 : _GEN_299) | p1_block_load_mask_17;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_53 =
      ldq_17_bits_addr_valid & ldq_17_bits_addr_is_virtual & ~ldq_retry_idx_block_17;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_18 =
      (will_fire_load_wakeup_0
         ? _GEN_234
         : can_fire_load_incoming_0 ? _GEN_258 : _GEN_301) | p1_block_load_mask_18;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_56 =
      ldq_18_bits_addr_valid & ldq_18_bits_addr_is_virtual & ~ldq_retry_idx_block_18;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_19 =
      (will_fire_load_wakeup_0
         ? _GEN_235
         : can_fire_load_incoming_0 ? _GEN_259 : _GEN_303) | p1_block_load_mask_19;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_59 =
      ldq_19_bits_addr_valid & ldq_19_bits_addr_is_virtual & ~ldq_retry_idx_block_19;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_20 =
      (will_fire_load_wakeup_0
         ? _GEN_236
         : can_fire_load_incoming_0 ? _GEN_260 : _GEN_305) | p1_block_load_mask_20;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_62 =
      ldq_20_bits_addr_valid & ldq_20_bits_addr_is_virtual & ~ldq_retry_idx_block_20;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_21 =
      (will_fire_load_wakeup_0
         ? _GEN_237
         : can_fire_load_incoming_0 ? _GEN_261 : _GEN_307) | p1_block_load_mask_21;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_65 =
      ldq_21_bits_addr_valid & ldq_21_bits_addr_is_virtual & ~ldq_retry_idx_block_21;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_22 =
      (will_fire_load_wakeup_0
         ? _GEN_238
         : can_fire_load_incoming_0 ? _GEN_262 : _GEN_309) | p1_block_load_mask_22;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_68 =
      ldq_22_bits_addr_valid & ldq_22_bits_addr_is_virtual & ~ldq_retry_idx_block_22;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_23 =
      (will_fire_load_wakeup_0
         ? _GEN_239
         : can_fire_load_incoming_0 ? _GEN_263 : _GEN_311) | p1_block_load_mask_23;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _temp_bits_T = ldq_head == 5'h0;	// lsu.scala:215:29, util.scala:351:72
    _temp_bits_T_2 = ldq_head < 5'h2;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_4 = ldq_head < 5'h3;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_6 = ldq_head < 5'h4;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_8 = ldq_head < 5'h5;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_10 = ldq_head < 5'h6;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_12 = ldq_head < 5'h7;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_14 = ldq_head < 5'h8;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_16 = ldq_head < 5'h9;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_18 = ldq_head < 5'hA;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_20 = ldq_head < 5'hB;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_22 = ldq_head < 5'hC;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_24 = ldq_head < 5'hD;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_26 = ldq_head < 5'hE;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_28 = ldq_head < 5'hF;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_32 = ldq_head < 5'h11;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_34 = ldq_head < 5'h12;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_36 = ldq_head < 5'h13;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_38 = ldq_head < 5'h14;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_40 = ldq_head < 5'h15;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_42 = ldq_head < 5'h16;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_44 = ldq_head < 5'h17;	// lsu.scala:215:29, util.scala:205:25, :351:72
    _temp_bits_T_46 = ldq_head[4:3] != 2'h3;	// lsu.scala:215:29, util.scala:351:72
    _stq_retry_idx_T = stq_0_bits_addr_valid & stq_0_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_1 = stq_1_bits_addr_valid & stq_1_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_2 = stq_2_bits_addr_valid & stq_2_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_3 = stq_3_bits_addr_valid & stq_3_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_4 = stq_4_bits_addr_valid & stq_4_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_5 = stq_5_bits_addr_valid & stq_5_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_6 = stq_6_bits_addr_valid & stq_6_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_7 = stq_7_bits_addr_valid & stq_7_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_8 = stq_8_bits_addr_valid & stq_8_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_9 = stq_9_bits_addr_valid & stq_9_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_10 = stq_10_bits_addr_valid & stq_10_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_11 = stq_11_bits_addr_valid & stq_11_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_12 = stq_12_bits_addr_valid & stq_12_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_13 = stq_13_bits_addr_valid & stq_13_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_14 = stq_14_bits_addr_valid & stq_14_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_15 = stq_15_bits_addr_valid & stq_15_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_16 = stq_16_bits_addr_valid & stq_16_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_17 = stq_17_bits_addr_valid & stq_17_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_18 = stq_18_bits_addr_valid & stq_18_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_19 = stq_19_bits_addr_valid & stq_19_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_20 = stq_20_bits_addr_valid & stq_20_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_21 = stq_21_bits_addr_valid & stq_21_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_22 = stq_22_bits_addr_valid & stq_22_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _ldq_wakeup_idx_T_7 =
      ldq_0_bits_addr_valid & ~ldq_0_bits_executed & ~ldq_0_bits_succeeded
      & ~ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_15 =
      ldq_1_bits_addr_valid & ~ldq_1_bits_executed & ~ldq_1_bits_succeeded
      & ~ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_23 =
      ldq_2_bits_addr_valid & ~ldq_2_bits_executed & ~ldq_2_bits_succeeded
      & ~ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_31 =
      ldq_3_bits_addr_valid & ~ldq_3_bits_executed & ~ldq_3_bits_succeeded
      & ~ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_39 =
      ldq_4_bits_addr_valid & ~ldq_4_bits_executed & ~ldq_4_bits_succeeded
      & ~ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_47 =
      ldq_5_bits_addr_valid & ~ldq_5_bits_executed & ~ldq_5_bits_succeeded
      & ~ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_55 =
      ldq_6_bits_addr_valid & ~ldq_6_bits_executed & ~ldq_6_bits_succeeded
      & ~ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_63 =
      ldq_7_bits_addr_valid & ~ldq_7_bits_executed & ~ldq_7_bits_succeeded
      & ~ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_71 =
      ldq_8_bits_addr_valid & ~ldq_8_bits_executed & ~ldq_8_bits_succeeded
      & ~ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_79 =
      ldq_9_bits_addr_valid & ~ldq_9_bits_executed & ~ldq_9_bits_succeeded
      & ~ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_87 =
      ldq_10_bits_addr_valid & ~ldq_10_bits_executed & ~ldq_10_bits_succeeded
      & ~ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_95 =
      ldq_11_bits_addr_valid & ~ldq_11_bits_executed & ~ldq_11_bits_succeeded
      & ~ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_103 =
      ldq_12_bits_addr_valid & ~ldq_12_bits_executed & ~ldq_12_bits_succeeded
      & ~ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_111 =
      ldq_13_bits_addr_valid & ~ldq_13_bits_executed & ~ldq_13_bits_succeeded
      & ~ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_119 =
      ldq_14_bits_addr_valid & ~ldq_14_bits_executed & ~ldq_14_bits_succeeded
      & ~ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_127 =
      ldq_15_bits_addr_valid & ~ldq_15_bits_executed & ~ldq_15_bits_succeeded
      & ~ldq_15_bits_addr_is_virtual & ~ldq_retry_idx_block_15;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_135 =
      ldq_16_bits_addr_valid & ~ldq_16_bits_executed & ~ldq_16_bits_succeeded
      & ~ldq_16_bits_addr_is_virtual & ~ldq_retry_idx_block_16;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_143 =
      ldq_17_bits_addr_valid & ~ldq_17_bits_executed & ~ldq_17_bits_succeeded
      & ~ldq_17_bits_addr_is_virtual & ~ldq_retry_idx_block_17;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_151 =
      ldq_18_bits_addr_valid & ~ldq_18_bits_executed & ~ldq_18_bits_succeeded
      & ~ldq_18_bits_addr_is_virtual & ~ldq_retry_idx_block_18;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_159 =
      ldq_19_bits_addr_valid & ~ldq_19_bits_executed & ~ldq_19_bits_succeeded
      & ~ldq_19_bits_addr_is_virtual & ~ldq_retry_idx_block_19;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_167 =
      ldq_20_bits_addr_valid & ~ldq_20_bits_executed & ~ldq_20_bits_succeeded
      & ~ldq_20_bits_addr_is_virtual & ~ldq_retry_idx_block_20;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_175 =
      ldq_21_bits_addr_valid & ~ldq_21_bits_executed & ~ldq_21_bits_succeeded
      & ~ldq_21_bits_addr_is_virtual & ~ldq_retry_idx_block_21;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_183 =
      ldq_22_bits_addr_valid & ~ldq_22_bits_executed & ~ldq_22_bits_succeeded
      & ~ldq_22_bits_addr_is_virtual & ~ldq_retry_idx_block_22;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    ma_st_0 = _stq_idx_T & io_core_exe_0_req_bits_mxcpt_valid;	// lsu.scala:660:{56,87}
    pf_ld_0 =
      ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_ld
      & _mem_xcpt_uops_WIRE_0_uses_ldq;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :661:75
    pf_st_0 =
      ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_st
      & _mem_xcpt_uops_WIRE_0_uses_stq;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :662:75
    ae_ld_0 =
      ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_ae_ld
      & _mem_xcpt_uops_WIRE_0_uses_ldq;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :663:75
    dmem_req_fire_0 = dmem_req_0_valid & io_dmem_req_ready;	// lsu.scala:752:55, :766:39, :767:30, :773:43
    ldq_idx =
      can_fire_load_incoming_0 ? io_core_exe_0_req_bits_uop_ldq_idx : ldq_retry_idx;	// lsu.scala:415:30, :441:63, :837:24
    _GEN_1243 = _GEN_315 & ldq_idx == 5'h0;	// lsu.scala:220:29, :304:5, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1244 =
      _GEN_1243 | ~_GEN_1051
      & (dis_ld_val_1
           ? ~_GEN_930 & ldq_0_bits_addr_valid
           : ~_GEN_855 & ldq_0_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1245 = _GEN_315 & ldq_idx == 5'h1;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1246 =
      _GEN_1245 | ~_GEN_1053
      & (dis_ld_val_1
           ? ~_GEN_932 & ldq_1_bits_addr_valid
           : ~_GEN_856 & ldq_1_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1247 = _GEN_315 & ldq_idx == 5'h2;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1248 =
      _GEN_1247 | ~_GEN_1055
      & (dis_ld_val_1
           ? ~_GEN_934 & ldq_2_bits_addr_valid
           : ~_GEN_857 & ldq_2_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1249 = _GEN_315 & ldq_idx == 5'h3;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1250 =
      _GEN_1249 | ~_GEN_1057
      & (dis_ld_val_1
           ? ~_GEN_936 & ldq_3_bits_addr_valid
           : ~_GEN_858 & ldq_3_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1251 = _GEN_315 & ldq_idx == 5'h4;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1252 =
      _GEN_1251 | ~_GEN_1059
      & (dis_ld_val_1
           ? ~_GEN_938 & ldq_4_bits_addr_valid
           : ~_GEN_859 & ldq_4_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1253 = _GEN_315 & ldq_idx == 5'h5;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1254 =
      _GEN_1253 | ~_GEN_1061
      & (dis_ld_val_1
           ? ~_GEN_940 & ldq_5_bits_addr_valid
           : ~_GEN_860 & ldq_5_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1255 = _GEN_315 & ldq_idx == 5'h6;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1256 =
      _GEN_1255 | ~_GEN_1063
      & (dis_ld_val_1
           ? ~_GEN_942 & ldq_6_bits_addr_valid
           : ~_GEN_861 & ldq_6_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1257 = _GEN_315 & ldq_idx == 5'h7;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1258 =
      _GEN_1257 | ~_GEN_1065
      & (dis_ld_val_1
           ? ~_GEN_944 & ldq_7_bits_addr_valid
           : ~_GEN_862 & ldq_7_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1259 = _GEN_315 & ldq_idx == 5'h8;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1260 =
      _GEN_1259 | ~_GEN_1067
      & (dis_ld_val_1
           ? ~_GEN_946 & ldq_8_bits_addr_valid
           : ~_GEN_863 & ldq_8_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1261 = _GEN_315 & ldq_idx == 5'h9;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1262 =
      _GEN_1261 | ~_GEN_1069
      & (dis_ld_val_1
           ? ~_GEN_948 & ldq_9_bits_addr_valid
           : ~_GEN_864 & ldq_9_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1263 = _GEN_315 & ldq_idx == 5'hA;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1264 =
      _GEN_1263 | ~_GEN_1071
      & (dis_ld_val_1
           ? ~_GEN_950 & ldq_10_bits_addr_valid
           : ~_GEN_865 & ldq_10_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1265 = _GEN_315 & ldq_idx == 5'hB;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1266 =
      _GEN_1265 | ~_GEN_1073
      & (dis_ld_val_1
           ? ~_GEN_952 & ldq_11_bits_addr_valid
           : ~_GEN_866 & ldq_11_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1267 = _GEN_315 & ldq_idx == 5'hC;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1268 =
      _GEN_1267 | ~_GEN_1075
      & (dis_ld_val_1
           ? ~_GEN_954 & ldq_12_bits_addr_valid
           : ~_GEN_867 & ldq_12_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1269 = _GEN_315 & ldq_idx == 5'hD;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1270 =
      _GEN_1269 | ~_GEN_1077
      & (dis_ld_val_1
           ? ~_GEN_956 & ldq_13_bits_addr_valid
           : ~_GEN_868 & ldq_13_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1271 = _GEN_315 & ldq_idx == 5'hE;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1272 =
      _GEN_1271 | ~_GEN_1079
      & (dis_ld_val_1
           ? ~_GEN_958 & ldq_14_bits_addr_valid
           : ~_GEN_869 & ldq_14_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1273 = _GEN_315 & ldq_idx == 5'hF;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1274 =
      _GEN_1273 | ~_GEN_1081
      & (dis_ld_val_1
           ? ~_GEN_960 & ldq_15_bits_addr_valid
           : ~_GEN_870 & ldq_15_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1275 = _GEN_315 & ldq_idx == 5'h10;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1276 =
      _GEN_1275 | ~_GEN_1083
      & (dis_ld_val_1
           ? ~_GEN_962 & ldq_16_bits_addr_valid
           : ~_GEN_871 & ldq_16_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1277 = _GEN_315 & ldq_idx == 5'h11;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1278 =
      _GEN_1277 | ~_GEN_1085
      & (dis_ld_val_1
           ? ~_GEN_964 & ldq_17_bits_addr_valid
           : ~_GEN_872 & ldq_17_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1279 = _GEN_315 & ldq_idx == 5'h12;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1280 =
      _GEN_1279 | ~_GEN_1087
      & (dis_ld_val_1
           ? ~_GEN_966 & ldq_18_bits_addr_valid
           : ~_GEN_873 & ldq_18_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1281 = _GEN_315 & ldq_idx == 5'h13;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1282 =
      _GEN_1281 | ~_GEN_1089
      & (dis_ld_val_1
           ? ~_GEN_968 & ldq_19_bits_addr_valid
           : ~_GEN_874 & ldq_19_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1283 = _GEN_315 & ldq_idx == 5'h14;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1284 =
      _GEN_1283 | ~_GEN_1091
      & (dis_ld_val_1
           ? ~_GEN_970 & ldq_20_bits_addr_valid
           : ~_GEN_875 & ldq_20_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1285 = _GEN_315 & ldq_idx == 5'h15;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1286 =
      _GEN_1285 | ~_GEN_1093
      & (dis_ld_val_1
           ? ~_GEN_972 & ldq_21_bits_addr_valid
           : ~_GEN_876 & ldq_21_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1287 = _GEN_315 & ldq_idx == 5'h16;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_1288 =
      _GEN_1287 | ~_GEN_1095
      & (dis_ld_val_1
           ? ~_GEN_974 & ldq_22_bits_addr_valid
           : ~_GEN_877 & ldq_22_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_1289 = _GEN_315 & ldq_idx == 5'h17;	// lsu.scala:220:29, :304:5, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45, util.scala:205:25
    _GEN_1290 =
      _GEN_1289 | ~_GEN_1097
      & (dis_ld_val_1
           ? ~_GEN_976 & ldq_23_bits_addr_valid
           : ~_GEN_878 & ldq_23_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _ldq_bits_addr_is_uncacheable_T_1 = ~_dtlb_io_resp_0_cacheable & ~exe_tlb_miss_0;	// lsu.scala:249:20, :708:58, :711:43, :842:{71,74}
    stq_idx = _stq_idx_T ? io_core_exe_0_req_bits_uop_stq_idx : stq_retry_idx;	// lsu.scala:422:30, :660:56, :850:24
    _GEN_1291 = _GEN_321 & stq_idx == 5'h0;	// lsu.scala:304:5, :848:67, :849:5, :850:24, :853:36
    _GEN_1292 =
      _GEN_1291 ? ~pf_st_0 : _GEN_1195 & _GEN_1025 & _GEN_903 & stq_0_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1293 = _GEN_321 & stq_idx == 5'h1;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1294 =
      _GEN_1293 ? ~pf_st_0 : _GEN_1196 & _GEN_1026 & _GEN_904 & stq_1_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1295 = _GEN_321 & stq_idx == 5'h2;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1296 =
      _GEN_1295 ? ~pf_st_0 : _GEN_1197 & _GEN_1027 & _GEN_905 & stq_2_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1297 = _GEN_321 & stq_idx == 5'h3;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1298 =
      _GEN_1297 ? ~pf_st_0 : _GEN_1198 & _GEN_1028 & _GEN_906 & stq_3_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1299 = _GEN_321 & stq_idx == 5'h4;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1300 =
      _GEN_1299 ? ~pf_st_0 : _GEN_1199 & _GEN_1029 & _GEN_907 & stq_4_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1301 = _GEN_321 & stq_idx == 5'h5;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1302 =
      _GEN_1301 ? ~pf_st_0 : _GEN_1200 & _GEN_1030 & _GEN_908 & stq_5_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1303 = _GEN_321 & stq_idx == 5'h6;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1304 =
      _GEN_1303 ? ~pf_st_0 : _GEN_1201 & _GEN_1031 & _GEN_909 & stq_6_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1305 = _GEN_321 & stq_idx == 5'h7;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1306 =
      _GEN_1305 ? ~pf_st_0 : _GEN_1202 & _GEN_1032 & _GEN_910 & stq_7_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1307 = _GEN_321 & stq_idx == 5'h8;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1308 =
      _GEN_1307 ? ~pf_st_0 : _GEN_1203 & _GEN_1033 & _GEN_911 & stq_8_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1309 = _GEN_321 & stq_idx == 5'h9;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1310 =
      _GEN_1309 ? ~pf_st_0 : _GEN_1204 & _GEN_1034 & _GEN_912 & stq_9_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1311 = _GEN_321 & stq_idx == 5'hA;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1312 =
      _GEN_1311 ? ~pf_st_0 : _GEN_1205 & _GEN_1035 & _GEN_913 & stq_10_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1313 = _GEN_321 & stq_idx == 5'hB;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1314 =
      _GEN_1313 ? ~pf_st_0 : _GEN_1206 & _GEN_1036 & _GEN_914 & stq_11_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1315 = _GEN_321 & stq_idx == 5'hC;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1316 =
      _GEN_1315 ? ~pf_st_0 : _GEN_1207 & _GEN_1037 & _GEN_915 & stq_12_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1317 = _GEN_321 & stq_idx == 5'hD;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1318 =
      _GEN_1317 ? ~pf_st_0 : _GEN_1208 & _GEN_1038 & _GEN_916 & stq_13_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1319 = _GEN_321 & stq_idx == 5'hE;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1320 =
      _GEN_1319 ? ~pf_st_0 : _GEN_1209 & _GEN_1039 & _GEN_917 & stq_14_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1321 = _GEN_321 & stq_idx == 5'hF;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1322 =
      _GEN_1321 ? ~pf_st_0 : _GEN_1210 & _GEN_1040 & _GEN_918 & stq_15_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1323 = _GEN_321 & stq_idx == 5'h10;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1324 =
      _GEN_1323 ? ~pf_st_0 : _GEN_1211 & _GEN_1041 & _GEN_919 & stq_16_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1325 = _GEN_321 & stq_idx == 5'h11;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1326 =
      _GEN_1325 ? ~pf_st_0 : _GEN_1212 & _GEN_1042 & _GEN_920 & stq_17_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1327 = _GEN_321 & stq_idx == 5'h12;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1328 =
      _GEN_1327 ? ~pf_st_0 : _GEN_1213 & _GEN_1043 & _GEN_921 & stq_18_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1329 = _GEN_321 & stq_idx == 5'h13;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1330 =
      _GEN_1329 ? ~pf_st_0 : _GEN_1214 & _GEN_1044 & _GEN_922 & stq_19_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1331 = _GEN_321 & stq_idx == 5'h14;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1332 =
      _GEN_1331 ? ~pf_st_0 : _GEN_1215 & _GEN_1045 & _GEN_923 & stq_20_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1333 = _GEN_321 & stq_idx == 5'h15;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1334 =
      _GEN_1333 ? ~pf_st_0 : _GEN_1216 & _GEN_1046 & _GEN_924 & stq_21_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1335 = _GEN_321 & stq_idx == 5'h16;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_1336 =
      _GEN_1335 ? ~pf_st_0 : _GEN_1217 & _GEN_1047 & _GEN_925 & stq_22_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1337 = _GEN_321 & stq_idx == 5'h17;	// lsu.scala:304:5, :848:67, :849:5, :850:24, :853:36, util.scala:205:25
    _GEN_1338 =
      _GEN_1337 ? ~pf_st_0 : _GEN_1218 & _GEN_1048 & _GEN_926 & stq_23_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_1340 = _GEN_1339 | _GEN_1195 & _GEN_1025 & _GEN_903 & stq_0_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1342 = _GEN_1341 | _GEN_1196 & _GEN_1026 & _GEN_904 & stq_1_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1344 = _GEN_1343 | _GEN_1197 & _GEN_1027 & _GEN_905 & stq_2_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1346 = _GEN_1345 | _GEN_1198 & _GEN_1028 & _GEN_906 & stq_3_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1348 = _GEN_1347 | _GEN_1199 & _GEN_1029 & _GEN_907 & stq_4_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1350 = _GEN_1349 | _GEN_1200 & _GEN_1030 & _GEN_908 & stq_5_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1352 = _GEN_1351 | _GEN_1201 & _GEN_1031 & _GEN_909 & stq_6_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1354 = _GEN_1353 | _GEN_1202 & _GEN_1032 & _GEN_910 & stq_7_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1356 = _GEN_1355 | _GEN_1203 & _GEN_1033 & _GEN_911 & stq_8_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1358 = _GEN_1357 | _GEN_1204 & _GEN_1034 & _GEN_912 & stq_9_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1360 = _GEN_1359 | _GEN_1205 & _GEN_1035 & _GEN_913 & stq_10_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1362 = _GEN_1361 | _GEN_1206 & _GEN_1036 & _GEN_914 & stq_11_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1364 = _GEN_1363 | _GEN_1207 & _GEN_1037 & _GEN_915 & stq_12_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1366 = _GEN_1365 | _GEN_1208 & _GEN_1038 & _GEN_916 & stq_13_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1368 = _GEN_1367 | _GEN_1209 & _GEN_1039 & _GEN_917 & stq_14_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1370 = _GEN_1369 | _GEN_1210 & _GEN_1040 & _GEN_918 & stq_15_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1372 = _GEN_1371 | _GEN_1211 & _GEN_1041 & _GEN_919 & stq_16_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1374 = _GEN_1373 | _GEN_1212 & _GEN_1042 & _GEN_920 & stq_17_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1376 = _GEN_1375 | _GEN_1213 & _GEN_1043 & _GEN_921 & stq_18_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1378 = _GEN_1377 | _GEN_1214 & _GEN_1044 & _GEN_922 & stq_19_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1380 = _GEN_1379 | _GEN_1215 & _GEN_1045 & _GEN_923 & stq_20_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1382 = _GEN_1381 | _GEN_1216 & _GEN_1046 & _GEN_924 & stq_21_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1384 = _GEN_1383 | _GEN_1217 & _GEN_1047 & _GEN_925 & stq_22_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_1386 = _GEN_1385 | _GEN_1218 & _GEN_1048 & _GEN_926 & stq_23_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    l_forward_stq_idx =
      l_forwarders_0 ? wb_forward_stq_idx_0 : ldq_0_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1387 =
      ~ldq_0_bits_forward_std_val | l_forward_stq_idx != lcam_stq_idx_0
      & (l_forward_stq_idx < lcam_stq_idx_0
         ^ l_forward_stq_idx < ldq_0_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_0_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1388 = _GEN_329 & ~s1_executing_loads_0 & ldq_0_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_24 =
      ~_GEN_327 & (_GEN_332 ? _GEN_1387 : _GEN_333 & searcher_is_older & _GEN_1388);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_1 =
      l_forwarders_1_0 ? wb_forward_stq_idx_0 : ldq_1_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1412 =
      ~ldq_1_bits_forward_std_val | l_forward_stq_idx_1 != lcam_stq_idx_0
      & (l_forward_stq_idx_1 < lcam_stq_idx_0
         ^ l_forward_stq_idx_1 < ldq_1_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_1_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1413 = _GEN_340 & ~s1_executing_loads_1 & ldq_1_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_25 =
      ~_GEN_338 & (_GEN_342 ? _GEN_1412 : _GEN_343 & searcher_is_older_1 & _GEN_1413);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_2 =
      l_forwarders_2_0 ? wb_forward_stq_idx_0 : ldq_2_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1414 =
      ~ldq_2_bits_forward_std_val | l_forward_stq_idx_2 != lcam_stq_idx_0
      & (l_forward_stq_idx_2 < lcam_stq_idx_0
         ^ l_forward_stq_idx_2 < ldq_2_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_2_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1415 = _GEN_351 & ~s1_executing_loads_2 & ldq_2_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_26 =
      ~_GEN_349 & (_GEN_353 ? _GEN_1414 : _GEN_354 & searcher_is_older_2 & _GEN_1415);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_3 =
      l_forwarders_3_0 ? wb_forward_stq_idx_0 : ldq_3_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1416 =
      ~ldq_3_bits_forward_std_val | l_forward_stq_idx_3 != lcam_stq_idx_0
      & (l_forward_stq_idx_3 < lcam_stq_idx_0
         ^ l_forward_stq_idx_3 < ldq_3_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_3_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1417 = _GEN_362 & ~s1_executing_loads_3 & ldq_3_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_27 =
      ~_GEN_360 & (_GEN_364 ? _GEN_1416 : _GEN_365 & searcher_is_older_3 & _GEN_1417);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_4 =
      l_forwarders_4_0 ? wb_forward_stq_idx_0 : ldq_4_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1418 =
      ~ldq_4_bits_forward_std_val | l_forward_stq_idx_4 != lcam_stq_idx_0
      & (l_forward_stq_idx_4 < lcam_stq_idx_0
         ^ l_forward_stq_idx_4 < ldq_4_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_4_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1419 = _GEN_373 & ~s1_executing_loads_4 & ldq_4_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_28 =
      ~_GEN_371 & (_GEN_375 ? _GEN_1418 : _GEN_376 & searcher_is_older_4 & _GEN_1419);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_5 =
      l_forwarders_5_0 ? wb_forward_stq_idx_0 : ldq_5_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1420 =
      ~ldq_5_bits_forward_std_val | l_forward_stq_idx_5 != lcam_stq_idx_0
      & (l_forward_stq_idx_5 < lcam_stq_idx_0
         ^ l_forward_stq_idx_5 < ldq_5_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_5_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1421 = _GEN_384 & ~s1_executing_loads_5 & ldq_5_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_29 =
      ~_GEN_382 & (_GEN_386 ? _GEN_1420 : _GEN_387 & searcher_is_older_5 & _GEN_1421);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_6 =
      l_forwarders_6_0 ? wb_forward_stq_idx_0 : ldq_6_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1422 =
      ~ldq_6_bits_forward_std_val | l_forward_stq_idx_6 != lcam_stq_idx_0
      & (l_forward_stq_idx_6 < lcam_stq_idx_0
         ^ l_forward_stq_idx_6 < ldq_6_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_6_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1423 = _GEN_395 & ~s1_executing_loads_6 & ldq_6_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_30 =
      ~_GEN_393 & (_GEN_397 ? _GEN_1422 : _GEN_398 & searcher_is_older_6 & _GEN_1423);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_7 =
      l_forwarders_7_0 ? wb_forward_stq_idx_0 : ldq_7_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1424 =
      ~ldq_7_bits_forward_std_val | l_forward_stq_idx_7 != lcam_stq_idx_0
      & (l_forward_stq_idx_7 < lcam_stq_idx_0
         ^ l_forward_stq_idx_7 < ldq_7_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_7_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1425 = _GEN_406 & ~s1_executing_loads_7 & ldq_7_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_31 =
      ~_GEN_404 & (_GEN_408 ? _GEN_1424 : _GEN_409 & searcher_is_older_7 & _GEN_1425);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_8 =
      l_forwarders_8_0 ? wb_forward_stq_idx_0 : ldq_8_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1426 =
      ~ldq_8_bits_forward_std_val | l_forward_stq_idx_8 != lcam_stq_idx_0
      & (l_forward_stq_idx_8 < lcam_stq_idx_0
         ^ l_forward_stq_idx_8 < ldq_8_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_8_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1427 = _GEN_417 & ~s1_executing_loads_8 & ldq_8_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_32 =
      ~_GEN_415 & (_GEN_419 ? _GEN_1426 : _GEN_420 & searcher_is_older_8 & _GEN_1427);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_9 =
      l_forwarders_9_0 ? wb_forward_stq_idx_0 : ldq_9_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1428 =
      ~ldq_9_bits_forward_std_val | l_forward_stq_idx_9 != lcam_stq_idx_0
      & (l_forward_stq_idx_9 < lcam_stq_idx_0
         ^ l_forward_stq_idx_9 < ldq_9_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_9_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1429 = _GEN_428 & ~s1_executing_loads_9 & ldq_9_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_33 =
      ~_GEN_426 & (_GEN_430 ? _GEN_1428 : _GEN_431 & searcher_is_older_9 & _GEN_1429);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_10 =
      l_forwarders_10_0 ? wb_forward_stq_idx_0 : ldq_10_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1430 =
      ~ldq_10_bits_forward_std_val | l_forward_stq_idx_10 != lcam_stq_idx_0
      & (l_forward_stq_idx_10 < lcam_stq_idx_0
         ^ l_forward_stq_idx_10 < ldq_10_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_10_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1431 = _GEN_439 & ~s1_executing_loads_10 & ldq_10_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_34 =
      ~_GEN_437 & (_GEN_441 ? _GEN_1430 : _GEN_442 & searcher_is_older_10 & _GEN_1431);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_11 =
      l_forwarders_11_0 ? wb_forward_stq_idx_0 : ldq_11_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1432 =
      ~ldq_11_bits_forward_std_val | l_forward_stq_idx_11 != lcam_stq_idx_0
      & (l_forward_stq_idx_11 < lcam_stq_idx_0
         ^ l_forward_stq_idx_11 < ldq_11_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_11_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1433 = _GEN_450 & ~s1_executing_loads_11 & ldq_11_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_35 =
      ~_GEN_448 & (_GEN_452 ? _GEN_1432 : _GEN_453 & searcher_is_older_11 & _GEN_1433);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_12 =
      l_forwarders_12_0 ? wb_forward_stq_idx_0 : ldq_12_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1434 =
      ~ldq_12_bits_forward_std_val | l_forward_stq_idx_12 != lcam_stq_idx_0
      & (l_forward_stq_idx_12 < lcam_stq_idx_0
         ^ l_forward_stq_idx_12 < ldq_12_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_12_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1435 = _GEN_461 & ~s1_executing_loads_12 & ldq_12_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_36 =
      ~_GEN_459 & (_GEN_463 ? _GEN_1434 : _GEN_464 & searcher_is_older_12 & _GEN_1435);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_13 =
      l_forwarders_13_0 ? wb_forward_stq_idx_0 : ldq_13_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1436 =
      ~ldq_13_bits_forward_std_val | l_forward_stq_idx_13 != lcam_stq_idx_0
      & (l_forward_stq_idx_13 < lcam_stq_idx_0
         ^ l_forward_stq_idx_13 < ldq_13_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_13_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1437 = _GEN_472 & ~s1_executing_loads_13 & ldq_13_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_37 =
      ~_GEN_470 & (_GEN_474 ? _GEN_1436 : _GEN_475 & searcher_is_older_13 & _GEN_1437);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_14 =
      l_forwarders_14_0 ? wb_forward_stq_idx_0 : ldq_14_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1438 =
      ~ldq_14_bits_forward_std_val | l_forward_stq_idx_14 != lcam_stq_idx_0
      & (l_forward_stq_idx_14 < lcam_stq_idx_0
         ^ l_forward_stq_idx_14 < ldq_14_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_14_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1439 = _GEN_483 & ~s1_executing_loads_14 & ldq_14_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_38 =
      ~_GEN_481 & (_GEN_485 ? _GEN_1438 : _GEN_486 & searcher_is_older_14 & _GEN_1439);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_15 =
      l_forwarders_15_0 ? wb_forward_stq_idx_0 : ldq_15_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1440 =
      ~ldq_15_bits_forward_std_val | l_forward_stq_idx_15 != lcam_stq_idx_0
      & (l_forward_stq_idx_15 < lcam_stq_idx_0
         ^ l_forward_stq_idx_15 < ldq_15_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_15_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1441 = _GEN_494 & ~s1_executing_loads_15 & ldq_15_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_39 =
      ~_GEN_492 & (_GEN_496 ? _GEN_1440 : _GEN_497 & searcher_is_older_15 & _GEN_1441);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_16 =
      l_forwarders_16_0 ? wb_forward_stq_idx_0 : ldq_16_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1442 =
      ~ldq_16_bits_forward_std_val | l_forward_stq_idx_16 != lcam_stq_idx_0
      & (l_forward_stq_idx_16 < lcam_stq_idx_0
         ^ l_forward_stq_idx_16 < ldq_16_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_16_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1443 = _GEN_505 & ~s1_executing_loads_16 & ldq_16_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_40 =
      ~_GEN_503 & (_GEN_507 ? _GEN_1442 : _GEN_508 & searcher_is_older_16 & _GEN_1443);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_17 =
      l_forwarders_17_0 ? wb_forward_stq_idx_0 : ldq_17_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1444 =
      ~ldq_17_bits_forward_std_val | l_forward_stq_idx_17 != lcam_stq_idx_0
      & (l_forward_stq_idx_17 < lcam_stq_idx_0
         ^ l_forward_stq_idx_17 < ldq_17_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_17_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1445 = _GEN_516 & ~s1_executing_loads_17 & ldq_17_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_41 =
      ~_GEN_514 & (_GEN_518 ? _GEN_1444 : _GEN_519 & searcher_is_older_17 & _GEN_1445);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_18 =
      l_forwarders_18_0 ? wb_forward_stq_idx_0 : ldq_18_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1446 =
      ~ldq_18_bits_forward_std_val | l_forward_stq_idx_18 != lcam_stq_idx_0
      & (l_forward_stq_idx_18 < lcam_stq_idx_0
         ^ l_forward_stq_idx_18 < ldq_18_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_18_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1447 = _GEN_527 & ~s1_executing_loads_18 & ldq_18_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_42 =
      ~_GEN_525 & (_GEN_529 ? _GEN_1446 : _GEN_530 & searcher_is_older_18 & _GEN_1447);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_19 =
      l_forwarders_19_0 ? wb_forward_stq_idx_0 : ldq_19_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1448 =
      ~ldq_19_bits_forward_std_val | l_forward_stq_idx_19 != lcam_stq_idx_0
      & (l_forward_stq_idx_19 < lcam_stq_idx_0
         ^ l_forward_stq_idx_19 < ldq_19_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_19_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1449 = _GEN_538 & ~s1_executing_loads_19 & ldq_19_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_43 =
      ~_GEN_536 & (_GEN_540 ? _GEN_1448 : _GEN_541 & searcher_is_older_19 & _GEN_1449);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_20 =
      l_forwarders_20_0 ? wb_forward_stq_idx_0 : ldq_20_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1450 =
      ~ldq_20_bits_forward_std_val | l_forward_stq_idx_20 != lcam_stq_idx_0
      & (l_forward_stq_idx_20 < lcam_stq_idx_0
         ^ l_forward_stq_idx_20 < ldq_20_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_20_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1451 = _GEN_549 & ~s1_executing_loads_20 & ldq_20_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_44 =
      ~_GEN_547 & (_GEN_551 ? _GEN_1450 : _GEN_552 & searcher_is_older_20 & _GEN_1451);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_21 =
      l_forwarders_21_0 ? wb_forward_stq_idx_0 : ldq_21_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1452 =
      ~ldq_21_bits_forward_std_val | l_forward_stq_idx_21 != lcam_stq_idx_0
      & (l_forward_stq_idx_21 < lcam_stq_idx_0
         ^ l_forward_stq_idx_21 < ldq_21_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_21_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1453 = _GEN_560 & ~s1_executing_loads_21 & ldq_21_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_45 =
      ~_GEN_558 & (_GEN_562 ? _GEN_1452 : _GEN_563 & searcher_is_older_21 & _GEN_1453);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_22 =
      l_forwarders_22_0 ? wb_forward_stq_idx_0 : ldq_22_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1454 =
      ~ldq_22_bits_forward_std_val | l_forward_stq_idx_22 != lcam_stq_idx_0
      & (l_forward_stq_idx_22 < lcam_stq_idx_0
         ^ l_forward_stq_idx_22 < ldq_22_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_22_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1455 = _GEN_571 & ~s1_executing_loads_22 & ldq_22_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_46 =
      ~_GEN_569 & (_GEN_573 ? _GEN_1454 : _GEN_574 & searcher_is_older_22 & _GEN_1455);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_23 =
      l_forwarders_23_0 ? wb_forward_stq_idx_0 : ldq_23_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_1456 =
      ~ldq_23_bits_forward_std_val | l_forward_stq_idx_23 != lcam_stq_idx_0
      & (l_forward_stq_idx_23 < lcam_stq_idx_0
         ^ l_forward_stq_idx_23 < ldq_23_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_23_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_1457 = _GEN_582 & ~s1_executing_loads_23 & ldq_23_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_47 =
      ~_GEN_580 & (_GEN_584 ? _GEN_1456 : _GEN_585 & searcher_is_older_23 & _GEN_1457);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    _GEN_1458 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23
       | ~(_GEN_586 & _GEN_587 & ~(|lcam_ldq_idx_0)))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22
         | ~(_GEN_575 & _GEN_576 & ~(|lcam_ldq_idx_0)))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21
         | ~(_GEN_564 & _GEN_565 & ~(|lcam_ldq_idx_0)))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20
         | ~(_GEN_553 & _GEN_554 & ~(|lcam_ldq_idx_0)))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19
         | ~(_GEN_542 & _GEN_543 & ~(|lcam_ldq_idx_0)))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18
         | ~(_GEN_531 & _GEN_532 & ~(|lcam_ldq_idx_0)))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17
         | ~(_GEN_520 & _GEN_521 & ~(|lcam_ldq_idx_0)))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16
         | ~(_GEN_509 & _GEN_510 & ~(|lcam_ldq_idx_0)))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15
         | ~(_GEN_498 & _GEN_499 & ~(|lcam_ldq_idx_0)))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14
         | ~(_GEN_487 & _GEN_488 & ~(|lcam_ldq_idx_0)))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13
         | ~(_GEN_476 & _GEN_477 & ~(|lcam_ldq_idx_0)))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12
         | ~(_GEN_465 & _GEN_466 & ~(|lcam_ldq_idx_0)))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11
         | ~(_GEN_454 & _GEN_455 & ~(|lcam_ldq_idx_0)))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10
         | ~(_GEN_443 & _GEN_444 & ~(|lcam_ldq_idx_0)))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9
         | ~(_GEN_432 & _GEN_433 & ~(|lcam_ldq_idx_0)))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8
         | ~(_GEN_421 & _GEN_422 & ~(|lcam_ldq_idx_0)))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7
         | ~(_GEN_410 & _GEN_411 & ~(|lcam_ldq_idx_0)))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6
         | ~(_GEN_399 & _GEN_400 & ~(|lcam_ldq_idx_0)))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5
         | ~(_GEN_388 & _GEN_389 & ~(|lcam_ldq_idx_0)))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4
         | ~(_GEN_377 & _GEN_378 & ~(|lcam_ldq_idx_0)))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3
         | ~(_GEN_366 & _GEN_367 & ~(|lcam_ldq_idx_0)))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2
         | ~(_GEN_355 & _GEN_356 & ~(|lcam_ldq_idx_0)))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1
         | ~(_GEN_344 & _GEN_345 & ~(|lcam_ldq_idx_0))) & s1_executing_loads_0;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1459 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1389))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1389))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1389))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1389))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1389))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1389))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1389))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1389))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1389))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1389))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1389))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1389))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1389))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1389))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1389))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1389))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1389))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1389))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1389))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1389))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1389))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1389))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1389))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1389)) & s1_executing_loads_1;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1460 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1390))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1390))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1390))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1390))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1390))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1390))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1390))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1390))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1390))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1390))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1390))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1390))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1390))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1390))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1390))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1390))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1390))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1390))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1390))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1390))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1390))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1390))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1390))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1390)) & s1_executing_loads_2;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1461 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1391))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1391))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1391))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1391))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1391))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1391))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1391))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1391))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1391))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1391))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1391))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1391))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1391))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1391))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1391))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1391))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1391))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1391))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1391))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1391))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1391))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1391))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1391))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1391)) & s1_executing_loads_3;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1462 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1392))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1392))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1392))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1392))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1392))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1392))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1392))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1392))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1392))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1392))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1392))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1392))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1392))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1392))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1392))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1392))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1392))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1392))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1392))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1392))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1392))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1392))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1392))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1392)) & s1_executing_loads_4;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1463 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1393))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1393))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1393))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1393))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1393))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1393))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1393))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1393))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1393))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1393))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1393))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1393))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1393))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1393))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1393))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1393))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1393))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1393))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1393))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1393))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1393))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1393))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1393))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1393)) & s1_executing_loads_5;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1464 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1394))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1394))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1394))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1394))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1394))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1394))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1394))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1394))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1394))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1394))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1394))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1394))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1394))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1394))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1394))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1394))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1394))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1394))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1394))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1394))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1394))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1394))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1394))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1394)) & s1_executing_loads_6;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1465 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1395))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1395))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1395))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1395))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1395))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1395))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1395))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1395))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1395))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1395))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1395))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1395))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1395))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1395))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1395))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1395))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1395))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1395))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1395))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1395))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1395))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1395))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1395))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1395)) & s1_executing_loads_7;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1466 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1396))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1396))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1396))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1396))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1396))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1396))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1396))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1396))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1396))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1396))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1396))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1396))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1396))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1396))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1396))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1396))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1396))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1396))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1396))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1396))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1396))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1396))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1396))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1396)) & s1_executing_loads_8;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1467 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1397))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1397))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1397))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1397))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1397))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1397))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1397))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1397))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1397))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1397))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1397))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1397))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1397))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1397))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1397))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1397))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1397))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1397))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1397))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1397))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1397))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1397))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1397))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1397)) & s1_executing_loads_9;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1468 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1398))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1398))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1398))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1398))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1398))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1398))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1398))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1398))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1398))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1398))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1398))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1398))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1398))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1398))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1398))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1398))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1398))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1398))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1398))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1398))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1398))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1398))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1398))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1398)) & s1_executing_loads_10;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1469 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1399))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1399))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1399))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1399))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1399))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1399))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1399))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1399))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1399))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1399))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1399))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1399))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1399))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1399))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1399))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1399))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1399))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1399))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1399))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1399))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1399))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1399))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1399))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1399)) & s1_executing_loads_11;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1470 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1400))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1400))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1400))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1400))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1400))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1400))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1400))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1400))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1400))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1400))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1400))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1400))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1400))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1400))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1400))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1400))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1400))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1400))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1400))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1400))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1400))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1400))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1400))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1400)) & s1_executing_loads_12;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1471 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1401))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1401))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1401))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1401))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1401))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1401))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1401))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1401))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1401))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1401))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1401))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1401))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1401))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1401))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1401))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1401))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1401))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1401))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1401))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1401))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1401))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1401))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1401))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1401)) & s1_executing_loads_13;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1472 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1402))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1402))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1402))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1402))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1402))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1402))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1402))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1402))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1402))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1402))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1402))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1402))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1402))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1402))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1402))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1402))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1402))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1402))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1402))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1402))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1402))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1402))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1402))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1402)) & s1_executing_loads_14;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1473 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1403))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1403))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1403))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1403))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1403))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1403))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1403))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1403))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1403))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1403))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1403))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1403))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1403))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1403))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1403))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1403))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1403))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1403))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1403))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1403))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1403))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1403))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1403))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1403)) & s1_executing_loads_15;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1474 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1404))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1404))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1404))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1404))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1404))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1404))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1404))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1404))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1404))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1404))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1404))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1404))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1404))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1404))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1404))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1404))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1404))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1404))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1404))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1404))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1404))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1404))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1404))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1404)) & s1_executing_loads_16;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1475 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1405))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1405))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1405))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1405))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1405))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1405))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1405))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1405))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1405))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1405))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1405))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1405))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1405))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1405))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1405))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1405))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1405))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1405))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1405))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1405))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1405))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1405))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1405))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1405)) & s1_executing_loads_17;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1476 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1406))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1406))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1406))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1406))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1406))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1406))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1406))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1406))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1406))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1406))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1406))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1406))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1406))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1406))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1406))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1406))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1406))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1406))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1406))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1406))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1406))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1406))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1406))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1406)) & s1_executing_loads_18;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1477 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1407))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1407))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1407))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1407))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1407))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1407))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1407))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1407))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1407))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1407))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1407))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1407))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1407))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1407))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1407))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1407))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1407))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1407))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1407))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1407))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1407))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1407))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1407))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1407)) & s1_executing_loads_19;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1478 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1408))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1408))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1408))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1408))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1408))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1408))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1408))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1408))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1408))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1408))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1408))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1408))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1408))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1408))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1408))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1408))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1408))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1408))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1408))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1408))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1408))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1408))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1408))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1408)) & s1_executing_loads_20;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1479 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1409))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1409))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1409))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1409))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1409))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1409))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1409))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1409))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1409))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1409))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1409))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1409))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1409))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1409))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1409))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1409))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1409))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1409))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1409))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1409))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1409))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1409))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1409))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1409)) & s1_executing_loads_21;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1480 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1410))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1410))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1410))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1410))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1410))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1410))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1410))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1410))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1410))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1410))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1410))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1410))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1410))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1410))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1410))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1410))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1410))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1410))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1410))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1410))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1410))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1410))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1410))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1410)) & s1_executing_loads_22;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1481 =
      (_GEN_588 | ~_GEN_585 | searcher_is_older_23 | ~(_GEN_586 & _GEN_587 & _GEN_1411))
      & (_GEN_577 | ~_GEN_574 | searcher_is_older_22 | ~(_GEN_575 & _GEN_576 & _GEN_1411))
      & (_GEN_566 | ~_GEN_563 | searcher_is_older_21 | ~(_GEN_564 & _GEN_565 & _GEN_1411))
      & (_GEN_555 | ~_GEN_552 | searcher_is_older_20 | ~(_GEN_553 & _GEN_554 & _GEN_1411))
      & (_GEN_544 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1411))
      & (_GEN_533 | ~_GEN_530 | searcher_is_older_18 | ~(_GEN_531 & _GEN_532 & _GEN_1411))
      & (_GEN_522 | ~_GEN_519 | searcher_is_older_17 | ~(_GEN_520 & _GEN_521 & _GEN_1411))
      & (_GEN_511 | ~_GEN_508 | searcher_is_older_16 | ~(_GEN_509 & _GEN_510 & _GEN_1411))
      & (_GEN_500 | ~_GEN_497 | searcher_is_older_15 | ~(_GEN_498 & _GEN_499 & _GEN_1411))
      & (_GEN_489 | ~_GEN_486 | searcher_is_older_14 | ~(_GEN_487 & _GEN_488 & _GEN_1411))
      & (_GEN_478 | ~_GEN_475 | searcher_is_older_13 | ~(_GEN_476 & _GEN_477 & _GEN_1411))
      & (_GEN_467 | ~_GEN_464 | searcher_is_older_12 | ~(_GEN_465 & _GEN_466 & _GEN_1411))
      & (_GEN_456 | ~_GEN_453 | searcher_is_older_11 | ~(_GEN_454 & _GEN_455 & _GEN_1411))
      & (_GEN_445 | ~_GEN_442 | searcher_is_older_10 | ~(_GEN_443 & _GEN_444 & _GEN_1411))
      & (_GEN_434 | ~_GEN_431 | searcher_is_older_9 | ~(_GEN_432 & _GEN_433 & _GEN_1411))
      & (_GEN_423 | ~_GEN_420 | searcher_is_older_8 | ~(_GEN_421 & _GEN_422 & _GEN_1411))
      & (_GEN_412 | ~_GEN_409 | searcher_is_older_7 | ~(_GEN_410 & _GEN_411 & _GEN_1411))
      & (_GEN_401 | ~_GEN_398 | searcher_is_older_6 | ~(_GEN_399 & _GEN_400 & _GEN_1411))
      & (_GEN_390 | ~_GEN_387 | searcher_is_older_5 | ~(_GEN_388 & _GEN_389 & _GEN_1411))
      & (_GEN_379 | ~_GEN_376 | searcher_is_older_4 | ~(_GEN_377 & _GEN_378 & _GEN_1411))
      & (_GEN_368 | ~_GEN_365 | searcher_is_older_3 | ~(_GEN_366 & _GEN_367 & _GEN_1411))
      & (_GEN_357 | ~_GEN_354 | searcher_is_older_2 | ~(_GEN_355 & _GEN_356 & _GEN_1411))
      & (_GEN_346 | ~_GEN_343 | searcher_is_older_1 | ~(_GEN_344 & _GEN_345 & _GEN_1411))
      & (_GEN_335 | ~_GEN_333 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_334 & _GEN_1411)) & s1_executing_loads_23;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    _GEN_1483 =
      _GEN_592
        ? (_GEN_1482
             ? (|lcam_ldq_idx_0) & _GEN_1458
             : ~(_GEN_596 & ~(|lcam_ldq_idx_0)) & _GEN_1458)
        : _GEN_1458;	// lsu.scala:1036:26, :1091:36, :1102:37, :1116:37, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1484 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1389 & _GEN_1459 : ~(_GEN_596 & _GEN_1389) & _GEN_1459)
        : _GEN_1459;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1485 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1390 & _GEN_1460 : ~(_GEN_596 & _GEN_1390) & _GEN_1460)
        : _GEN_1460;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1486 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1391 & _GEN_1461 : ~(_GEN_596 & _GEN_1391) & _GEN_1461)
        : _GEN_1461;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1487 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1392 & _GEN_1462 : ~(_GEN_596 & _GEN_1392) & _GEN_1462)
        : _GEN_1462;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1488 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1393 & _GEN_1463 : ~(_GEN_596 & _GEN_1393) & _GEN_1463)
        : _GEN_1463;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1489 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1394 & _GEN_1464 : ~(_GEN_596 & _GEN_1394) & _GEN_1464)
        : _GEN_1464;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1490 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1395 & _GEN_1465 : ~(_GEN_596 & _GEN_1395) & _GEN_1465)
        : _GEN_1465;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1491 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1396 & _GEN_1466 : ~(_GEN_596 & _GEN_1396) & _GEN_1466)
        : _GEN_1466;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1492 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1397 & _GEN_1467 : ~(_GEN_596 & _GEN_1397) & _GEN_1467)
        : _GEN_1467;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1493 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1398 & _GEN_1468 : ~(_GEN_596 & _GEN_1398) & _GEN_1468)
        : _GEN_1468;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1494 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1399 & _GEN_1469 : ~(_GEN_596 & _GEN_1399) & _GEN_1469)
        : _GEN_1469;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1495 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1400 & _GEN_1470 : ~(_GEN_596 & _GEN_1400) & _GEN_1470)
        : _GEN_1470;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1496 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1401 & _GEN_1471 : ~(_GEN_596 & _GEN_1401) & _GEN_1471)
        : _GEN_1471;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1497 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1402 & _GEN_1472 : ~(_GEN_596 & _GEN_1402) & _GEN_1472)
        : _GEN_1472;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1498 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1403 & _GEN_1473 : ~(_GEN_596 & _GEN_1403) & _GEN_1473)
        : _GEN_1473;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1499 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1404 & _GEN_1474 : ~(_GEN_596 & _GEN_1404) & _GEN_1474)
        : _GEN_1474;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1500 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1405 & _GEN_1475 : ~(_GEN_596 & _GEN_1405) & _GEN_1475)
        : _GEN_1475;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1501 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1406 & _GEN_1476 : ~(_GEN_596 & _GEN_1406) & _GEN_1476)
        : _GEN_1476;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1502 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1407 & _GEN_1477 : ~(_GEN_596 & _GEN_1407) & _GEN_1477)
        : _GEN_1477;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1503 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1408 & _GEN_1478 : ~(_GEN_596 & _GEN_1408) & _GEN_1478)
        : _GEN_1478;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1504 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1409 & _GEN_1479 : ~(_GEN_596 & _GEN_1409) & _GEN_1479)
        : _GEN_1479;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1505 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1410 & _GEN_1480 : ~(_GEN_596 & _GEN_1410) & _GEN_1480)
        : _GEN_1480;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1506 =
      _GEN_592
        ? (_GEN_1482 ? ~_GEN_1411 & _GEN_1481 : ~(_GEN_596 & _GEN_1411) & _GEN_1481)
        : _GEN_1481;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1508 =
      _GEN_599
        ? (_GEN_1507
             ? (|lcam_ldq_idx_0) & _GEN_1483
             : ~(_GEN_603 & ~(|lcam_ldq_idx_0)) & _GEN_1483)
        : _GEN_1483;	// lsu.scala:1036:26, :1091:36, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1509 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1389 & _GEN_1484 : ~(_GEN_603 & _GEN_1389) & _GEN_1484)
        : _GEN_1484;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1510 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1390 & _GEN_1485 : ~(_GEN_603 & _GEN_1390) & _GEN_1485)
        : _GEN_1485;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1511 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1391 & _GEN_1486 : ~(_GEN_603 & _GEN_1391) & _GEN_1486)
        : _GEN_1486;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1512 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1392 & _GEN_1487 : ~(_GEN_603 & _GEN_1392) & _GEN_1487)
        : _GEN_1487;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1513 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1393 & _GEN_1488 : ~(_GEN_603 & _GEN_1393) & _GEN_1488)
        : _GEN_1488;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1514 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1394 & _GEN_1489 : ~(_GEN_603 & _GEN_1394) & _GEN_1489)
        : _GEN_1489;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1515 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1395 & _GEN_1490 : ~(_GEN_603 & _GEN_1395) & _GEN_1490)
        : _GEN_1490;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1516 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1396 & _GEN_1491 : ~(_GEN_603 & _GEN_1396) & _GEN_1491)
        : _GEN_1491;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1517 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1397 & _GEN_1492 : ~(_GEN_603 & _GEN_1397) & _GEN_1492)
        : _GEN_1492;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1518 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1398 & _GEN_1493 : ~(_GEN_603 & _GEN_1398) & _GEN_1493)
        : _GEN_1493;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1519 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1399 & _GEN_1494 : ~(_GEN_603 & _GEN_1399) & _GEN_1494)
        : _GEN_1494;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1520 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1400 & _GEN_1495 : ~(_GEN_603 & _GEN_1400) & _GEN_1495)
        : _GEN_1495;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1521 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1401 & _GEN_1496 : ~(_GEN_603 & _GEN_1401) & _GEN_1496)
        : _GEN_1496;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1522 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1402 & _GEN_1497 : ~(_GEN_603 & _GEN_1402) & _GEN_1497)
        : _GEN_1497;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1523 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1403 & _GEN_1498 : ~(_GEN_603 & _GEN_1403) & _GEN_1498)
        : _GEN_1498;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1524 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1404 & _GEN_1499 : ~(_GEN_603 & _GEN_1404) & _GEN_1499)
        : _GEN_1499;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1525 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1405 & _GEN_1500 : ~(_GEN_603 & _GEN_1405) & _GEN_1500)
        : _GEN_1500;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1526 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1406 & _GEN_1501 : ~(_GEN_603 & _GEN_1406) & _GEN_1501)
        : _GEN_1501;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1527 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1407 & _GEN_1502 : ~(_GEN_603 & _GEN_1407) & _GEN_1502)
        : _GEN_1502;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1528 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1408 & _GEN_1503 : ~(_GEN_603 & _GEN_1408) & _GEN_1503)
        : _GEN_1503;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1529 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1409 & _GEN_1504 : ~(_GEN_603 & _GEN_1409) & _GEN_1504)
        : _GEN_1504;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1530 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1410 & _GEN_1505 : ~(_GEN_603 & _GEN_1410) & _GEN_1505)
        : _GEN_1505;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1531 =
      _GEN_599
        ? (_GEN_1507 ? ~_GEN_1411 & _GEN_1506 : ~(_GEN_603 & _GEN_1411) & _GEN_1506)
        : _GEN_1506;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1533 =
      _GEN_606
        ? (_GEN_1532
             ? (|lcam_ldq_idx_0) & _GEN_1508
             : ~(_GEN_610 & ~(|lcam_ldq_idx_0)) & _GEN_1508)
        : _GEN_1508;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1534 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1389 & _GEN_1509 : ~(_GEN_610 & _GEN_1389) & _GEN_1509)
        : _GEN_1509;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1535 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1390 & _GEN_1510 : ~(_GEN_610 & _GEN_1390) & _GEN_1510)
        : _GEN_1510;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1536 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1391 & _GEN_1511 : ~(_GEN_610 & _GEN_1391) & _GEN_1511)
        : _GEN_1511;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1537 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1392 & _GEN_1512 : ~(_GEN_610 & _GEN_1392) & _GEN_1512)
        : _GEN_1512;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1538 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1393 & _GEN_1513 : ~(_GEN_610 & _GEN_1393) & _GEN_1513)
        : _GEN_1513;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1539 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1394 & _GEN_1514 : ~(_GEN_610 & _GEN_1394) & _GEN_1514)
        : _GEN_1514;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1540 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1395 & _GEN_1515 : ~(_GEN_610 & _GEN_1395) & _GEN_1515)
        : _GEN_1515;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1541 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1396 & _GEN_1516 : ~(_GEN_610 & _GEN_1396) & _GEN_1516)
        : _GEN_1516;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1542 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1397 & _GEN_1517 : ~(_GEN_610 & _GEN_1397) & _GEN_1517)
        : _GEN_1517;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1543 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1398 & _GEN_1518 : ~(_GEN_610 & _GEN_1398) & _GEN_1518)
        : _GEN_1518;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1544 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1399 & _GEN_1519 : ~(_GEN_610 & _GEN_1399) & _GEN_1519)
        : _GEN_1519;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1545 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1400 & _GEN_1520 : ~(_GEN_610 & _GEN_1400) & _GEN_1520)
        : _GEN_1520;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1546 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1401 & _GEN_1521 : ~(_GEN_610 & _GEN_1401) & _GEN_1521)
        : _GEN_1521;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1547 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1402 & _GEN_1522 : ~(_GEN_610 & _GEN_1402) & _GEN_1522)
        : _GEN_1522;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1548 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1403 & _GEN_1523 : ~(_GEN_610 & _GEN_1403) & _GEN_1523)
        : _GEN_1523;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1549 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1404 & _GEN_1524 : ~(_GEN_610 & _GEN_1404) & _GEN_1524)
        : _GEN_1524;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1550 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1405 & _GEN_1525 : ~(_GEN_610 & _GEN_1405) & _GEN_1525)
        : _GEN_1525;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1551 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1406 & _GEN_1526 : ~(_GEN_610 & _GEN_1406) & _GEN_1526)
        : _GEN_1526;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1552 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1407 & _GEN_1527 : ~(_GEN_610 & _GEN_1407) & _GEN_1527)
        : _GEN_1527;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1553 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1408 & _GEN_1528 : ~(_GEN_610 & _GEN_1408) & _GEN_1528)
        : _GEN_1528;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1554 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1409 & _GEN_1529 : ~(_GEN_610 & _GEN_1409) & _GEN_1529)
        : _GEN_1529;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1555 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1410 & _GEN_1530 : ~(_GEN_610 & _GEN_1410) & _GEN_1530)
        : _GEN_1530;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1556 =
      _GEN_606
        ? (_GEN_1532 ? ~_GEN_1411 & _GEN_1531 : ~(_GEN_610 & _GEN_1411) & _GEN_1531)
        : _GEN_1531;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1558 =
      _GEN_613
        ? (_GEN_1557
             ? (|lcam_ldq_idx_0) & _GEN_1533
             : ~(_GEN_617 & ~(|lcam_ldq_idx_0)) & _GEN_1533)
        : _GEN_1533;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1559 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1389 & _GEN_1534 : ~(_GEN_617 & _GEN_1389) & _GEN_1534)
        : _GEN_1534;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1560 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1390 & _GEN_1535 : ~(_GEN_617 & _GEN_1390) & _GEN_1535)
        : _GEN_1535;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1561 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1391 & _GEN_1536 : ~(_GEN_617 & _GEN_1391) & _GEN_1536)
        : _GEN_1536;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1562 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1392 & _GEN_1537 : ~(_GEN_617 & _GEN_1392) & _GEN_1537)
        : _GEN_1537;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1563 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1393 & _GEN_1538 : ~(_GEN_617 & _GEN_1393) & _GEN_1538)
        : _GEN_1538;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1564 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1394 & _GEN_1539 : ~(_GEN_617 & _GEN_1394) & _GEN_1539)
        : _GEN_1539;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1565 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1395 & _GEN_1540 : ~(_GEN_617 & _GEN_1395) & _GEN_1540)
        : _GEN_1540;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1566 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1396 & _GEN_1541 : ~(_GEN_617 & _GEN_1396) & _GEN_1541)
        : _GEN_1541;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1567 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1397 & _GEN_1542 : ~(_GEN_617 & _GEN_1397) & _GEN_1542)
        : _GEN_1542;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1568 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1398 & _GEN_1543 : ~(_GEN_617 & _GEN_1398) & _GEN_1543)
        : _GEN_1543;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1569 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1399 & _GEN_1544 : ~(_GEN_617 & _GEN_1399) & _GEN_1544)
        : _GEN_1544;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1570 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1400 & _GEN_1545 : ~(_GEN_617 & _GEN_1400) & _GEN_1545)
        : _GEN_1545;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1571 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1401 & _GEN_1546 : ~(_GEN_617 & _GEN_1401) & _GEN_1546)
        : _GEN_1546;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1572 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1402 & _GEN_1547 : ~(_GEN_617 & _GEN_1402) & _GEN_1547)
        : _GEN_1547;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1573 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1403 & _GEN_1548 : ~(_GEN_617 & _GEN_1403) & _GEN_1548)
        : _GEN_1548;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1574 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1404 & _GEN_1549 : ~(_GEN_617 & _GEN_1404) & _GEN_1549)
        : _GEN_1549;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1575 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1405 & _GEN_1550 : ~(_GEN_617 & _GEN_1405) & _GEN_1550)
        : _GEN_1550;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1576 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1406 & _GEN_1551 : ~(_GEN_617 & _GEN_1406) & _GEN_1551)
        : _GEN_1551;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1577 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1407 & _GEN_1552 : ~(_GEN_617 & _GEN_1407) & _GEN_1552)
        : _GEN_1552;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1578 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1408 & _GEN_1553 : ~(_GEN_617 & _GEN_1408) & _GEN_1553)
        : _GEN_1553;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1579 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1409 & _GEN_1554 : ~(_GEN_617 & _GEN_1409) & _GEN_1554)
        : _GEN_1554;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1580 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1410 & _GEN_1555 : ~(_GEN_617 & _GEN_1410) & _GEN_1555)
        : _GEN_1555;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1581 =
      _GEN_613
        ? (_GEN_1557 ? ~_GEN_1411 & _GEN_1556 : ~(_GEN_617 & _GEN_1411) & _GEN_1556)
        : _GEN_1556;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1583 =
      _GEN_620
        ? (_GEN_1582
             ? (|lcam_ldq_idx_0) & _GEN_1558
             : ~(_GEN_624 & ~(|lcam_ldq_idx_0)) & _GEN_1558)
        : _GEN_1558;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1584 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1389 & _GEN_1559 : ~(_GEN_624 & _GEN_1389) & _GEN_1559)
        : _GEN_1559;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1585 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1390 & _GEN_1560 : ~(_GEN_624 & _GEN_1390) & _GEN_1560)
        : _GEN_1560;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1586 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1391 & _GEN_1561 : ~(_GEN_624 & _GEN_1391) & _GEN_1561)
        : _GEN_1561;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1587 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1392 & _GEN_1562 : ~(_GEN_624 & _GEN_1392) & _GEN_1562)
        : _GEN_1562;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1588 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1393 & _GEN_1563 : ~(_GEN_624 & _GEN_1393) & _GEN_1563)
        : _GEN_1563;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1589 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1394 & _GEN_1564 : ~(_GEN_624 & _GEN_1394) & _GEN_1564)
        : _GEN_1564;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1590 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1395 & _GEN_1565 : ~(_GEN_624 & _GEN_1395) & _GEN_1565)
        : _GEN_1565;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1591 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1396 & _GEN_1566 : ~(_GEN_624 & _GEN_1396) & _GEN_1566)
        : _GEN_1566;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1592 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1397 & _GEN_1567 : ~(_GEN_624 & _GEN_1397) & _GEN_1567)
        : _GEN_1567;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1593 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1398 & _GEN_1568 : ~(_GEN_624 & _GEN_1398) & _GEN_1568)
        : _GEN_1568;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1594 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1399 & _GEN_1569 : ~(_GEN_624 & _GEN_1399) & _GEN_1569)
        : _GEN_1569;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1595 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1400 & _GEN_1570 : ~(_GEN_624 & _GEN_1400) & _GEN_1570)
        : _GEN_1570;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1596 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1401 & _GEN_1571 : ~(_GEN_624 & _GEN_1401) & _GEN_1571)
        : _GEN_1571;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1597 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1402 & _GEN_1572 : ~(_GEN_624 & _GEN_1402) & _GEN_1572)
        : _GEN_1572;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1598 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1403 & _GEN_1573 : ~(_GEN_624 & _GEN_1403) & _GEN_1573)
        : _GEN_1573;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1599 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1404 & _GEN_1574 : ~(_GEN_624 & _GEN_1404) & _GEN_1574)
        : _GEN_1574;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1600 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1405 & _GEN_1575 : ~(_GEN_624 & _GEN_1405) & _GEN_1575)
        : _GEN_1575;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1601 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1406 & _GEN_1576 : ~(_GEN_624 & _GEN_1406) & _GEN_1576)
        : _GEN_1576;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1602 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1407 & _GEN_1577 : ~(_GEN_624 & _GEN_1407) & _GEN_1577)
        : _GEN_1577;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1603 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1408 & _GEN_1578 : ~(_GEN_624 & _GEN_1408) & _GEN_1578)
        : _GEN_1578;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1604 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1409 & _GEN_1579 : ~(_GEN_624 & _GEN_1409) & _GEN_1579)
        : _GEN_1579;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1605 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1410 & _GEN_1580 : ~(_GEN_624 & _GEN_1410) & _GEN_1580)
        : _GEN_1580;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1606 =
      _GEN_620
        ? (_GEN_1582 ? ~_GEN_1411 & _GEN_1581 : ~(_GEN_624 & _GEN_1411) & _GEN_1581)
        : _GEN_1581;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1608 =
      _GEN_627
        ? (_GEN_1607
             ? (|lcam_ldq_idx_0) & _GEN_1583
             : ~(_GEN_631 & ~(|lcam_ldq_idx_0)) & _GEN_1583)
        : _GEN_1583;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1609 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1389 & _GEN_1584 : ~(_GEN_631 & _GEN_1389) & _GEN_1584)
        : _GEN_1584;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1610 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1390 & _GEN_1585 : ~(_GEN_631 & _GEN_1390) & _GEN_1585)
        : _GEN_1585;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1611 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1391 & _GEN_1586 : ~(_GEN_631 & _GEN_1391) & _GEN_1586)
        : _GEN_1586;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1612 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1392 & _GEN_1587 : ~(_GEN_631 & _GEN_1392) & _GEN_1587)
        : _GEN_1587;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1613 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1393 & _GEN_1588 : ~(_GEN_631 & _GEN_1393) & _GEN_1588)
        : _GEN_1588;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1614 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1394 & _GEN_1589 : ~(_GEN_631 & _GEN_1394) & _GEN_1589)
        : _GEN_1589;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1615 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1395 & _GEN_1590 : ~(_GEN_631 & _GEN_1395) & _GEN_1590)
        : _GEN_1590;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1616 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1396 & _GEN_1591 : ~(_GEN_631 & _GEN_1396) & _GEN_1591)
        : _GEN_1591;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1617 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1397 & _GEN_1592 : ~(_GEN_631 & _GEN_1397) & _GEN_1592)
        : _GEN_1592;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1618 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1398 & _GEN_1593 : ~(_GEN_631 & _GEN_1398) & _GEN_1593)
        : _GEN_1593;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1619 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1399 & _GEN_1594 : ~(_GEN_631 & _GEN_1399) & _GEN_1594)
        : _GEN_1594;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1620 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1400 & _GEN_1595 : ~(_GEN_631 & _GEN_1400) & _GEN_1595)
        : _GEN_1595;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1621 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1401 & _GEN_1596 : ~(_GEN_631 & _GEN_1401) & _GEN_1596)
        : _GEN_1596;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1622 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1402 & _GEN_1597 : ~(_GEN_631 & _GEN_1402) & _GEN_1597)
        : _GEN_1597;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1623 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1403 & _GEN_1598 : ~(_GEN_631 & _GEN_1403) & _GEN_1598)
        : _GEN_1598;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1624 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1404 & _GEN_1599 : ~(_GEN_631 & _GEN_1404) & _GEN_1599)
        : _GEN_1599;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1625 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1405 & _GEN_1600 : ~(_GEN_631 & _GEN_1405) & _GEN_1600)
        : _GEN_1600;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1626 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1406 & _GEN_1601 : ~(_GEN_631 & _GEN_1406) & _GEN_1601)
        : _GEN_1601;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1627 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1407 & _GEN_1602 : ~(_GEN_631 & _GEN_1407) & _GEN_1602)
        : _GEN_1602;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1628 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1408 & _GEN_1603 : ~(_GEN_631 & _GEN_1408) & _GEN_1603)
        : _GEN_1603;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1629 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1409 & _GEN_1604 : ~(_GEN_631 & _GEN_1409) & _GEN_1604)
        : _GEN_1604;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1630 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1410 & _GEN_1605 : ~(_GEN_631 & _GEN_1410) & _GEN_1605)
        : _GEN_1605;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1631 =
      _GEN_627
        ? (_GEN_1607 ? ~_GEN_1411 & _GEN_1606 : ~(_GEN_631 & _GEN_1411) & _GEN_1606)
        : _GEN_1606;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1633 =
      _GEN_634
        ? (_GEN_1632
             ? (|lcam_ldq_idx_0) & _GEN_1608
             : ~(_GEN_638 & ~(|lcam_ldq_idx_0)) & _GEN_1608)
        : _GEN_1608;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1634 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1389 & _GEN_1609 : ~(_GEN_638 & _GEN_1389) & _GEN_1609)
        : _GEN_1609;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1635 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1390 & _GEN_1610 : ~(_GEN_638 & _GEN_1390) & _GEN_1610)
        : _GEN_1610;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1636 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1391 & _GEN_1611 : ~(_GEN_638 & _GEN_1391) & _GEN_1611)
        : _GEN_1611;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1637 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1392 & _GEN_1612 : ~(_GEN_638 & _GEN_1392) & _GEN_1612)
        : _GEN_1612;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1638 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1393 & _GEN_1613 : ~(_GEN_638 & _GEN_1393) & _GEN_1613)
        : _GEN_1613;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1639 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1394 & _GEN_1614 : ~(_GEN_638 & _GEN_1394) & _GEN_1614)
        : _GEN_1614;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1640 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1395 & _GEN_1615 : ~(_GEN_638 & _GEN_1395) & _GEN_1615)
        : _GEN_1615;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1641 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1396 & _GEN_1616 : ~(_GEN_638 & _GEN_1396) & _GEN_1616)
        : _GEN_1616;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1642 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1397 & _GEN_1617 : ~(_GEN_638 & _GEN_1397) & _GEN_1617)
        : _GEN_1617;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1643 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1398 & _GEN_1618 : ~(_GEN_638 & _GEN_1398) & _GEN_1618)
        : _GEN_1618;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1644 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1399 & _GEN_1619 : ~(_GEN_638 & _GEN_1399) & _GEN_1619)
        : _GEN_1619;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1645 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1400 & _GEN_1620 : ~(_GEN_638 & _GEN_1400) & _GEN_1620)
        : _GEN_1620;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1646 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1401 & _GEN_1621 : ~(_GEN_638 & _GEN_1401) & _GEN_1621)
        : _GEN_1621;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1647 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1402 & _GEN_1622 : ~(_GEN_638 & _GEN_1402) & _GEN_1622)
        : _GEN_1622;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1648 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1403 & _GEN_1623 : ~(_GEN_638 & _GEN_1403) & _GEN_1623)
        : _GEN_1623;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1649 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1404 & _GEN_1624 : ~(_GEN_638 & _GEN_1404) & _GEN_1624)
        : _GEN_1624;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1650 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1405 & _GEN_1625 : ~(_GEN_638 & _GEN_1405) & _GEN_1625)
        : _GEN_1625;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1651 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1406 & _GEN_1626 : ~(_GEN_638 & _GEN_1406) & _GEN_1626)
        : _GEN_1626;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1652 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1407 & _GEN_1627 : ~(_GEN_638 & _GEN_1407) & _GEN_1627)
        : _GEN_1627;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1653 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1408 & _GEN_1628 : ~(_GEN_638 & _GEN_1408) & _GEN_1628)
        : _GEN_1628;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1654 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1409 & _GEN_1629 : ~(_GEN_638 & _GEN_1409) & _GEN_1629)
        : _GEN_1629;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1655 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1410 & _GEN_1630 : ~(_GEN_638 & _GEN_1410) & _GEN_1630)
        : _GEN_1630;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1656 =
      _GEN_634
        ? (_GEN_1632 ? ~_GEN_1411 & _GEN_1631 : ~(_GEN_638 & _GEN_1411) & _GEN_1631)
        : _GEN_1631;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1658 =
      _GEN_641
        ? (_GEN_1657
             ? (|lcam_ldq_idx_0) & _GEN_1633
             : ~(_GEN_645 & ~(|lcam_ldq_idx_0)) & _GEN_1633)
        : _GEN_1633;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1659 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1389 & _GEN_1634 : ~(_GEN_645 & _GEN_1389) & _GEN_1634)
        : _GEN_1634;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1660 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1390 & _GEN_1635 : ~(_GEN_645 & _GEN_1390) & _GEN_1635)
        : _GEN_1635;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1661 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1391 & _GEN_1636 : ~(_GEN_645 & _GEN_1391) & _GEN_1636)
        : _GEN_1636;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1662 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1392 & _GEN_1637 : ~(_GEN_645 & _GEN_1392) & _GEN_1637)
        : _GEN_1637;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1663 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1393 & _GEN_1638 : ~(_GEN_645 & _GEN_1393) & _GEN_1638)
        : _GEN_1638;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1664 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1394 & _GEN_1639 : ~(_GEN_645 & _GEN_1394) & _GEN_1639)
        : _GEN_1639;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1665 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1395 & _GEN_1640 : ~(_GEN_645 & _GEN_1395) & _GEN_1640)
        : _GEN_1640;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1666 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1396 & _GEN_1641 : ~(_GEN_645 & _GEN_1396) & _GEN_1641)
        : _GEN_1641;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1667 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1397 & _GEN_1642 : ~(_GEN_645 & _GEN_1397) & _GEN_1642)
        : _GEN_1642;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1668 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1398 & _GEN_1643 : ~(_GEN_645 & _GEN_1398) & _GEN_1643)
        : _GEN_1643;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1669 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1399 & _GEN_1644 : ~(_GEN_645 & _GEN_1399) & _GEN_1644)
        : _GEN_1644;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1670 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1400 & _GEN_1645 : ~(_GEN_645 & _GEN_1400) & _GEN_1645)
        : _GEN_1645;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1671 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1401 & _GEN_1646 : ~(_GEN_645 & _GEN_1401) & _GEN_1646)
        : _GEN_1646;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1672 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1402 & _GEN_1647 : ~(_GEN_645 & _GEN_1402) & _GEN_1647)
        : _GEN_1647;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1673 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1403 & _GEN_1648 : ~(_GEN_645 & _GEN_1403) & _GEN_1648)
        : _GEN_1648;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1674 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1404 & _GEN_1649 : ~(_GEN_645 & _GEN_1404) & _GEN_1649)
        : _GEN_1649;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1675 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1405 & _GEN_1650 : ~(_GEN_645 & _GEN_1405) & _GEN_1650)
        : _GEN_1650;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1676 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1406 & _GEN_1651 : ~(_GEN_645 & _GEN_1406) & _GEN_1651)
        : _GEN_1651;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1677 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1407 & _GEN_1652 : ~(_GEN_645 & _GEN_1407) & _GEN_1652)
        : _GEN_1652;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1678 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1408 & _GEN_1653 : ~(_GEN_645 & _GEN_1408) & _GEN_1653)
        : _GEN_1653;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1679 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1409 & _GEN_1654 : ~(_GEN_645 & _GEN_1409) & _GEN_1654)
        : _GEN_1654;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1680 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1410 & _GEN_1655 : ~(_GEN_645 & _GEN_1410) & _GEN_1655)
        : _GEN_1655;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1681 =
      _GEN_641
        ? (_GEN_1657 ? ~_GEN_1411 & _GEN_1656 : ~(_GEN_645 & _GEN_1411) & _GEN_1656)
        : _GEN_1656;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1683 =
      _GEN_648
        ? (_GEN_1682
             ? (|lcam_ldq_idx_0) & _GEN_1658
             : ~(_GEN_652 & ~(|lcam_ldq_idx_0)) & _GEN_1658)
        : _GEN_1658;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1684 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1389 & _GEN_1659 : ~(_GEN_652 & _GEN_1389) & _GEN_1659)
        : _GEN_1659;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1685 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1390 & _GEN_1660 : ~(_GEN_652 & _GEN_1390) & _GEN_1660)
        : _GEN_1660;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1686 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1391 & _GEN_1661 : ~(_GEN_652 & _GEN_1391) & _GEN_1661)
        : _GEN_1661;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1687 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1392 & _GEN_1662 : ~(_GEN_652 & _GEN_1392) & _GEN_1662)
        : _GEN_1662;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1688 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1393 & _GEN_1663 : ~(_GEN_652 & _GEN_1393) & _GEN_1663)
        : _GEN_1663;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1689 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1394 & _GEN_1664 : ~(_GEN_652 & _GEN_1394) & _GEN_1664)
        : _GEN_1664;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1690 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1395 & _GEN_1665 : ~(_GEN_652 & _GEN_1395) & _GEN_1665)
        : _GEN_1665;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1691 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1396 & _GEN_1666 : ~(_GEN_652 & _GEN_1396) & _GEN_1666)
        : _GEN_1666;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1692 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1397 & _GEN_1667 : ~(_GEN_652 & _GEN_1397) & _GEN_1667)
        : _GEN_1667;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1693 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1398 & _GEN_1668 : ~(_GEN_652 & _GEN_1398) & _GEN_1668)
        : _GEN_1668;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1694 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1399 & _GEN_1669 : ~(_GEN_652 & _GEN_1399) & _GEN_1669)
        : _GEN_1669;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1695 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1400 & _GEN_1670 : ~(_GEN_652 & _GEN_1400) & _GEN_1670)
        : _GEN_1670;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1696 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1401 & _GEN_1671 : ~(_GEN_652 & _GEN_1401) & _GEN_1671)
        : _GEN_1671;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1697 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1402 & _GEN_1672 : ~(_GEN_652 & _GEN_1402) & _GEN_1672)
        : _GEN_1672;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1698 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1403 & _GEN_1673 : ~(_GEN_652 & _GEN_1403) & _GEN_1673)
        : _GEN_1673;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1699 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1404 & _GEN_1674 : ~(_GEN_652 & _GEN_1404) & _GEN_1674)
        : _GEN_1674;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1700 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1405 & _GEN_1675 : ~(_GEN_652 & _GEN_1405) & _GEN_1675)
        : _GEN_1675;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1701 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1406 & _GEN_1676 : ~(_GEN_652 & _GEN_1406) & _GEN_1676)
        : _GEN_1676;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1702 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1407 & _GEN_1677 : ~(_GEN_652 & _GEN_1407) & _GEN_1677)
        : _GEN_1677;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1703 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1408 & _GEN_1678 : ~(_GEN_652 & _GEN_1408) & _GEN_1678)
        : _GEN_1678;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1704 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1409 & _GEN_1679 : ~(_GEN_652 & _GEN_1409) & _GEN_1679)
        : _GEN_1679;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1705 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1410 & _GEN_1680 : ~(_GEN_652 & _GEN_1410) & _GEN_1680)
        : _GEN_1680;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1706 =
      _GEN_648
        ? (_GEN_1682 ? ~_GEN_1411 & _GEN_1681 : ~(_GEN_652 & _GEN_1411) & _GEN_1681)
        : _GEN_1681;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1708 =
      _GEN_655
        ? (_GEN_1707
             ? (|lcam_ldq_idx_0) & _GEN_1683
             : ~(_GEN_659 & ~(|lcam_ldq_idx_0)) & _GEN_1683)
        : _GEN_1683;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1709 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1389 & _GEN_1684 : ~(_GEN_659 & _GEN_1389) & _GEN_1684)
        : _GEN_1684;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1710 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1390 & _GEN_1685 : ~(_GEN_659 & _GEN_1390) & _GEN_1685)
        : _GEN_1685;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1711 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1391 & _GEN_1686 : ~(_GEN_659 & _GEN_1391) & _GEN_1686)
        : _GEN_1686;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1712 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1392 & _GEN_1687 : ~(_GEN_659 & _GEN_1392) & _GEN_1687)
        : _GEN_1687;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1713 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1393 & _GEN_1688 : ~(_GEN_659 & _GEN_1393) & _GEN_1688)
        : _GEN_1688;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1714 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1394 & _GEN_1689 : ~(_GEN_659 & _GEN_1394) & _GEN_1689)
        : _GEN_1689;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1715 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1395 & _GEN_1690 : ~(_GEN_659 & _GEN_1395) & _GEN_1690)
        : _GEN_1690;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1716 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1396 & _GEN_1691 : ~(_GEN_659 & _GEN_1396) & _GEN_1691)
        : _GEN_1691;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1717 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1397 & _GEN_1692 : ~(_GEN_659 & _GEN_1397) & _GEN_1692)
        : _GEN_1692;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1718 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1398 & _GEN_1693 : ~(_GEN_659 & _GEN_1398) & _GEN_1693)
        : _GEN_1693;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1719 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1399 & _GEN_1694 : ~(_GEN_659 & _GEN_1399) & _GEN_1694)
        : _GEN_1694;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1720 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1400 & _GEN_1695 : ~(_GEN_659 & _GEN_1400) & _GEN_1695)
        : _GEN_1695;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1721 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1401 & _GEN_1696 : ~(_GEN_659 & _GEN_1401) & _GEN_1696)
        : _GEN_1696;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1722 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1402 & _GEN_1697 : ~(_GEN_659 & _GEN_1402) & _GEN_1697)
        : _GEN_1697;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1723 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1403 & _GEN_1698 : ~(_GEN_659 & _GEN_1403) & _GEN_1698)
        : _GEN_1698;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1724 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1404 & _GEN_1699 : ~(_GEN_659 & _GEN_1404) & _GEN_1699)
        : _GEN_1699;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1725 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1405 & _GEN_1700 : ~(_GEN_659 & _GEN_1405) & _GEN_1700)
        : _GEN_1700;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1726 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1406 & _GEN_1701 : ~(_GEN_659 & _GEN_1406) & _GEN_1701)
        : _GEN_1701;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1727 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1407 & _GEN_1702 : ~(_GEN_659 & _GEN_1407) & _GEN_1702)
        : _GEN_1702;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1728 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1408 & _GEN_1703 : ~(_GEN_659 & _GEN_1408) & _GEN_1703)
        : _GEN_1703;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1729 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1409 & _GEN_1704 : ~(_GEN_659 & _GEN_1409) & _GEN_1704)
        : _GEN_1704;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1730 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1410 & _GEN_1705 : ~(_GEN_659 & _GEN_1410) & _GEN_1705)
        : _GEN_1705;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1731 =
      _GEN_655
        ? (_GEN_1707 ? ~_GEN_1411 & _GEN_1706 : ~(_GEN_659 & _GEN_1411) & _GEN_1706)
        : _GEN_1706;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1733 =
      _GEN_662
        ? (_GEN_1732
             ? (|lcam_ldq_idx_0) & _GEN_1708
             : ~(_GEN_666 & ~(|lcam_ldq_idx_0)) & _GEN_1708)
        : _GEN_1708;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1734 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1389 & _GEN_1709 : ~(_GEN_666 & _GEN_1389) & _GEN_1709)
        : _GEN_1709;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1735 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1390 & _GEN_1710 : ~(_GEN_666 & _GEN_1390) & _GEN_1710)
        : _GEN_1710;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1736 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1391 & _GEN_1711 : ~(_GEN_666 & _GEN_1391) & _GEN_1711)
        : _GEN_1711;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1737 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1392 & _GEN_1712 : ~(_GEN_666 & _GEN_1392) & _GEN_1712)
        : _GEN_1712;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1738 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1393 & _GEN_1713 : ~(_GEN_666 & _GEN_1393) & _GEN_1713)
        : _GEN_1713;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1739 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1394 & _GEN_1714 : ~(_GEN_666 & _GEN_1394) & _GEN_1714)
        : _GEN_1714;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1740 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1395 & _GEN_1715 : ~(_GEN_666 & _GEN_1395) & _GEN_1715)
        : _GEN_1715;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1741 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1396 & _GEN_1716 : ~(_GEN_666 & _GEN_1396) & _GEN_1716)
        : _GEN_1716;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1742 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1397 & _GEN_1717 : ~(_GEN_666 & _GEN_1397) & _GEN_1717)
        : _GEN_1717;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1743 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1398 & _GEN_1718 : ~(_GEN_666 & _GEN_1398) & _GEN_1718)
        : _GEN_1718;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1744 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1399 & _GEN_1719 : ~(_GEN_666 & _GEN_1399) & _GEN_1719)
        : _GEN_1719;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1745 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1400 & _GEN_1720 : ~(_GEN_666 & _GEN_1400) & _GEN_1720)
        : _GEN_1720;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1746 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1401 & _GEN_1721 : ~(_GEN_666 & _GEN_1401) & _GEN_1721)
        : _GEN_1721;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1747 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1402 & _GEN_1722 : ~(_GEN_666 & _GEN_1402) & _GEN_1722)
        : _GEN_1722;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1748 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1403 & _GEN_1723 : ~(_GEN_666 & _GEN_1403) & _GEN_1723)
        : _GEN_1723;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1749 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1404 & _GEN_1724 : ~(_GEN_666 & _GEN_1404) & _GEN_1724)
        : _GEN_1724;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1750 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1405 & _GEN_1725 : ~(_GEN_666 & _GEN_1405) & _GEN_1725)
        : _GEN_1725;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1751 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1406 & _GEN_1726 : ~(_GEN_666 & _GEN_1406) & _GEN_1726)
        : _GEN_1726;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1752 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1407 & _GEN_1727 : ~(_GEN_666 & _GEN_1407) & _GEN_1727)
        : _GEN_1727;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1753 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1408 & _GEN_1728 : ~(_GEN_666 & _GEN_1408) & _GEN_1728)
        : _GEN_1728;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1754 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1409 & _GEN_1729 : ~(_GEN_666 & _GEN_1409) & _GEN_1729)
        : _GEN_1729;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1755 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1410 & _GEN_1730 : ~(_GEN_666 & _GEN_1410) & _GEN_1730)
        : _GEN_1730;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1756 =
      _GEN_662
        ? (_GEN_1732 ? ~_GEN_1411 & _GEN_1731 : ~(_GEN_666 & _GEN_1411) & _GEN_1731)
        : _GEN_1731;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1758 =
      _GEN_669
        ? (_GEN_1757
             ? (|lcam_ldq_idx_0) & _GEN_1733
             : ~(_GEN_673 & ~(|lcam_ldq_idx_0)) & _GEN_1733)
        : _GEN_1733;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1759 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1389 & _GEN_1734 : ~(_GEN_673 & _GEN_1389) & _GEN_1734)
        : _GEN_1734;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1760 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1390 & _GEN_1735 : ~(_GEN_673 & _GEN_1390) & _GEN_1735)
        : _GEN_1735;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1761 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1391 & _GEN_1736 : ~(_GEN_673 & _GEN_1391) & _GEN_1736)
        : _GEN_1736;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1762 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1392 & _GEN_1737 : ~(_GEN_673 & _GEN_1392) & _GEN_1737)
        : _GEN_1737;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1763 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1393 & _GEN_1738 : ~(_GEN_673 & _GEN_1393) & _GEN_1738)
        : _GEN_1738;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1764 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1394 & _GEN_1739 : ~(_GEN_673 & _GEN_1394) & _GEN_1739)
        : _GEN_1739;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1765 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1395 & _GEN_1740 : ~(_GEN_673 & _GEN_1395) & _GEN_1740)
        : _GEN_1740;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1766 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1396 & _GEN_1741 : ~(_GEN_673 & _GEN_1396) & _GEN_1741)
        : _GEN_1741;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1767 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1397 & _GEN_1742 : ~(_GEN_673 & _GEN_1397) & _GEN_1742)
        : _GEN_1742;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1768 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1398 & _GEN_1743 : ~(_GEN_673 & _GEN_1398) & _GEN_1743)
        : _GEN_1743;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1769 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1399 & _GEN_1744 : ~(_GEN_673 & _GEN_1399) & _GEN_1744)
        : _GEN_1744;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1770 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1400 & _GEN_1745 : ~(_GEN_673 & _GEN_1400) & _GEN_1745)
        : _GEN_1745;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1771 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1401 & _GEN_1746 : ~(_GEN_673 & _GEN_1401) & _GEN_1746)
        : _GEN_1746;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1772 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1402 & _GEN_1747 : ~(_GEN_673 & _GEN_1402) & _GEN_1747)
        : _GEN_1747;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1773 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1403 & _GEN_1748 : ~(_GEN_673 & _GEN_1403) & _GEN_1748)
        : _GEN_1748;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1774 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1404 & _GEN_1749 : ~(_GEN_673 & _GEN_1404) & _GEN_1749)
        : _GEN_1749;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1775 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1405 & _GEN_1750 : ~(_GEN_673 & _GEN_1405) & _GEN_1750)
        : _GEN_1750;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1776 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1406 & _GEN_1751 : ~(_GEN_673 & _GEN_1406) & _GEN_1751)
        : _GEN_1751;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1777 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1407 & _GEN_1752 : ~(_GEN_673 & _GEN_1407) & _GEN_1752)
        : _GEN_1752;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1778 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1408 & _GEN_1753 : ~(_GEN_673 & _GEN_1408) & _GEN_1753)
        : _GEN_1753;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1779 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1409 & _GEN_1754 : ~(_GEN_673 & _GEN_1409) & _GEN_1754)
        : _GEN_1754;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1780 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1410 & _GEN_1755 : ~(_GEN_673 & _GEN_1410) & _GEN_1755)
        : _GEN_1755;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1781 =
      _GEN_669
        ? (_GEN_1757 ? ~_GEN_1411 & _GEN_1756 : ~(_GEN_673 & _GEN_1411) & _GEN_1756)
        : _GEN_1756;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1783 =
      _GEN_676
        ? (_GEN_1782
             ? (|lcam_ldq_idx_0) & _GEN_1758
             : ~(_GEN_680 & ~(|lcam_ldq_idx_0)) & _GEN_1758)
        : _GEN_1758;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1784 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1389 & _GEN_1759 : ~(_GEN_680 & _GEN_1389) & _GEN_1759)
        : _GEN_1759;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1785 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1390 & _GEN_1760 : ~(_GEN_680 & _GEN_1390) & _GEN_1760)
        : _GEN_1760;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1786 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1391 & _GEN_1761 : ~(_GEN_680 & _GEN_1391) & _GEN_1761)
        : _GEN_1761;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1787 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1392 & _GEN_1762 : ~(_GEN_680 & _GEN_1392) & _GEN_1762)
        : _GEN_1762;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1788 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1393 & _GEN_1763 : ~(_GEN_680 & _GEN_1393) & _GEN_1763)
        : _GEN_1763;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1789 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1394 & _GEN_1764 : ~(_GEN_680 & _GEN_1394) & _GEN_1764)
        : _GEN_1764;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1790 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1395 & _GEN_1765 : ~(_GEN_680 & _GEN_1395) & _GEN_1765)
        : _GEN_1765;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1791 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1396 & _GEN_1766 : ~(_GEN_680 & _GEN_1396) & _GEN_1766)
        : _GEN_1766;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1792 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1397 & _GEN_1767 : ~(_GEN_680 & _GEN_1397) & _GEN_1767)
        : _GEN_1767;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1793 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1398 & _GEN_1768 : ~(_GEN_680 & _GEN_1398) & _GEN_1768)
        : _GEN_1768;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1794 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1399 & _GEN_1769 : ~(_GEN_680 & _GEN_1399) & _GEN_1769)
        : _GEN_1769;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1795 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1400 & _GEN_1770 : ~(_GEN_680 & _GEN_1400) & _GEN_1770)
        : _GEN_1770;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1796 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1401 & _GEN_1771 : ~(_GEN_680 & _GEN_1401) & _GEN_1771)
        : _GEN_1771;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1797 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1402 & _GEN_1772 : ~(_GEN_680 & _GEN_1402) & _GEN_1772)
        : _GEN_1772;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1798 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1403 & _GEN_1773 : ~(_GEN_680 & _GEN_1403) & _GEN_1773)
        : _GEN_1773;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1799 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1404 & _GEN_1774 : ~(_GEN_680 & _GEN_1404) & _GEN_1774)
        : _GEN_1774;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1800 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1405 & _GEN_1775 : ~(_GEN_680 & _GEN_1405) & _GEN_1775)
        : _GEN_1775;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1801 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1406 & _GEN_1776 : ~(_GEN_680 & _GEN_1406) & _GEN_1776)
        : _GEN_1776;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1802 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1407 & _GEN_1777 : ~(_GEN_680 & _GEN_1407) & _GEN_1777)
        : _GEN_1777;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1803 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1408 & _GEN_1778 : ~(_GEN_680 & _GEN_1408) & _GEN_1778)
        : _GEN_1778;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1804 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1409 & _GEN_1779 : ~(_GEN_680 & _GEN_1409) & _GEN_1779)
        : _GEN_1779;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1805 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1410 & _GEN_1780 : ~(_GEN_680 & _GEN_1410) & _GEN_1780)
        : _GEN_1780;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1806 =
      _GEN_676
        ? (_GEN_1782 ? ~_GEN_1411 & _GEN_1781 : ~(_GEN_680 & _GEN_1411) & _GEN_1781)
        : _GEN_1781;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1808 =
      _GEN_683
        ? (_GEN_1807
             ? (|lcam_ldq_idx_0) & _GEN_1783
             : ~(_GEN_687 & ~(|lcam_ldq_idx_0)) & _GEN_1783)
        : _GEN_1783;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1809 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1389 & _GEN_1784 : ~(_GEN_687 & _GEN_1389) & _GEN_1784)
        : _GEN_1784;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1810 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1390 & _GEN_1785 : ~(_GEN_687 & _GEN_1390) & _GEN_1785)
        : _GEN_1785;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1811 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1391 & _GEN_1786 : ~(_GEN_687 & _GEN_1391) & _GEN_1786)
        : _GEN_1786;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1812 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1392 & _GEN_1787 : ~(_GEN_687 & _GEN_1392) & _GEN_1787)
        : _GEN_1787;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1813 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1393 & _GEN_1788 : ~(_GEN_687 & _GEN_1393) & _GEN_1788)
        : _GEN_1788;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1814 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1394 & _GEN_1789 : ~(_GEN_687 & _GEN_1394) & _GEN_1789)
        : _GEN_1789;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1815 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1395 & _GEN_1790 : ~(_GEN_687 & _GEN_1395) & _GEN_1790)
        : _GEN_1790;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1816 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1396 & _GEN_1791 : ~(_GEN_687 & _GEN_1396) & _GEN_1791)
        : _GEN_1791;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1817 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1397 & _GEN_1792 : ~(_GEN_687 & _GEN_1397) & _GEN_1792)
        : _GEN_1792;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1818 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1398 & _GEN_1793 : ~(_GEN_687 & _GEN_1398) & _GEN_1793)
        : _GEN_1793;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1819 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1399 & _GEN_1794 : ~(_GEN_687 & _GEN_1399) & _GEN_1794)
        : _GEN_1794;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1820 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1400 & _GEN_1795 : ~(_GEN_687 & _GEN_1400) & _GEN_1795)
        : _GEN_1795;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1821 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1401 & _GEN_1796 : ~(_GEN_687 & _GEN_1401) & _GEN_1796)
        : _GEN_1796;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1822 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1402 & _GEN_1797 : ~(_GEN_687 & _GEN_1402) & _GEN_1797)
        : _GEN_1797;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1823 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1403 & _GEN_1798 : ~(_GEN_687 & _GEN_1403) & _GEN_1798)
        : _GEN_1798;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1824 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1404 & _GEN_1799 : ~(_GEN_687 & _GEN_1404) & _GEN_1799)
        : _GEN_1799;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1825 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1405 & _GEN_1800 : ~(_GEN_687 & _GEN_1405) & _GEN_1800)
        : _GEN_1800;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1826 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1406 & _GEN_1801 : ~(_GEN_687 & _GEN_1406) & _GEN_1801)
        : _GEN_1801;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1827 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1407 & _GEN_1802 : ~(_GEN_687 & _GEN_1407) & _GEN_1802)
        : _GEN_1802;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1828 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1408 & _GEN_1803 : ~(_GEN_687 & _GEN_1408) & _GEN_1803)
        : _GEN_1803;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1829 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1409 & _GEN_1804 : ~(_GEN_687 & _GEN_1409) & _GEN_1804)
        : _GEN_1804;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1830 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1410 & _GEN_1805 : ~(_GEN_687 & _GEN_1410) & _GEN_1805)
        : _GEN_1805;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1831 =
      _GEN_683
        ? (_GEN_1807 ? ~_GEN_1411 & _GEN_1806 : ~(_GEN_687 & _GEN_1411) & _GEN_1806)
        : _GEN_1806;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1833 =
      _GEN_690
        ? (_GEN_1832
             ? (|lcam_ldq_idx_0) & _GEN_1808
             : ~(_GEN_694 & ~(|lcam_ldq_idx_0)) & _GEN_1808)
        : _GEN_1808;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1834 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1389 & _GEN_1809 : ~(_GEN_694 & _GEN_1389) & _GEN_1809)
        : _GEN_1809;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1835 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1390 & _GEN_1810 : ~(_GEN_694 & _GEN_1390) & _GEN_1810)
        : _GEN_1810;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1836 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1391 & _GEN_1811 : ~(_GEN_694 & _GEN_1391) & _GEN_1811)
        : _GEN_1811;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1837 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1392 & _GEN_1812 : ~(_GEN_694 & _GEN_1392) & _GEN_1812)
        : _GEN_1812;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1838 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1393 & _GEN_1813 : ~(_GEN_694 & _GEN_1393) & _GEN_1813)
        : _GEN_1813;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1839 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1394 & _GEN_1814 : ~(_GEN_694 & _GEN_1394) & _GEN_1814)
        : _GEN_1814;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1840 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1395 & _GEN_1815 : ~(_GEN_694 & _GEN_1395) & _GEN_1815)
        : _GEN_1815;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1841 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1396 & _GEN_1816 : ~(_GEN_694 & _GEN_1396) & _GEN_1816)
        : _GEN_1816;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1842 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1397 & _GEN_1817 : ~(_GEN_694 & _GEN_1397) & _GEN_1817)
        : _GEN_1817;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1843 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1398 & _GEN_1818 : ~(_GEN_694 & _GEN_1398) & _GEN_1818)
        : _GEN_1818;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1844 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1399 & _GEN_1819 : ~(_GEN_694 & _GEN_1399) & _GEN_1819)
        : _GEN_1819;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1845 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1400 & _GEN_1820 : ~(_GEN_694 & _GEN_1400) & _GEN_1820)
        : _GEN_1820;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1846 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1401 & _GEN_1821 : ~(_GEN_694 & _GEN_1401) & _GEN_1821)
        : _GEN_1821;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1847 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1402 & _GEN_1822 : ~(_GEN_694 & _GEN_1402) & _GEN_1822)
        : _GEN_1822;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1848 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1403 & _GEN_1823 : ~(_GEN_694 & _GEN_1403) & _GEN_1823)
        : _GEN_1823;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1849 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1404 & _GEN_1824 : ~(_GEN_694 & _GEN_1404) & _GEN_1824)
        : _GEN_1824;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1850 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1405 & _GEN_1825 : ~(_GEN_694 & _GEN_1405) & _GEN_1825)
        : _GEN_1825;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1851 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1406 & _GEN_1826 : ~(_GEN_694 & _GEN_1406) & _GEN_1826)
        : _GEN_1826;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1852 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1407 & _GEN_1827 : ~(_GEN_694 & _GEN_1407) & _GEN_1827)
        : _GEN_1827;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1853 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1408 & _GEN_1828 : ~(_GEN_694 & _GEN_1408) & _GEN_1828)
        : _GEN_1828;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1854 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1409 & _GEN_1829 : ~(_GEN_694 & _GEN_1409) & _GEN_1829)
        : _GEN_1829;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1855 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1410 & _GEN_1830 : ~(_GEN_694 & _GEN_1410) & _GEN_1830)
        : _GEN_1830;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1856 =
      _GEN_690
        ? (_GEN_1832 ? ~_GEN_1411 & _GEN_1831 : ~(_GEN_694 & _GEN_1411) & _GEN_1831)
        : _GEN_1831;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1858 =
      _GEN_697
        ? (_GEN_1857
             ? (|lcam_ldq_idx_0) & _GEN_1833
             : ~(_GEN_701 & ~(|lcam_ldq_idx_0)) & _GEN_1833)
        : _GEN_1833;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1859 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1389 & _GEN_1834 : ~(_GEN_701 & _GEN_1389) & _GEN_1834)
        : _GEN_1834;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1860 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1390 & _GEN_1835 : ~(_GEN_701 & _GEN_1390) & _GEN_1835)
        : _GEN_1835;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1861 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1391 & _GEN_1836 : ~(_GEN_701 & _GEN_1391) & _GEN_1836)
        : _GEN_1836;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1862 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1392 & _GEN_1837 : ~(_GEN_701 & _GEN_1392) & _GEN_1837)
        : _GEN_1837;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1863 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1393 & _GEN_1838 : ~(_GEN_701 & _GEN_1393) & _GEN_1838)
        : _GEN_1838;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1864 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1394 & _GEN_1839 : ~(_GEN_701 & _GEN_1394) & _GEN_1839)
        : _GEN_1839;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1865 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1395 & _GEN_1840 : ~(_GEN_701 & _GEN_1395) & _GEN_1840)
        : _GEN_1840;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1866 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1396 & _GEN_1841 : ~(_GEN_701 & _GEN_1396) & _GEN_1841)
        : _GEN_1841;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1867 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1397 & _GEN_1842 : ~(_GEN_701 & _GEN_1397) & _GEN_1842)
        : _GEN_1842;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1868 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1398 & _GEN_1843 : ~(_GEN_701 & _GEN_1398) & _GEN_1843)
        : _GEN_1843;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1869 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1399 & _GEN_1844 : ~(_GEN_701 & _GEN_1399) & _GEN_1844)
        : _GEN_1844;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1870 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1400 & _GEN_1845 : ~(_GEN_701 & _GEN_1400) & _GEN_1845)
        : _GEN_1845;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1871 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1401 & _GEN_1846 : ~(_GEN_701 & _GEN_1401) & _GEN_1846)
        : _GEN_1846;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1872 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1402 & _GEN_1847 : ~(_GEN_701 & _GEN_1402) & _GEN_1847)
        : _GEN_1847;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1873 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1403 & _GEN_1848 : ~(_GEN_701 & _GEN_1403) & _GEN_1848)
        : _GEN_1848;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1874 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1404 & _GEN_1849 : ~(_GEN_701 & _GEN_1404) & _GEN_1849)
        : _GEN_1849;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1875 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1405 & _GEN_1850 : ~(_GEN_701 & _GEN_1405) & _GEN_1850)
        : _GEN_1850;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1876 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1406 & _GEN_1851 : ~(_GEN_701 & _GEN_1406) & _GEN_1851)
        : _GEN_1851;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1877 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1407 & _GEN_1852 : ~(_GEN_701 & _GEN_1407) & _GEN_1852)
        : _GEN_1852;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1878 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1408 & _GEN_1853 : ~(_GEN_701 & _GEN_1408) & _GEN_1853)
        : _GEN_1853;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1879 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1409 & _GEN_1854 : ~(_GEN_701 & _GEN_1409) & _GEN_1854)
        : _GEN_1854;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1880 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1410 & _GEN_1855 : ~(_GEN_701 & _GEN_1410) & _GEN_1855)
        : _GEN_1855;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1881 =
      _GEN_697
        ? (_GEN_1857 ? ~_GEN_1411 & _GEN_1856 : ~(_GEN_701 & _GEN_1411) & _GEN_1856)
        : _GEN_1856;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1883 =
      _GEN_704
        ? (_GEN_1882
             ? (|lcam_ldq_idx_0) & _GEN_1858
             : ~(_GEN_708 & ~(|lcam_ldq_idx_0)) & _GEN_1858)
        : _GEN_1858;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1884 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1389 & _GEN_1859 : ~(_GEN_708 & _GEN_1389) & _GEN_1859)
        : _GEN_1859;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1885 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1390 & _GEN_1860 : ~(_GEN_708 & _GEN_1390) & _GEN_1860)
        : _GEN_1860;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1886 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1391 & _GEN_1861 : ~(_GEN_708 & _GEN_1391) & _GEN_1861)
        : _GEN_1861;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1887 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1392 & _GEN_1862 : ~(_GEN_708 & _GEN_1392) & _GEN_1862)
        : _GEN_1862;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1888 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1393 & _GEN_1863 : ~(_GEN_708 & _GEN_1393) & _GEN_1863)
        : _GEN_1863;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1889 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1394 & _GEN_1864 : ~(_GEN_708 & _GEN_1394) & _GEN_1864)
        : _GEN_1864;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1890 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1395 & _GEN_1865 : ~(_GEN_708 & _GEN_1395) & _GEN_1865)
        : _GEN_1865;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1891 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1396 & _GEN_1866 : ~(_GEN_708 & _GEN_1396) & _GEN_1866)
        : _GEN_1866;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1892 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1397 & _GEN_1867 : ~(_GEN_708 & _GEN_1397) & _GEN_1867)
        : _GEN_1867;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1893 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1398 & _GEN_1868 : ~(_GEN_708 & _GEN_1398) & _GEN_1868)
        : _GEN_1868;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1894 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1399 & _GEN_1869 : ~(_GEN_708 & _GEN_1399) & _GEN_1869)
        : _GEN_1869;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1895 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1400 & _GEN_1870 : ~(_GEN_708 & _GEN_1400) & _GEN_1870)
        : _GEN_1870;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1896 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1401 & _GEN_1871 : ~(_GEN_708 & _GEN_1401) & _GEN_1871)
        : _GEN_1871;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1897 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1402 & _GEN_1872 : ~(_GEN_708 & _GEN_1402) & _GEN_1872)
        : _GEN_1872;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1898 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1403 & _GEN_1873 : ~(_GEN_708 & _GEN_1403) & _GEN_1873)
        : _GEN_1873;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1899 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1404 & _GEN_1874 : ~(_GEN_708 & _GEN_1404) & _GEN_1874)
        : _GEN_1874;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1900 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1405 & _GEN_1875 : ~(_GEN_708 & _GEN_1405) & _GEN_1875)
        : _GEN_1875;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1901 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1406 & _GEN_1876 : ~(_GEN_708 & _GEN_1406) & _GEN_1876)
        : _GEN_1876;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1902 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1407 & _GEN_1877 : ~(_GEN_708 & _GEN_1407) & _GEN_1877)
        : _GEN_1877;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1903 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1408 & _GEN_1878 : ~(_GEN_708 & _GEN_1408) & _GEN_1878)
        : _GEN_1878;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1904 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1409 & _GEN_1879 : ~(_GEN_708 & _GEN_1409) & _GEN_1879)
        : _GEN_1879;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1905 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1410 & _GEN_1880 : ~(_GEN_708 & _GEN_1410) & _GEN_1880)
        : _GEN_1880;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1906 =
      _GEN_704
        ? (_GEN_1882 ? ~_GEN_1411 & _GEN_1881 : ~(_GEN_708 & _GEN_1411) & _GEN_1881)
        : _GEN_1881;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1908 =
      _GEN_711
        ? (_GEN_1907
             ? (|lcam_ldq_idx_0) & _GEN_1883
             : ~(_GEN_715 & ~(|lcam_ldq_idx_0)) & _GEN_1883)
        : _GEN_1883;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1909 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1389 & _GEN_1884 : ~(_GEN_715 & _GEN_1389) & _GEN_1884)
        : _GEN_1884;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1910 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1390 & _GEN_1885 : ~(_GEN_715 & _GEN_1390) & _GEN_1885)
        : _GEN_1885;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1911 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1391 & _GEN_1886 : ~(_GEN_715 & _GEN_1391) & _GEN_1886)
        : _GEN_1886;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1912 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1392 & _GEN_1887 : ~(_GEN_715 & _GEN_1392) & _GEN_1887)
        : _GEN_1887;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1913 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1393 & _GEN_1888 : ~(_GEN_715 & _GEN_1393) & _GEN_1888)
        : _GEN_1888;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1914 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1394 & _GEN_1889 : ~(_GEN_715 & _GEN_1394) & _GEN_1889)
        : _GEN_1889;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1915 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1395 & _GEN_1890 : ~(_GEN_715 & _GEN_1395) & _GEN_1890)
        : _GEN_1890;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1916 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1396 & _GEN_1891 : ~(_GEN_715 & _GEN_1396) & _GEN_1891)
        : _GEN_1891;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1917 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1397 & _GEN_1892 : ~(_GEN_715 & _GEN_1397) & _GEN_1892)
        : _GEN_1892;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1918 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1398 & _GEN_1893 : ~(_GEN_715 & _GEN_1398) & _GEN_1893)
        : _GEN_1893;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1919 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1399 & _GEN_1894 : ~(_GEN_715 & _GEN_1399) & _GEN_1894)
        : _GEN_1894;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1920 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1400 & _GEN_1895 : ~(_GEN_715 & _GEN_1400) & _GEN_1895)
        : _GEN_1895;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1921 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1401 & _GEN_1896 : ~(_GEN_715 & _GEN_1401) & _GEN_1896)
        : _GEN_1896;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1922 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1402 & _GEN_1897 : ~(_GEN_715 & _GEN_1402) & _GEN_1897)
        : _GEN_1897;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1923 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1403 & _GEN_1898 : ~(_GEN_715 & _GEN_1403) & _GEN_1898)
        : _GEN_1898;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1924 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1404 & _GEN_1899 : ~(_GEN_715 & _GEN_1404) & _GEN_1899)
        : _GEN_1899;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1925 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1405 & _GEN_1900 : ~(_GEN_715 & _GEN_1405) & _GEN_1900)
        : _GEN_1900;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1926 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1406 & _GEN_1901 : ~(_GEN_715 & _GEN_1406) & _GEN_1901)
        : _GEN_1901;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1927 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1407 & _GEN_1902 : ~(_GEN_715 & _GEN_1407) & _GEN_1902)
        : _GEN_1902;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1928 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1408 & _GEN_1903 : ~(_GEN_715 & _GEN_1408) & _GEN_1903)
        : _GEN_1903;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1929 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1409 & _GEN_1904 : ~(_GEN_715 & _GEN_1409) & _GEN_1904)
        : _GEN_1904;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1930 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1410 & _GEN_1905 : ~(_GEN_715 & _GEN_1410) & _GEN_1905)
        : _GEN_1905;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1931 =
      _GEN_711
        ? (_GEN_1907 ? ~_GEN_1411 & _GEN_1906 : ~(_GEN_715 & _GEN_1411) & _GEN_1906)
        : _GEN_1906;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1933 =
      _GEN_718
        ? (_GEN_1932
             ? (|lcam_ldq_idx_0) & _GEN_1908
             : ~(_GEN_722 & ~(|lcam_ldq_idx_0)) & _GEN_1908)
        : _GEN_1908;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1934 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1389 & _GEN_1909 : ~(_GEN_722 & _GEN_1389) & _GEN_1909)
        : _GEN_1909;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1935 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1390 & _GEN_1910 : ~(_GEN_722 & _GEN_1390) & _GEN_1910)
        : _GEN_1910;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1936 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1391 & _GEN_1911 : ~(_GEN_722 & _GEN_1391) & _GEN_1911)
        : _GEN_1911;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1937 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1392 & _GEN_1912 : ~(_GEN_722 & _GEN_1392) & _GEN_1912)
        : _GEN_1912;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1938 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1393 & _GEN_1913 : ~(_GEN_722 & _GEN_1393) & _GEN_1913)
        : _GEN_1913;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1939 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1394 & _GEN_1914 : ~(_GEN_722 & _GEN_1394) & _GEN_1914)
        : _GEN_1914;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1940 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1395 & _GEN_1915 : ~(_GEN_722 & _GEN_1395) & _GEN_1915)
        : _GEN_1915;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1941 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1396 & _GEN_1916 : ~(_GEN_722 & _GEN_1396) & _GEN_1916)
        : _GEN_1916;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1942 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1397 & _GEN_1917 : ~(_GEN_722 & _GEN_1397) & _GEN_1917)
        : _GEN_1917;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1943 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1398 & _GEN_1918 : ~(_GEN_722 & _GEN_1398) & _GEN_1918)
        : _GEN_1918;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1944 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1399 & _GEN_1919 : ~(_GEN_722 & _GEN_1399) & _GEN_1919)
        : _GEN_1919;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1945 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1400 & _GEN_1920 : ~(_GEN_722 & _GEN_1400) & _GEN_1920)
        : _GEN_1920;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1946 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1401 & _GEN_1921 : ~(_GEN_722 & _GEN_1401) & _GEN_1921)
        : _GEN_1921;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1947 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1402 & _GEN_1922 : ~(_GEN_722 & _GEN_1402) & _GEN_1922)
        : _GEN_1922;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1948 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1403 & _GEN_1923 : ~(_GEN_722 & _GEN_1403) & _GEN_1923)
        : _GEN_1923;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1949 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1404 & _GEN_1924 : ~(_GEN_722 & _GEN_1404) & _GEN_1924)
        : _GEN_1924;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1950 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1405 & _GEN_1925 : ~(_GEN_722 & _GEN_1405) & _GEN_1925)
        : _GEN_1925;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1951 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1406 & _GEN_1926 : ~(_GEN_722 & _GEN_1406) & _GEN_1926)
        : _GEN_1926;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1952 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1407 & _GEN_1927 : ~(_GEN_722 & _GEN_1407) & _GEN_1927)
        : _GEN_1927;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1953 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1408 & _GEN_1928 : ~(_GEN_722 & _GEN_1408) & _GEN_1928)
        : _GEN_1928;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1954 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1409 & _GEN_1929 : ~(_GEN_722 & _GEN_1409) & _GEN_1929)
        : _GEN_1929;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1955 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1410 & _GEN_1930 : ~(_GEN_722 & _GEN_1410) & _GEN_1930)
        : _GEN_1930;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1956 =
      _GEN_718
        ? (_GEN_1932 ? ~_GEN_1411 & _GEN_1931 : ~(_GEN_722 & _GEN_1411) & _GEN_1931)
        : _GEN_1931;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1958 =
      _GEN_725
        ? (_GEN_1957
             ? (|lcam_ldq_idx_0) & _GEN_1933
             : ~(_GEN_729 & ~(|lcam_ldq_idx_0)) & _GEN_1933)
        : _GEN_1933;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1959 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1389 & _GEN_1934 : ~(_GEN_729 & _GEN_1389) & _GEN_1934)
        : _GEN_1934;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1960 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1390 & _GEN_1935 : ~(_GEN_729 & _GEN_1390) & _GEN_1935)
        : _GEN_1935;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1961 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1391 & _GEN_1936 : ~(_GEN_729 & _GEN_1391) & _GEN_1936)
        : _GEN_1936;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1962 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1392 & _GEN_1937 : ~(_GEN_729 & _GEN_1392) & _GEN_1937)
        : _GEN_1937;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1963 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1393 & _GEN_1938 : ~(_GEN_729 & _GEN_1393) & _GEN_1938)
        : _GEN_1938;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1964 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1394 & _GEN_1939 : ~(_GEN_729 & _GEN_1394) & _GEN_1939)
        : _GEN_1939;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1965 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1395 & _GEN_1940 : ~(_GEN_729 & _GEN_1395) & _GEN_1940)
        : _GEN_1940;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1966 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1396 & _GEN_1941 : ~(_GEN_729 & _GEN_1396) & _GEN_1941)
        : _GEN_1941;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1967 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1397 & _GEN_1942 : ~(_GEN_729 & _GEN_1397) & _GEN_1942)
        : _GEN_1942;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1968 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1398 & _GEN_1943 : ~(_GEN_729 & _GEN_1398) & _GEN_1943)
        : _GEN_1943;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1969 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1399 & _GEN_1944 : ~(_GEN_729 & _GEN_1399) & _GEN_1944)
        : _GEN_1944;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1970 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1400 & _GEN_1945 : ~(_GEN_729 & _GEN_1400) & _GEN_1945)
        : _GEN_1945;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1971 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1401 & _GEN_1946 : ~(_GEN_729 & _GEN_1401) & _GEN_1946)
        : _GEN_1946;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1972 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1402 & _GEN_1947 : ~(_GEN_729 & _GEN_1402) & _GEN_1947)
        : _GEN_1947;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1973 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1403 & _GEN_1948 : ~(_GEN_729 & _GEN_1403) & _GEN_1948)
        : _GEN_1948;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1974 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1404 & _GEN_1949 : ~(_GEN_729 & _GEN_1404) & _GEN_1949)
        : _GEN_1949;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1975 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1405 & _GEN_1950 : ~(_GEN_729 & _GEN_1405) & _GEN_1950)
        : _GEN_1950;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1976 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1406 & _GEN_1951 : ~(_GEN_729 & _GEN_1406) & _GEN_1951)
        : _GEN_1951;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1977 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1407 & _GEN_1952 : ~(_GEN_729 & _GEN_1407) & _GEN_1952)
        : _GEN_1952;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1978 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1408 & _GEN_1953 : ~(_GEN_729 & _GEN_1408) & _GEN_1953)
        : _GEN_1953;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1979 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1409 & _GEN_1954 : ~(_GEN_729 & _GEN_1409) & _GEN_1954)
        : _GEN_1954;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1980 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1410 & _GEN_1955 : ~(_GEN_729 & _GEN_1410) & _GEN_1955)
        : _GEN_1955;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1981 =
      _GEN_725
        ? (_GEN_1957 ? ~_GEN_1411 & _GEN_1956 : ~(_GEN_729 & _GEN_1411) & _GEN_1956)
        : _GEN_1956;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1983 =
      _GEN_732
        ? (_GEN_1982
             ? (|lcam_ldq_idx_0) & _GEN_1958
             : ~(_GEN_736 & ~(|lcam_ldq_idx_0)) & _GEN_1958)
        : _GEN_1958;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1984 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1389 & _GEN_1959 : ~(_GEN_736 & _GEN_1389) & _GEN_1959)
        : _GEN_1959;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1985 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1390 & _GEN_1960 : ~(_GEN_736 & _GEN_1390) & _GEN_1960)
        : _GEN_1960;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1986 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1391 & _GEN_1961 : ~(_GEN_736 & _GEN_1391) & _GEN_1961)
        : _GEN_1961;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1987 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1392 & _GEN_1962 : ~(_GEN_736 & _GEN_1392) & _GEN_1962)
        : _GEN_1962;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1988 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1393 & _GEN_1963 : ~(_GEN_736 & _GEN_1393) & _GEN_1963)
        : _GEN_1963;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1989 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1394 & _GEN_1964 : ~(_GEN_736 & _GEN_1394) & _GEN_1964)
        : _GEN_1964;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1990 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1395 & _GEN_1965 : ~(_GEN_736 & _GEN_1395) & _GEN_1965)
        : _GEN_1965;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1991 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1396 & _GEN_1966 : ~(_GEN_736 & _GEN_1396) & _GEN_1966)
        : _GEN_1966;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1992 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1397 & _GEN_1967 : ~(_GEN_736 & _GEN_1397) & _GEN_1967)
        : _GEN_1967;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1993 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1398 & _GEN_1968 : ~(_GEN_736 & _GEN_1398) & _GEN_1968)
        : _GEN_1968;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1994 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1399 & _GEN_1969 : ~(_GEN_736 & _GEN_1399) & _GEN_1969)
        : _GEN_1969;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1995 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1400 & _GEN_1970 : ~(_GEN_736 & _GEN_1400) & _GEN_1970)
        : _GEN_1970;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1996 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1401 & _GEN_1971 : ~(_GEN_736 & _GEN_1401) & _GEN_1971)
        : _GEN_1971;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1997 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1402 & _GEN_1972 : ~(_GEN_736 & _GEN_1402) & _GEN_1972)
        : _GEN_1972;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1998 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1403 & _GEN_1973 : ~(_GEN_736 & _GEN_1403) & _GEN_1973)
        : _GEN_1973;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1999 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1404 & _GEN_1974 : ~(_GEN_736 & _GEN_1404) & _GEN_1974)
        : _GEN_1974;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2000 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1405 & _GEN_1975 : ~(_GEN_736 & _GEN_1405) & _GEN_1975)
        : _GEN_1975;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2001 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1406 & _GEN_1976 : ~(_GEN_736 & _GEN_1406) & _GEN_1976)
        : _GEN_1976;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2002 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1407 & _GEN_1977 : ~(_GEN_736 & _GEN_1407) & _GEN_1977)
        : _GEN_1977;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2003 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1408 & _GEN_1978 : ~(_GEN_736 & _GEN_1408) & _GEN_1978)
        : _GEN_1978;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2004 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1409 & _GEN_1979 : ~(_GEN_736 & _GEN_1409) & _GEN_1979)
        : _GEN_1979;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2005 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1410 & _GEN_1980 : ~(_GEN_736 & _GEN_1410) & _GEN_1980)
        : _GEN_1980;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2006 =
      _GEN_732
        ? (_GEN_1982 ? ~_GEN_1411 & _GEN_1981 : ~(_GEN_736 & _GEN_1411) & _GEN_1981)
        : _GEN_1981;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2008 =
      _GEN_739
        ? (_GEN_2007
             ? (|lcam_ldq_idx_0) & _GEN_1983
             : ~(_GEN_743 & ~(|lcam_ldq_idx_0)) & _GEN_1983)
        : _GEN_1983;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2009 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1389 & _GEN_1984 : ~(_GEN_743 & _GEN_1389) & _GEN_1984)
        : _GEN_1984;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2010 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1390 & _GEN_1985 : ~(_GEN_743 & _GEN_1390) & _GEN_1985)
        : _GEN_1985;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2011 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1391 & _GEN_1986 : ~(_GEN_743 & _GEN_1391) & _GEN_1986)
        : _GEN_1986;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2012 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1392 & _GEN_1987 : ~(_GEN_743 & _GEN_1392) & _GEN_1987)
        : _GEN_1987;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2013 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1393 & _GEN_1988 : ~(_GEN_743 & _GEN_1393) & _GEN_1988)
        : _GEN_1988;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2014 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1394 & _GEN_1989 : ~(_GEN_743 & _GEN_1394) & _GEN_1989)
        : _GEN_1989;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2015 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1395 & _GEN_1990 : ~(_GEN_743 & _GEN_1395) & _GEN_1990)
        : _GEN_1990;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2016 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1396 & _GEN_1991 : ~(_GEN_743 & _GEN_1396) & _GEN_1991)
        : _GEN_1991;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2017 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1397 & _GEN_1992 : ~(_GEN_743 & _GEN_1397) & _GEN_1992)
        : _GEN_1992;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2018 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1398 & _GEN_1993 : ~(_GEN_743 & _GEN_1398) & _GEN_1993)
        : _GEN_1993;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2019 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1399 & _GEN_1994 : ~(_GEN_743 & _GEN_1399) & _GEN_1994)
        : _GEN_1994;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2020 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1400 & _GEN_1995 : ~(_GEN_743 & _GEN_1400) & _GEN_1995)
        : _GEN_1995;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2021 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1401 & _GEN_1996 : ~(_GEN_743 & _GEN_1401) & _GEN_1996)
        : _GEN_1996;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2022 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1402 & _GEN_1997 : ~(_GEN_743 & _GEN_1402) & _GEN_1997)
        : _GEN_1997;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2023 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1403 & _GEN_1998 : ~(_GEN_743 & _GEN_1403) & _GEN_1998)
        : _GEN_1998;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2024 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1404 & _GEN_1999 : ~(_GEN_743 & _GEN_1404) & _GEN_1999)
        : _GEN_1999;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2025 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1405 & _GEN_2000 : ~(_GEN_743 & _GEN_1405) & _GEN_2000)
        : _GEN_2000;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2026 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1406 & _GEN_2001 : ~(_GEN_743 & _GEN_1406) & _GEN_2001)
        : _GEN_2001;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2027 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1407 & _GEN_2002 : ~(_GEN_743 & _GEN_1407) & _GEN_2002)
        : _GEN_2002;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2028 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1408 & _GEN_2003 : ~(_GEN_743 & _GEN_1408) & _GEN_2003)
        : _GEN_2003;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2029 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1409 & _GEN_2004 : ~(_GEN_743 & _GEN_1409) & _GEN_2004)
        : _GEN_2004;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2030 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1410 & _GEN_2005 : ~(_GEN_743 & _GEN_1410) & _GEN_2005)
        : _GEN_2005;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2031 =
      _GEN_739
        ? (_GEN_2007 ? ~_GEN_1411 & _GEN_2006 : ~(_GEN_743 & _GEN_1411) & _GEN_2006)
        : _GEN_2006;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2033 =
      _GEN_746
        ? (_GEN_2032
             ? (|lcam_ldq_idx_0) & _GEN_2008
             : ~(_GEN_750 & ~(|lcam_ldq_idx_0)) & _GEN_2008)
        : _GEN_2008;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2034 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1389 & _GEN_2009 : ~(_GEN_750 & _GEN_1389) & _GEN_2009)
        : _GEN_2009;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2035 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1390 & _GEN_2010 : ~(_GEN_750 & _GEN_1390) & _GEN_2010)
        : _GEN_2010;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2036 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1391 & _GEN_2011 : ~(_GEN_750 & _GEN_1391) & _GEN_2011)
        : _GEN_2011;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2037 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1392 & _GEN_2012 : ~(_GEN_750 & _GEN_1392) & _GEN_2012)
        : _GEN_2012;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2038 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1393 & _GEN_2013 : ~(_GEN_750 & _GEN_1393) & _GEN_2013)
        : _GEN_2013;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2039 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1394 & _GEN_2014 : ~(_GEN_750 & _GEN_1394) & _GEN_2014)
        : _GEN_2014;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2040 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1395 & _GEN_2015 : ~(_GEN_750 & _GEN_1395) & _GEN_2015)
        : _GEN_2015;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2041 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1396 & _GEN_2016 : ~(_GEN_750 & _GEN_1396) & _GEN_2016)
        : _GEN_2016;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2042 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1397 & _GEN_2017 : ~(_GEN_750 & _GEN_1397) & _GEN_2017)
        : _GEN_2017;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2043 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1398 & _GEN_2018 : ~(_GEN_750 & _GEN_1398) & _GEN_2018)
        : _GEN_2018;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2044 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1399 & _GEN_2019 : ~(_GEN_750 & _GEN_1399) & _GEN_2019)
        : _GEN_2019;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2045 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1400 & _GEN_2020 : ~(_GEN_750 & _GEN_1400) & _GEN_2020)
        : _GEN_2020;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2046 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1401 & _GEN_2021 : ~(_GEN_750 & _GEN_1401) & _GEN_2021)
        : _GEN_2021;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2047 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1402 & _GEN_2022 : ~(_GEN_750 & _GEN_1402) & _GEN_2022)
        : _GEN_2022;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2048 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1403 & _GEN_2023 : ~(_GEN_750 & _GEN_1403) & _GEN_2023)
        : _GEN_2023;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2049 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1404 & _GEN_2024 : ~(_GEN_750 & _GEN_1404) & _GEN_2024)
        : _GEN_2024;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2050 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1405 & _GEN_2025 : ~(_GEN_750 & _GEN_1405) & _GEN_2025)
        : _GEN_2025;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2051 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1406 & _GEN_2026 : ~(_GEN_750 & _GEN_1406) & _GEN_2026)
        : _GEN_2026;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2052 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1407 & _GEN_2027 : ~(_GEN_750 & _GEN_1407) & _GEN_2027)
        : _GEN_2027;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2053 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1408 & _GEN_2028 : ~(_GEN_750 & _GEN_1408) & _GEN_2028)
        : _GEN_2028;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2054 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1409 & _GEN_2029 : ~(_GEN_750 & _GEN_1409) & _GEN_2029)
        : _GEN_2029;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2055 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1410 & _GEN_2030 : ~(_GEN_750 & _GEN_1410) & _GEN_2030)
        : _GEN_2030;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_2056 =
      _GEN_746
        ? (_GEN_2032 ? ~_GEN_1411 & _GEN_2031 : ~(_GEN_750 & _GEN_1411) & _GEN_2031)
        : _GEN_2031;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    mem_forward_valid_0 =
      _GEN_2058[_forwarding_age_logic_0_io_forwarding_idx]
      & (io_core_brupdate_b1_mispredict_mask
         & (do_st_search_0
              ? (_lcam_stq_idx_T
                   ? mem_stq_incoming_e_0_bits_uop_br_mask
                   : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_br_mask : 16'h0)
              : do_ld_search_0
                  ? (fired_load_incoming_REG
                       ? mem_ldq_incoming_e_0_bits_uop_br_mask
                       : fired_load_retry_REG
                           ? mem_ldq_retry_e_bits_uop_br_mask
                           : fired_load_wakeup_REG
                               ? mem_ldq_wakeup_e_bits_uop_br_mask
                               : 16'h0)
                  : 16'h0)) == 16'h0 & ~io_core_exception & ~REG_1;	// lsu.scala:669:22, :894:51, :901:51, :902:51, :904:51, :909:37, :910:37, :911:37, :912:37, :913:37, :915:33, :916:33, :917:33, :919:{33,57}, :921:33, :1014:108, :1016:106, :1029:37, :1030:37, :1178:57, :1187:86, :1189:{53,56,64}, util.scala:118:{51,59}
    l_idx =
      _temp_bits_WIRE_1_24 & _temp_bits_T
        ? 6'h0
        : _temp_bits_WIRE_1_25 & _temp_bits_T_2
            ? 6'h1
            : _temp_bits_WIRE_1_26 & _temp_bits_T_4
                ? 6'h2
                : _temp_bits_WIRE_1_27 & _temp_bits_T_6
                    ? 6'h3
                    : _temp_bits_WIRE_1_28 & _temp_bits_T_8
                        ? 6'h4
                        : _temp_bits_WIRE_1_29 & _temp_bits_T_10
                            ? 6'h5
                            : _temp_bits_WIRE_1_30 & _temp_bits_T_12
                                ? 6'h6
                                : _temp_bits_WIRE_1_31 & _temp_bits_T_14
                                    ? 6'h7
                                    : _temp_bits_WIRE_1_32 & _temp_bits_T_16
                                        ? 6'h8
                                        : _temp_bits_WIRE_1_33 & _temp_bits_T_18
                                            ? 6'h9
                                            : _temp_bits_WIRE_1_34 & _temp_bits_T_20
                                                ? 6'hA
                                                : _temp_bits_WIRE_1_35 & _temp_bits_T_22
                                                    ? 6'hB
                                                    : _temp_bits_WIRE_1_36
                                                      & _temp_bits_T_24
                                                        ? 6'hC
                                                        : _temp_bits_WIRE_1_37
                                                          & _temp_bits_T_26
                                                            ? 6'hD
                                                            : _temp_bits_WIRE_1_38
                                                              & _temp_bits_T_28
                                                                ? 6'hE
                                                                : _temp_bits_WIRE_1_39
                                                                  & ~(ldq_head[4])
                                                                    ? 6'hF
                                                                    : _temp_bits_WIRE_1_40
                                                                      & _temp_bits_T_32
                                                                        ? 6'h10
                                                                        : _temp_bits_WIRE_1_41
                                                                          & _temp_bits_T_34
                                                                            ? 6'h11
                                                                            : _temp_bits_WIRE_1_42
                                                                              & _temp_bits_T_36
                                                                                ? 6'h12
                                                                                : _temp_bits_WIRE_1_43
                                                                                  & _temp_bits_T_38
                                                                                    ? 6'h13
                                                                                    : _temp_bits_WIRE_1_44
                                                                                      & _temp_bits_T_40
                                                                                        ? 6'h14
                                                                                        : _temp_bits_WIRE_1_45
                                                                                          & _temp_bits_T_42
                                                                                            ? 6'h15
                                                                                            : _temp_bits_WIRE_1_46
                                                                                              & _temp_bits_T_44
                                                                                                ? 6'h16
                                                                                                : _temp_bits_WIRE_1_47
                                                                                                  & _temp_bits_T_46
                                                                                                    ? 6'h17
                                                                                                    : _temp_bits_WIRE_1_24
                                                                                                        ? 6'h18
                                                                                                        : _temp_bits_WIRE_1_25
                                                                                                            ? 6'h19
                                                                                                            : _temp_bits_WIRE_1_26
                                                                                                                ? 6'h1A
                                                                                                                : _temp_bits_WIRE_1_27
                                                                                                                    ? 6'h1B
                                                                                                                    : _temp_bits_WIRE_1_28
                                                                                                                        ? 6'h1C
                                                                                                                        : _temp_bits_WIRE_1_29
                                                                                                                            ? 6'h1D
                                                                                                                            : _temp_bits_WIRE_1_30
                                                                                                                                ? 6'h1E
                                                                                                                                : _temp_bits_WIRE_1_31
                                                                                                                                    ? 6'h1F
                                                                                                                                    : _temp_bits_WIRE_1_32
                                                                                                                                        ? 6'h20
                                                                                                                                        : _temp_bits_WIRE_1_33
                                                                                                                                            ? 6'h21
                                                                                                                                            : _temp_bits_WIRE_1_34
                                                                                                                                                ? 6'h22
                                                                                                                                                : _temp_bits_WIRE_1_35
                                                                                                                                                    ? 6'h23
                                                                                                                                                    : _temp_bits_WIRE_1_36
                                                                                                                                                        ? 6'h24
                                                                                                                                                        : _temp_bits_WIRE_1_37
                                                                                                                                                            ? 6'h25
                                                                                                                                                            : _temp_bits_WIRE_1_38
                                                                                                                                                                ? 6'h26
                                                                                                                                                                : _temp_bits_WIRE_1_39
                                                                                                                                                                    ? 6'h27
                                                                                                                                                                    : _temp_bits_WIRE_1_40
                                                                                                                                                                        ? 6'h28
                                                                                                                                                                        : _temp_bits_WIRE_1_41
                                                                                                                                                                            ? 6'h29
                                                                                                                                                                            : _temp_bits_WIRE_1_42
                                                                                                                                                                                ? 6'h2A
                                                                                                                                                                                : _temp_bits_WIRE_1_43
                                                                                                                                                                                    ? 6'h2B
                                                                                                                                                                                    : _temp_bits_WIRE_1_44
                                                                                                                                                                                        ? 6'h2C
                                                                                                                                                                                        : _temp_bits_WIRE_1_45
                                                                                                                                                                                            ? 6'h2D
                                                                                                                                                                                            : {5'h17,
                                                                                                                                                                                               ~_temp_bits_WIRE_1_46};	// Mux.scala:47:69, lsu.scala:215:29, :1091:36, :1102:37, :1229:21, util.scala:205:25, :351:72
    ld_xcpt_valid =
      _temp_bits_WIRE_1_24 | _temp_bits_WIRE_1_25 | _temp_bits_WIRE_1_26
      | _temp_bits_WIRE_1_27 | _temp_bits_WIRE_1_28 | _temp_bits_WIRE_1_29
      | _temp_bits_WIRE_1_30 | _temp_bits_WIRE_1_31 | _temp_bits_WIRE_1_32
      | _temp_bits_WIRE_1_33 | _temp_bits_WIRE_1_34 | _temp_bits_WIRE_1_35
      | _temp_bits_WIRE_1_36 | _temp_bits_WIRE_1_37 | _temp_bits_WIRE_1_38
      | _temp_bits_WIRE_1_39 | _temp_bits_WIRE_1_40 | _temp_bits_WIRE_1_41
      | _temp_bits_WIRE_1_42 | _temp_bits_WIRE_1_43 | _temp_bits_WIRE_1_44
      | _temp_bits_WIRE_1_45 | _temp_bits_WIRE_1_46 | _temp_bits_WIRE_1_47;	// lsu.scala:1091:36, :1102:37, :1238:44
    _ld_xcpt_uop_T_3 = l_idx > 6'h17 ? l_idx[4:0] + 5'h8 : l_idx[4:0];	// Mux.scala:47:69, lsu.scala:305:44, :1239:{30,37,63}
    use_mem_xcpt =
      mem_xcpt_valids_0
      & (mem_xcpt_uops_0_rob_idx < _GEN_148[_ld_xcpt_uop_T_3]
         ^ mem_xcpt_uops_0_rob_idx < io_core_rob_head_idx
         ^ _GEN_148[_ld_xcpt_uop_T_3] < io_core_rob_head_idx) | ~ld_xcpt_valid;	// lsu.scala:465:79, :667:32, :671:32, :1238:44, :1239:30, :1241:{38,115,118}, util.scala:363:{52,64,72,78}
    xcpt_uop_br_mask =
      use_mem_xcpt ? mem_xcpt_uops_0_br_mask : _GEN_110[_ld_xcpt_uop_T_3];	// lsu.scala:264:49, :671:32, :1239:30, :1241:115, :1243:21, util.scala:363:52
    _GEN_2060 = _GEN_788 & _GEN_2059 & ~(|wb_forward_ldq_idx_0);	// lsu.scala:1065:36, :1075:88, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2061 = _GEN_787 | ~_GEN_2060;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2062 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h1;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2063 = _GEN_787 | ~_GEN_2062;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2064 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h2;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2065 = _GEN_787 | ~_GEN_2064;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2066 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h3;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2067 = _GEN_787 | ~_GEN_2066;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2068 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h4;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2069 = _GEN_787 | ~_GEN_2068;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2070 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h5;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2071 = _GEN_787 | ~_GEN_2070;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2072 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h6;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2073 = _GEN_787 | ~_GEN_2072;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2074 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h7;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2075 = _GEN_787 | ~_GEN_2074;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2076 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h8;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2077 = _GEN_787 | ~_GEN_2076;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2078 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h9;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2079 = _GEN_787 | ~_GEN_2078;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2080 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'hA;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2081 = _GEN_787 | ~_GEN_2080;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2082 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'hB;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2083 = _GEN_787 | ~_GEN_2082;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2084 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'hC;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2085 = _GEN_787 | ~_GEN_2084;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2086 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'hD;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2087 = _GEN_787 | ~_GEN_2086;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2088 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'hE;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2089 = _GEN_787 | ~_GEN_2088;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2090 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'hF;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2091 = _GEN_787 | ~_GEN_2090;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2092 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h10;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2093 = _GEN_787 | ~_GEN_2092;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2094 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h11;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2095 = _GEN_787 | ~_GEN_2094;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2096 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h12;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2097 = _GEN_787 | ~_GEN_2096;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2098 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h13;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2099 = _GEN_787 | ~_GEN_2098;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2100 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h14;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2101 = _GEN_787 | ~_GEN_2100;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2102 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h15;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2103 = _GEN_787 | ~_GEN_2102;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2104 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h16;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_2105 = _GEN_787 | ~_GEN_2104;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2106 = _GEN_788 & _GEN_2059 & wb_forward_ldq_idx_0 == 5'h17;	// lsu.scala:1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35, util.scala:205:25
    _GEN_2107 = _GEN_787 | ~_GEN_2106;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_2108 = stq_0_valid & (|_GEN_802);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2109 = stq_1_valid & (|_GEN_803);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2110 = stq_2_valid & (|_GEN_804);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2111 = stq_3_valid & (|_GEN_805);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2112 = stq_4_valid & (|_GEN_806);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2113 = stq_5_valid & (|_GEN_807);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2114 = stq_6_valid & (|_GEN_808);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2115 = stq_7_valid & (|_GEN_809);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2116 = stq_8_valid & (|_GEN_810);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2117 = stq_9_valid & (|_GEN_811);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2118 = stq_10_valid & (|_GEN_812);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2119 = stq_11_valid & (|_GEN_813);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2120 = stq_12_valid & (|_GEN_814);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2121 = stq_13_valid & (|_GEN_815);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2122 = stq_14_valid & (|_GEN_816);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2123 = stq_15_valid & (|_GEN_817);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2124 = stq_16_valid & (|_GEN_818);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2125 = stq_17_valid & (|_GEN_819);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2126 = stq_18_valid & (|_GEN_820);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2127 = stq_19_valid & (|_GEN_821);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2128 = stq_20_valid & (|_GEN_822);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2129 = stq_21_valid & (|_GEN_823);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2130 = stq_22_valid & (|_GEN_824);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2131 = stq_23_valid & (|_GEN_825);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_2132 =
      ldq_0_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_0_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2133 =
      ldq_1_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_1_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2134 =
      ldq_2_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_2_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2135 =
      ldq_3_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_3_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2136 =
      ldq_4_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_4_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2137 =
      ldq_5_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_5_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2138 =
      ldq_6_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_6_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2139 =
      ldq_7_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_7_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2140 =
      ldq_8_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_8_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2141 =
      ldq_9_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_9_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2142 =
      ldq_10_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_10_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2143 =
      ldq_11_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_11_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2144 =
      ldq_12_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_12_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2145 =
      ldq_13_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_13_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2146 =
      ldq_14_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_14_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2147 =
      ldq_15_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_15_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2148 =
      ldq_16_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_16_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2149 =
      ldq_17_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_17_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2150 =
      ldq_18_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_18_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2151 =
      ldq_19_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_19_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2152 =
      ldq_20_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_20_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2153 =
      ldq_21_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_21_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2154 =
      ldq_22_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_22_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2155 =
      ldq_23_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_23_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_2204 = _GEN_2156 | _GEN_2132;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2206 = _GEN_2158 | _GEN_2133;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2207 = _GEN_2160 | _GEN_2134;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2208 = _GEN_2162 | _GEN_2135;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2209 = _GEN_2164 | _GEN_2136;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2210 = _GEN_2166 | _GEN_2137;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2211 = _GEN_2168 | _GEN_2138;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2212 = _GEN_2170 | _GEN_2139;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2213 = _GEN_2172 | _GEN_2140;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2214 = _GEN_2174 | _GEN_2141;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2215 = _GEN_2176 | _GEN_2142;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2216 = _GEN_2178 | _GEN_2143;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2217 = _GEN_2180 | _GEN_2144;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2218 = _GEN_2182 | _GEN_2145;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2219 = _GEN_2184 | _GEN_2146;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2220 = _GEN_2186 | _GEN_2147;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2221 = _GEN_2188 | _GEN_2148;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2222 = _GEN_2190 | _GEN_2149;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2223 = _GEN_2192 | _GEN_2150;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2224 = _GEN_2194 | _GEN_2151;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2225 = _GEN_2196 | _GEN_2152;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2226 = _GEN_2198 | _GEN_2153;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2227 = _GEN_2200 | _GEN_2154;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2228 = _GEN_2202 | _GEN_2155;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_2349 = stq_head == 5'h0;	// lsu.scala:217:29, :1506:35
    _GEN_2350 = _GEN_2349 | _GEN_2108;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2351 = stq_head == 5'h1;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2352 = _GEN_2351 | _GEN_2109;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2353 = stq_head == 5'h2;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2354 = _GEN_2353 | _GEN_2110;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2355 = stq_head == 5'h3;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2356 = _GEN_2355 | _GEN_2111;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2357 = stq_head == 5'h4;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2358 = _GEN_2357 | _GEN_2112;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2359 = stq_head == 5'h5;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2360 = _GEN_2359 | _GEN_2113;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2361 = stq_head == 5'h6;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2362 = _GEN_2361 | _GEN_2114;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2363 = stq_head == 5'h7;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2364 = _GEN_2363 | _GEN_2115;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2365 = stq_head == 5'h8;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2366 = _GEN_2365 | _GEN_2116;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2367 = stq_head == 5'h9;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2368 = _GEN_2367 | _GEN_2117;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2369 = stq_head == 5'hA;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2370 = _GEN_2369 | _GEN_2118;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2371 = stq_head == 5'hB;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2372 = _GEN_2371 | _GEN_2119;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2373 = stq_head == 5'hC;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2374 = _GEN_2373 | _GEN_2120;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2375 = stq_head == 5'hD;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2376 = _GEN_2375 | _GEN_2121;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2377 = stq_head == 5'hE;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2378 = _GEN_2377 | _GEN_2122;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2379 = stq_head == 5'hF;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2380 = _GEN_2379 | _GEN_2123;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2381 = stq_head == 5'h10;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2382 = _GEN_2381 | _GEN_2124;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2383 = stq_head == 5'h11;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2384 = _GEN_2383 | _GEN_2125;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2385 = stq_head == 5'h12;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2386 = _GEN_2385 | _GEN_2126;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2387 = stq_head == 5'h13;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2388 = _GEN_2387 | _GEN_2127;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2389 = stq_head == 5'h14;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2390 = _GEN_2389 | _GEN_2128;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2391 = stq_head == 5'h15;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2392 = _GEN_2391 | _GEN_2129;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2393 = stq_head == 5'h16;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_2394 = _GEN_2393 | _GEN_2130;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2395 = stq_head == 5'h17;	// lsu.scala:217:29, :1506:35, util.scala:205:25
    _GEN_2396 = _GEN_2395 | _GEN_2131;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_2397 = clear_store & _GEN_2349;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2398 = clear_store & _GEN_2351;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2399 = clear_store & _GEN_2353;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2400 = clear_store & _GEN_2355;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2401 = clear_store & _GEN_2357;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2402 = clear_store & _GEN_2359;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2403 = clear_store & _GEN_2361;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2404 = clear_store & _GEN_2363;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2405 = clear_store & _GEN_2365;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2406 = clear_store & _GEN_2367;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2407 = clear_store & _GEN_2369;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2408 = clear_store & _GEN_2371;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2409 = clear_store & _GEN_2373;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2410 = clear_store & _GEN_2375;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2411 = clear_store & _GEN_2377;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2412 = clear_store & _GEN_2379;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2413 = clear_store & _GEN_2381;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2414 = clear_store & _GEN_2383;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2415 = clear_store & _GEN_2385;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2416 = clear_store & _GEN_2387;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2417 = clear_store & _GEN_2389;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2418 = clear_store & _GEN_2391;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2419 = clear_store & _GEN_2393;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2420 = clear_store & _GEN_2395;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_2421 = ~(|hella_state) & io_hellacache_req_valid;	// Decoupled.scala:40:37, lsu.scala:242:38, :593:24, :1527:21
    _GEN_2422 = ~(|hella_state) & _GEN_2421;	// Decoupled.scala:40:37, lsu.scala:242:38, :243:34, :593:24, :1527:{21,34}, :1529:37, :1530:19
    _GEN_2423 = (|hella_state) & _GEN_1;	// lsu.scala:242:38, :244:34, :593:24, :803:26, :1527:34, :1533:38
    _GEN_2424 = reset | io_core_exception;	// lsu.scala:1596:22
    _GEN_2425 = _GEN_2424 & reset;	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1603:16
    _GEN_2426 = ~stq_0_bits_committed & ~stq_0_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2427 = _GEN_2424 & (reset | _GEN_2426);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2428 = ~stq_1_bits_committed & ~stq_1_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2429 = _GEN_2424 & (reset | _GEN_2428);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2430 = ~stq_2_bits_committed & ~stq_2_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2431 = _GEN_2424 & (reset | _GEN_2430);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2432 = ~stq_3_bits_committed & ~stq_3_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2433 = _GEN_2424 & (reset | _GEN_2432);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2434 = ~stq_4_bits_committed & ~stq_4_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2435 = _GEN_2424 & (reset | _GEN_2434);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2436 = ~stq_5_bits_committed & ~stq_5_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2437 = _GEN_2424 & (reset | _GEN_2436);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2438 = ~stq_6_bits_committed & ~stq_6_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2439 = _GEN_2424 & (reset | _GEN_2438);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2440 = ~stq_7_bits_committed & ~stq_7_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2441 = _GEN_2424 & (reset | _GEN_2440);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2442 = ~stq_8_bits_committed & ~stq_8_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2443 = _GEN_2424 & (reset | _GEN_2442);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2444 = ~stq_9_bits_committed & ~stq_9_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2445 = _GEN_2424 & (reset | _GEN_2444);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2446 = ~stq_10_bits_committed & ~stq_10_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2447 = _GEN_2424 & (reset | _GEN_2446);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2448 = ~stq_11_bits_committed & ~stq_11_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2449 = _GEN_2424 & (reset | _GEN_2448);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2450 = ~stq_12_bits_committed & ~stq_12_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2451 = _GEN_2424 & (reset | _GEN_2450);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2452 = ~stq_13_bits_committed & ~stq_13_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2453 = _GEN_2424 & (reset | _GEN_2452);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2454 = ~stq_14_bits_committed & ~stq_14_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2455 = _GEN_2424 & (reset | _GEN_2454);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2456 = ~stq_15_bits_committed & ~stq_15_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2457 = _GEN_2424 & (reset | _GEN_2456);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2458 = ~stq_16_bits_committed & ~stq_16_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2459 = _GEN_2424 & (reset | _GEN_2458);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2460 = ~stq_17_bits_committed & ~stq_17_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2461 = _GEN_2424 & (reset | _GEN_2460);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2462 = ~stq_18_bits_committed & ~stq_18_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2463 = _GEN_2424 & (reset | _GEN_2462);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2464 = ~stq_19_bits_committed & ~stq_19_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2465 = _GEN_2424 & (reset | _GEN_2464);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2466 = ~stq_20_bits_committed & ~stq_20_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2467 = _GEN_2424 & (reset | _GEN_2466);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2468 = ~stq_21_bits_committed & ~stq_21_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2469 = _GEN_2424 & (reset | _GEN_2468);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2470 = ~stq_22_bits_committed & ~stq_22_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2471 = _GEN_2424 & (reset | _GEN_2470);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_2472 = ~stq_23_bits_committed & ~stq_23_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_2473 = _GEN_2424 & (reset | _GEN_2472);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    ldq_0_valid <=
      ~_GEN_2424 & _GEN_2325 & _GEN_2277
      & (_GEN_2205 ? ~_GEN_2132 & _GEN_1052 : ~_GEN_2204 & _GEN_1052);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1051) begin	// lsu.scala:304:5, :305:44
      ldq_0_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_0_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_0_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_0_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_0_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_0_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_0_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_0_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_0_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_977) begin	// lsu.scala:304:5, :306:44
      ldq_0_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_0_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_0_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_0_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_0_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_0_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_0_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_855) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_0_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_0_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_0_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_0_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_0_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_0_valid)	// lsu.scala:210:16
      ldq_0_bits_uop_br_mask <=
        ldq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1051)	// lsu.scala:304:5, :305:44
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_977)	// lsu.scala:304:5, :306:44
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_855)	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1243) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_0_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_0_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_0_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_0_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_0_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_0_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_0_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_0_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_0_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_0_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_0_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1051)	// lsu.scala:304:5, :305:44
      ldq_0_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_977)	// lsu.scala:304:5, :306:44
      ldq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_855)	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1099)	// lsu.scala:210:16, :304:5, :306:44
      ldq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_0_bits_uop_ppred_busy <= ~_GEN_1099 & ldq_0_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_0_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h0
      | (_GEN_1051
           ? io_core_dis_uops_2_bits_exception
           : _GEN_977
               ? io_core_dis_uops_1_bits_exception
               : _GEN_855 ? io_core_dis_uops_0_bits_exception : ldq_0_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_0_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2325 & _GEN_2277
      & (_GEN_2205 ? ~_GEN_2132 & _GEN_1244 : ~_GEN_2204 & _GEN_1244);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_0_bits_executed <=
      ~_GEN_2424 & _GEN_2325 & _GEN_2277 & _GEN_2229
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_761))
      & ((_GEN_753
            ? (_GEN_2057
                 ? (|lcam_ldq_idx_0) & _GEN_2033
                 : ~(_GEN_757 & ~(|lcam_ldq_idx_0)) & _GEN_2033)
            : _GEN_2033) | ~_GEN_1051
         & (dis_ld_val_1
              ? ~_GEN_930 & ldq_0_bits_executed
              : ~_GEN_855 & ldq_0_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_0_bits_succeeded <=
      _GEN_2325 & _GEN_2277 & _GEN_2229
      & (_GEN_2061
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h0
                ? _ldq_bits_succeeded_T
                : ~_GEN_1051
                  & (dis_ld_val_1
                       ? ~_GEN_930 & ldq_0_bits_succeeded
                       : ~_GEN_855 & ldq_0_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_0_bits_order_fail <=
      _GEN_2325 & _GEN_2277 & _GEN_2229
      & (_GEN_327
           ? _GEN_1123
           : _GEN_332
               ? _GEN_1387 | _GEN_1123
               : _GEN_333 & searcher_is_older & _GEN_1388 | _GEN_1123);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_0_bits_observed <=
      _GEN_327 | ~_GEN_1051
      & (dis_ld_val_1
           ? ~_GEN_930 & ldq_0_bits_observed
           : ~_GEN_855 & ldq_0_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_0_bits_forward_std_val <=
      _GEN_2325 & _GEN_2277 & _GEN_2229
      & (~_GEN_787 & _GEN_2060 | ~_GEN_1051
         & (dis_ld_val_1
              ? ~_GEN_930 & ldq_0_bits_forward_std_val
              : ~_GEN_855 & ldq_0_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2061) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_0_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_1_valid <=
      ~_GEN_2424 & _GEN_2326 & _GEN_2278
      & (_GEN_2205 ? ~_GEN_2133 & _GEN_1054 : ~_GEN_2206 & _GEN_1054);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1053) begin	// lsu.scala:304:5, :305:44
      ldq_1_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_1_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_1_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_1_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_1_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_1_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_1_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_1_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_1_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_978) begin	// lsu.scala:304:5, :306:44
      ldq_1_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_1_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_1_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_1_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_1_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_1_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_1_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_856) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_1_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_1_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_1_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_1_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_1_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_1_valid)	// lsu.scala:210:16
      ldq_1_bits_uop_br_mask <=
        ldq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1053)	// lsu.scala:304:5, :305:44
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_978)	// lsu.scala:304:5, :306:44
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_856)	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1245) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_1_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_1_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_1_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_1_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_1_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_1_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_1_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_1_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_1_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_1_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_1_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1053)	// lsu.scala:304:5, :305:44
      ldq_1_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_978)	// lsu.scala:304:5, :306:44
      ldq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_856)	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1100)	// lsu.scala:210:16, :304:5, :306:44
      ldq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_1_bits_uop_ppred_busy <= ~_GEN_1100 & ldq_1_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_1_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h1
      | (_GEN_1053
           ? io_core_dis_uops_2_bits_exception
           : _GEN_978
               ? io_core_dis_uops_1_bits_exception
               : _GEN_856 ? io_core_dis_uops_0_bits_exception : ldq_1_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_1_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2326 & _GEN_2278
      & (_GEN_2205 ? ~_GEN_2133 & _GEN_1246 : ~_GEN_2206 & _GEN_1246);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_1_bits_executed <=
      ~_GEN_2424 & _GEN_2326 & _GEN_2278 & _GEN_2230
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_762))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1389 & _GEN_2034 : ~(_GEN_757 & _GEN_1389) & _GEN_2034)
            : _GEN_2034) | ~_GEN_1053
         & (dis_ld_val_1
              ? ~_GEN_932 & ldq_1_bits_executed
              : ~_GEN_856 & ldq_1_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_1_bits_succeeded <=
      _GEN_2326 & _GEN_2278 & _GEN_2230
      & (_GEN_2063
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1
                ? _ldq_bits_succeeded_T
                : ~_GEN_1053
                  & (dis_ld_val_1
                       ? ~_GEN_932 & ldq_1_bits_succeeded
                       : ~_GEN_856 & ldq_1_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_1_bits_order_fail <=
      _GEN_2326 & _GEN_2278 & _GEN_2230
      & (_GEN_338
           ? _GEN_1124
           : _GEN_342
               ? _GEN_1412 | _GEN_1124
               : _GEN_343 & searcher_is_older_1 & _GEN_1413 | _GEN_1124);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_1_bits_observed <=
      _GEN_338 | ~_GEN_1053
      & (dis_ld_val_1
           ? ~_GEN_932 & ldq_1_bits_observed
           : ~_GEN_856 & ldq_1_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_1_bits_forward_std_val <=
      _GEN_2326 & _GEN_2278 & _GEN_2230
      & (~_GEN_787 & _GEN_2062 | ~_GEN_1053
         & (dis_ld_val_1
              ? ~_GEN_932 & ldq_1_bits_forward_std_val
              : ~_GEN_856 & ldq_1_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2063) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_1_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_2_valid <=
      ~_GEN_2424 & _GEN_2327 & _GEN_2279
      & (_GEN_2205 ? ~_GEN_2134 & _GEN_1056 : ~_GEN_2207 & _GEN_1056);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1055) begin	// lsu.scala:304:5, :305:44
      ldq_2_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_2_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_2_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_2_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_2_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_2_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_2_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_2_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_2_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_979) begin	// lsu.scala:304:5, :306:44
      ldq_2_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_2_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_2_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_2_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_2_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_2_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_2_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_857) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_2_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_2_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_2_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_2_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_2_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_2_valid)	// lsu.scala:210:16
      ldq_2_bits_uop_br_mask <=
        ldq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1055)	// lsu.scala:304:5, :305:44
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_979)	// lsu.scala:304:5, :306:44
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_857)	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1247) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_2_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_2_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_2_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_2_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_2_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_2_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_2_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_2_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_2_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_2_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_2_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1055)	// lsu.scala:304:5, :305:44
      ldq_2_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_979)	// lsu.scala:304:5, :306:44
      ldq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_857)	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1101)	// lsu.scala:210:16, :304:5, :306:44
      ldq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_2_bits_uop_ppred_busy <= ~_GEN_1101 & ldq_2_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_2_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h2
      | (_GEN_1055
           ? io_core_dis_uops_2_bits_exception
           : _GEN_979
               ? io_core_dis_uops_1_bits_exception
               : _GEN_857 ? io_core_dis_uops_0_bits_exception : ldq_2_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_2_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2327 & _GEN_2279
      & (_GEN_2205 ? ~_GEN_2134 & _GEN_1248 : ~_GEN_2207 & _GEN_1248);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_2_bits_executed <=
      ~_GEN_2424 & _GEN_2327 & _GEN_2279 & _GEN_2231
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_763))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1390 & _GEN_2035 : ~(_GEN_757 & _GEN_1390) & _GEN_2035)
            : _GEN_2035) | ~_GEN_1055
         & (dis_ld_val_1
              ? ~_GEN_934 & ldq_2_bits_executed
              : ~_GEN_857 & ldq_2_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_2_bits_succeeded <=
      _GEN_2327 & _GEN_2279 & _GEN_2231
      & (_GEN_2065
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h2
                ? _ldq_bits_succeeded_T
                : ~_GEN_1055
                  & (dis_ld_val_1
                       ? ~_GEN_934 & ldq_2_bits_succeeded
                       : ~_GEN_857 & ldq_2_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_2_bits_order_fail <=
      _GEN_2327 & _GEN_2279 & _GEN_2231
      & (_GEN_349
           ? _GEN_1125
           : _GEN_353
               ? _GEN_1414 | _GEN_1125
               : _GEN_354 & searcher_is_older_2 & _GEN_1415 | _GEN_1125);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_2_bits_observed <=
      _GEN_349 | ~_GEN_1055
      & (dis_ld_val_1
           ? ~_GEN_934 & ldq_2_bits_observed
           : ~_GEN_857 & ldq_2_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_2_bits_forward_std_val <=
      _GEN_2327 & _GEN_2279 & _GEN_2231
      & (~_GEN_787 & _GEN_2064 | ~_GEN_1055
         & (dis_ld_val_1
              ? ~_GEN_934 & ldq_2_bits_forward_std_val
              : ~_GEN_857 & ldq_2_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2065) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_2_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_3_valid <=
      ~_GEN_2424 & _GEN_2328 & _GEN_2280
      & (_GEN_2205 ? ~_GEN_2135 & _GEN_1058 : ~_GEN_2208 & _GEN_1058);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1057) begin	// lsu.scala:304:5, :305:44
      ldq_3_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_3_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_3_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_3_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_3_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_3_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_3_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_3_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_3_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_980) begin	// lsu.scala:304:5, :306:44
      ldq_3_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_3_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_3_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_3_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_3_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_3_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_3_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_858) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_3_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_3_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_3_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_3_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_3_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_3_valid)	// lsu.scala:210:16
      ldq_3_bits_uop_br_mask <=
        ldq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1057)	// lsu.scala:304:5, :305:44
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_980)	// lsu.scala:304:5, :306:44
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_858)	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1249) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_3_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_3_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_3_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_3_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_3_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_3_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_3_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_3_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_3_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_3_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_3_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1057)	// lsu.scala:304:5, :305:44
      ldq_3_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_980)	// lsu.scala:304:5, :306:44
      ldq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_858)	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1102)	// lsu.scala:210:16, :304:5, :306:44
      ldq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_3_bits_uop_ppred_busy <= ~_GEN_1102 & ldq_3_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_3_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h3
      | (_GEN_1057
           ? io_core_dis_uops_2_bits_exception
           : _GEN_980
               ? io_core_dis_uops_1_bits_exception
               : _GEN_858 ? io_core_dis_uops_0_bits_exception : ldq_3_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_3_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2328 & _GEN_2280
      & (_GEN_2205 ? ~_GEN_2135 & _GEN_1250 : ~_GEN_2208 & _GEN_1250);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_3_bits_executed <=
      ~_GEN_2424 & _GEN_2328 & _GEN_2280 & _GEN_2232
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_764))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1391 & _GEN_2036 : ~(_GEN_757 & _GEN_1391) & _GEN_2036)
            : _GEN_2036) | ~_GEN_1057
         & (dis_ld_val_1
              ? ~_GEN_936 & ldq_3_bits_executed
              : ~_GEN_858 & ldq_3_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_3_bits_succeeded <=
      _GEN_2328 & _GEN_2280 & _GEN_2232
      & (_GEN_2067
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h3
                ? _ldq_bits_succeeded_T
                : ~_GEN_1057
                  & (dis_ld_val_1
                       ? ~_GEN_936 & ldq_3_bits_succeeded
                       : ~_GEN_858 & ldq_3_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_3_bits_order_fail <=
      _GEN_2328 & _GEN_2280 & _GEN_2232
      & (_GEN_360
           ? _GEN_1126
           : _GEN_364
               ? _GEN_1416 | _GEN_1126
               : _GEN_365 & searcher_is_older_3 & _GEN_1417 | _GEN_1126);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_3_bits_observed <=
      _GEN_360 | ~_GEN_1057
      & (dis_ld_val_1
           ? ~_GEN_936 & ldq_3_bits_observed
           : ~_GEN_858 & ldq_3_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_3_bits_forward_std_val <=
      _GEN_2328 & _GEN_2280 & _GEN_2232
      & (~_GEN_787 & _GEN_2066 | ~_GEN_1057
         & (dis_ld_val_1
              ? ~_GEN_936 & ldq_3_bits_forward_std_val
              : ~_GEN_858 & ldq_3_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2067) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_3_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_4_valid <=
      ~_GEN_2424 & _GEN_2329 & _GEN_2281
      & (_GEN_2205 ? ~_GEN_2136 & _GEN_1060 : ~_GEN_2209 & _GEN_1060);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1059) begin	// lsu.scala:304:5, :305:44
      ldq_4_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_4_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_4_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_4_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_4_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_4_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_4_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_4_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_4_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_981) begin	// lsu.scala:304:5, :306:44
      ldq_4_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_4_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_4_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_4_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_4_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_4_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_4_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_859) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_4_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_4_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_4_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_4_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_4_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_4_valid)	// lsu.scala:210:16
      ldq_4_bits_uop_br_mask <=
        ldq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1059)	// lsu.scala:304:5, :305:44
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_981)	// lsu.scala:304:5, :306:44
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_859)	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1251) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_4_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_4_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_4_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_4_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_4_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_4_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_4_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_4_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_4_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_4_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_4_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1059)	// lsu.scala:304:5, :305:44
      ldq_4_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_981)	// lsu.scala:304:5, :306:44
      ldq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_859)	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1103)	// lsu.scala:210:16, :304:5, :306:44
      ldq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_4_bits_uop_ppred_busy <= ~_GEN_1103 & ldq_4_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_4_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h4
      | (_GEN_1059
           ? io_core_dis_uops_2_bits_exception
           : _GEN_981
               ? io_core_dis_uops_1_bits_exception
               : _GEN_859 ? io_core_dis_uops_0_bits_exception : ldq_4_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_4_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2329 & _GEN_2281
      & (_GEN_2205 ? ~_GEN_2136 & _GEN_1252 : ~_GEN_2209 & _GEN_1252);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_4_bits_executed <=
      ~_GEN_2424 & _GEN_2329 & _GEN_2281 & _GEN_2233
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_765))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1392 & _GEN_2037 : ~(_GEN_757 & _GEN_1392) & _GEN_2037)
            : _GEN_2037) | ~_GEN_1059
         & (dis_ld_val_1
              ? ~_GEN_938 & ldq_4_bits_executed
              : ~_GEN_859 & ldq_4_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_4_bits_succeeded <=
      _GEN_2329 & _GEN_2281 & _GEN_2233
      & (_GEN_2069
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h4
                ? _ldq_bits_succeeded_T
                : ~_GEN_1059
                  & (dis_ld_val_1
                       ? ~_GEN_938 & ldq_4_bits_succeeded
                       : ~_GEN_859 & ldq_4_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_4_bits_order_fail <=
      _GEN_2329 & _GEN_2281 & _GEN_2233
      & (_GEN_371
           ? _GEN_1127
           : _GEN_375
               ? _GEN_1418 | _GEN_1127
               : _GEN_376 & searcher_is_older_4 & _GEN_1419 | _GEN_1127);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_4_bits_observed <=
      _GEN_371 | ~_GEN_1059
      & (dis_ld_val_1
           ? ~_GEN_938 & ldq_4_bits_observed
           : ~_GEN_859 & ldq_4_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_4_bits_forward_std_val <=
      _GEN_2329 & _GEN_2281 & _GEN_2233
      & (~_GEN_787 & _GEN_2068 | ~_GEN_1059
         & (dis_ld_val_1
              ? ~_GEN_938 & ldq_4_bits_forward_std_val
              : ~_GEN_859 & ldq_4_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2069) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_4_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_5_valid <=
      ~_GEN_2424 & _GEN_2330 & _GEN_2282
      & (_GEN_2205 ? ~_GEN_2137 & _GEN_1062 : ~_GEN_2210 & _GEN_1062);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1061) begin	// lsu.scala:304:5, :305:44
      ldq_5_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_5_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_5_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_5_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_5_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_5_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_5_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_5_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_5_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_982) begin	// lsu.scala:304:5, :306:44
      ldq_5_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_5_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_5_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_5_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_5_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_5_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_5_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_860) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_5_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_5_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_5_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_5_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_5_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_5_valid)	// lsu.scala:210:16
      ldq_5_bits_uop_br_mask <=
        ldq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1061)	// lsu.scala:304:5, :305:44
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_982)	// lsu.scala:304:5, :306:44
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_860)	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1253) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_5_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_5_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_5_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_5_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_5_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_5_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_5_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_5_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_5_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_5_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_5_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1061)	// lsu.scala:304:5, :305:44
      ldq_5_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_982)	// lsu.scala:304:5, :306:44
      ldq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_860)	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1104)	// lsu.scala:210:16, :304:5, :306:44
      ldq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_5_bits_uop_ppred_busy <= ~_GEN_1104 & ldq_5_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_5_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h5
      | (_GEN_1061
           ? io_core_dis_uops_2_bits_exception
           : _GEN_982
               ? io_core_dis_uops_1_bits_exception
               : _GEN_860 ? io_core_dis_uops_0_bits_exception : ldq_5_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_5_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2330 & _GEN_2282
      & (_GEN_2205 ? ~_GEN_2137 & _GEN_1254 : ~_GEN_2210 & _GEN_1254);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_5_bits_executed <=
      ~_GEN_2424 & _GEN_2330 & _GEN_2282 & _GEN_2234
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_766))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1393 & _GEN_2038 : ~(_GEN_757 & _GEN_1393) & _GEN_2038)
            : _GEN_2038) | ~_GEN_1061
         & (dis_ld_val_1
              ? ~_GEN_940 & ldq_5_bits_executed
              : ~_GEN_860 & ldq_5_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_5_bits_succeeded <=
      _GEN_2330 & _GEN_2282 & _GEN_2234
      & (_GEN_2071
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h5
                ? _ldq_bits_succeeded_T
                : ~_GEN_1061
                  & (dis_ld_val_1
                       ? ~_GEN_940 & ldq_5_bits_succeeded
                       : ~_GEN_860 & ldq_5_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_5_bits_order_fail <=
      _GEN_2330 & _GEN_2282 & _GEN_2234
      & (_GEN_382
           ? _GEN_1128
           : _GEN_386
               ? _GEN_1420 | _GEN_1128
               : _GEN_387 & searcher_is_older_5 & _GEN_1421 | _GEN_1128);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_5_bits_observed <=
      _GEN_382 | ~_GEN_1061
      & (dis_ld_val_1
           ? ~_GEN_940 & ldq_5_bits_observed
           : ~_GEN_860 & ldq_5_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_5_bits_forward_std_val <=
      _GEN_2330 & _GEN_2282 & _GEN_2234
      & (~_GEN_787 & _GEN_2070 | ~_GEN_1061
         & (dis_ld_val_1
              ? ~_GEN_940 & ldq_5_bits_forward_std_val
              : ~_GEN_860 & ldq_5_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2071) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_5_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_6_valid <=
      ~_GEN_2424 & _GEN_2331 & _GEN_2283
      & (_GEN_2205 ? ~_GEN_2138 & _GEN_1064 : ~_GEN_2211 & _GEN_1064);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1063) begin	// lsu.scala:304:5, :305:44
      ldq_6_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_6_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_6_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_6_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_6_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_6_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_6_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_6_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_6_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_983) begin	// lsu.scala:304:5, :306:44
      ldq_6_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_6_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_6_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_6_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_6_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_6_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_6_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_861) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_6_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_6_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_6_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_6_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_6_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_6_valid)	// lsu.scala:210:16
      ldq_6_bits_uop_br_mask <=
        ldq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1063)	// lsu.scala:304:5, :305:44
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_983)	// lsu.scala:304:5, :306:44
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_861)	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1255) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_6_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_6_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_6_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_6_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_6_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_6_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_6_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_6_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_6_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_6_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_6_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1063)	// lsu.scala:304:5, :305:44
      ldq_6_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_983)	// lsu.scala:304:5, :306:44
      ldq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_861)	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1105)	// lsu.scala:210:16, :304:5, :306:44
      ldq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_6_bits_uop_ppred_busy <= ~_GEN_1105 & ldq_6_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_6_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h6
      | (_GEN_1063
           ? io_core_dis_uops_2_bits_exception
           : _GEN_983
               ? io_core_dis_uops_1_bits_exception
               : _GEN_861 ? io_core_dis_uops_0_bits_exception : ldq_6_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_6_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2331 & _GEN_2283
      & (_GEN_2205 ? ~_GEN_2138 & _GEN_1256 : ~_GEN_2211 & _GEN_1256);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_6_bits_executed <=
      ~_GEN_2424 & _GEN_2331 & _GEN_2283 & _GEN_2235
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_767))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1394 & _GEN_2039 : ~(_GEN_757 & _GEN_1394) & _GEN_2039)
            : _GEN_2039) | ~_GEN_1063
         & (dis_ld_val_1
              ? ~_GEN_942 & ldq_6_bits_executed
              : ~_GEN_861 & ldq_6_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_6_bits_succeeded <=
      _GEN_2331 & _GEN_2283 & _GEN_2235
      & (_GEN_2073
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h6
                ? _ldq_bits_succeeded_T
                : ~_GEN_1063
                  & (dis_ld_val_1
                       ? ~_GEN_942 & ldq_6_bits_succeeded
                       : ~_GEN_861 & ldq_6_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_6_bits_order_fail <=
      _GEN_2331 & _GEN_2283 & _GEN_2235
      & (_GEN_393
           ? _GEN_1129
           : _GEN_397
               ? _GEN_1422 | _GEN_1129
               : _GEN_398 & searcher_is_older_6 & _GEN_1423 | _GEN_1129);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_6_bits_observed <=
      _GEN_393 | ~_GEN_1063
      & (dis_ld_val_1
           ? ~_GEN_942 & ldq_6_bits_observed
           : ~_GEN_861 & ldq_6_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_6_bits_forward_std_val <=
      _GEN_2331 & _GEN_2283 & _GEN_2235
      & (~_GEN_787 & _GEN_2072 | ~_GEN_1063
         & (dis_ld_val_1
              ? ~_GEN_942 & ldq_6_bits_forward_std_val
              : ~_GEN_861 & ldq_6_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2073) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_6_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_7_valid <=
      ~_GEN_2424 & _GEN_2332 & _GEN_2284
      & (_GEN_2205 ? ~_GEN_2139 & _GEN_1066 : ~_GEN_2212 & _GEN_1066);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1065) begin	// lsu.scala:304:5, :305:44
      ldq_7_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_7_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_7_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_7_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_7_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_7_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_7_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_7_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_7_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_984) begin	// lsu.scala:304:5, :306:44
      ldq_7_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_7_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_7_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_7_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_7_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_7_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_7_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_862) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_7_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_7_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_7_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_7_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_7_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_7_valid)	// lsu.scala:210:16
      ldq_7_bits_uop_br_mask <=
        ldq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1065)	// lsu.scala:304:5, :305:44
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_984)	// lsu.scala:304:5, :306:44
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_862)	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1257) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_7_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_7_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_7_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_7_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_7_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_7_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_7_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_7_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_7_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_7_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_7_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1065)	// lsu.scala:304:5, :305:44
      ldq_7_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_984)	// lsu.scala:304:5, :306:44
      ldq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_862)	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1106)	// lsu.scala:210:16, :304:5, :306:44
      ldq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_7_bits_uop_ppred_busy <= ~_GEN_1106 & ldq_7_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_7_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h7
      | (_GEN_1065
           ? io_core_dis_uops_2_bits_exception
           : _GEN_984
               ? io_core_dis_uops_1_bits_exception
               : _GEN_862 ? io_core_dis_uops_0_bits_exception : ldq_7_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_7_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2332 & _GEN_2284
      & (_GEN_2205 ? ~_GEN_2139 & _GEN_1258 : ~_GEN_2212 & _GEN_1258);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_7_bits_executed <=
      ~_GEN_2424 & _GEN_2332 & _GEN_2284 & _GEN_2236
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_768))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1395 & _GEN_2040 : ~(_GEN_757 & _GEN_1395) & _GEN_2040)
            : _GEN_2040) | ~_GEN_1065
         & (dis_ld_val_1
              ? ~_GEN_944 & ldq_7_bits_executed
              : ~_GEN_862 & ldq_7_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_7_bits_succeeded <=
      _GEN_2332 & _GEN_2284 & _GEN_2236
      & (_GEN_2075
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h7
                ? _ldq_bits_succeeded_T
                : ~_GEN_1065
                  & (dis_ld_val_1
                       ? ~_GEN_944 & ldq_7_bits_succeeded
                       : ~_GEN_862 & ldq_7_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_7_bits_order_fail <=
      _GEN_2332 & _GEN_2284 & _GEN_2236
      & (_GEN_404
           ? _GEN_1130
           : _GEN_408
               ? _GEN_1424 | _GEN_1130
               : _GEN_409 & searcher_is_older_7 & _GEN_1425 | _GEN_1130);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_7_bits_observed <=
      _GEN_404 | ~_GEN_1065
      & (dis_ld_val_1
           ? ~_GEN_944 & ldq_7_bits_observed
           : ~_GEN_862 & ldq_7_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_7_bits_forward_std_val <=
      _GEN_2332 & _GEN_2284 & _GEN_2236
      & (~_GEN_787 & _GEN_2074 | ~_GEN_1065
         & (dis_ld_val_1
              ? ~_GEN_944 & ldq_7_bits_forward_std_val
              : ~_GEN_862 & ldq_7_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2075) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_7_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_8_valid <=
      ~_GEN_2424 & _GEN_2333 & _GEN_2285
      & (_GEN_2205 ? ~_GEN_2140 & _GEN_1068 : ~_GEN_2213 & _GEN_1068);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1067) begin	// lsu.scala:304:5, :305:44
      ldq_8_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_8_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_8_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_8_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_8_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_8_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_8_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_8_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_8_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_985) begin	// lsu.scala:304:5, :306:44
      ldq_8_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_8_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_8_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_8_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_8_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_8_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_8_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_863) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_8_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_8_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_8_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_8_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_8_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_8_valid)	// lsu.scala:210:16
      ldq_8_bits_uop_br_mask <=
        ldq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1067)	// lsu.scala:304:5, :305:44
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_985)	// lsu.scala:304:5, :306:44
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_863)	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1259) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_8_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_8_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_8_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_8_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_8_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_8_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_8_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_8_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_8_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_8_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_8_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1067)	// lsu.scala:304:5, :305:44
      ldq_8_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_985)	// lsu.scala:304:5, :306:44
      ldq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_863)	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1107)	// lsu.scala:210:16, :304:5, :306:44
      ldq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_8_bits_uop_ppred_busy <= ~_GEN_1107 & ldq_8_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_8_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h8
      | (_GEN_1067
           ? io_core_dis_uops_2_bits_exception
           : _GEN_985
               ? io_core_dis_uops_1_bits_exception
               : _GEN_863 ? io_core_dis_uops_0_bits_exception : ldq_8_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_8_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2333 & _GEN_2285
      & (_GEN_2205 ? ~_GEN_2140 & _GEN_1260 : ~_GEN_2213 & _GEN_1260);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_8_bits_executed <=
      ~_GEN_2424 & _GEN_2333 & _GEN_2285 & _GEN_2237
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_769))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1396 & _GEN_2041 : ~(_GEN_757 & _GEN_1396) & _GEN_2041)
            : _GEN_2041) | ~_GEN_1067
         & (dis_ld_val_1
              ? ~_GEN_946 & ldq_8_bits_executed
              : ~_GEN_863 & ldq_8_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_8_bits_succeeded <=
      _GEN_2333 & _GEN_2285 & _GEN_2237
      & (_GEN_2077
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h8
                ? _ldq_bits_succeeded_T
                : ~_GEN_1067
                  & (dis_ld_val_1
                       ? ~_GEN_946 & ldq_8_bits_succeeded
                       : ~_GEN_863 & ldq_8_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_8_bits_order_fail <=
      _GEN_2333 & _GEN_2285 & _GEN_2237
      & (_GEN_415
           ? _GEN_1131
           : _GEN_419
               ? _GEN_1426 | _GEN_1131
               : _GEN_420 & searcher_is_older_8 & _GEN_1427 | _GEN_1131);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_8_bits_observed <=
      _GEN_415 | ~_GEN_1067
      & (dis_ld_val_1
           ? ~_GEN_946 & ldq_8_bits_observed
           : ~_GEN_863 & ldq_8_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_8_bits_forward_std_val <=
      _GEN_2333 & _GEN_2285 & _GEN_2237
      & (~_GEN_787 & _GEN_2076 | ~_GEN_1067
         & (dis_ld_val_1
              ? ~_GEN_946 & ldq_8_bits_forward_std_val
              : ~_GEN_863 & ldq_8_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2077) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_8_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_9_valid <=
      ~_GEN_2424 & _GEN_2334 & _GEN_2286
      & (_GEN_2205 ? ~_GEN_2141 & _GEN_1070 : ~_GEN_2214 & _GEN_1070);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1069) begin	// lsu.scala:304:5, :305:44
      ldq_9_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_9_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_9_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_9_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_9_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_9_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_9_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_9_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_9_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_986) begin	// lsu.scala:304:5, :306:44
      ldq_9_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_9_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_9_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_9_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_9_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_9_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_9_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_864) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_9_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_9_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_9_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_9_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_9_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_9_valid)	// lsu.scala:210:16
      ldq_9_bits_uop_br_mask <=
        ldq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1069)	// lsu.scala:304:5, :305:44
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_986)	// lsu.scala:304:5, :306:44
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_864)	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1261) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_9_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_9_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_9_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_9_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_9_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_9_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_9_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_9_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_9_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_9_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_9_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1069)	// lsu.scala:304:5, :305:44
      ldq_9_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_986)	// lsu.scala:304:5, :306:44
      ldq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_864)	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1108)	// lsu.scala:210:16, :304:5, :306:44
      ldq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_9_bits_uop_ppred_busy <= ~_GEN_1108 & ldq_9_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_9_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h9
      | (_GEN_1069
           ? io_core_dis_uops_2_bits_exception
           : _GEN_986
               ? io_core_dis_uops_1_bits_exception
               : _GEN_864 ? io_core_dis_uops_0_bits_exception : ldq_9_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_9_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2334 & _GEN_2286
      & (_GEN_2205 ? ~_GEN_2141 & _GEN_1262 : ~_GEN_2214 & _GEN_1262);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_9_bits_executed <=
      ~_GEN_2424 & _GEN_2334 & _GEN_2286 & _GEN_2238
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_770))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1397 & _GEN_2042 : ~(_GEN_757 & _GEN_1397) & _GEN_2042)
            : _GEN_2042) | ~_GEN_1069
         & (dis_ld_val_1
              ? ~_GEN_948 & ldq_9_bits_executed
              : ~_GEN_864 & ldq_9_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_9_bits_succeeded <=
      _GEN_2334 & _GEN_2286 & _GEN_2238
      & (_GEN_2079
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h9
                ? _ldq_bits_succeeded_T
                : ~_GEN_1069
                  & (dis_ld_val_1
                       ? ~_GEN_948 & ldq_9_bits_succeeded
                       : ~_GEN_864 & ldq_9_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_9_bits_order_fail <=
      _GEN_2334 & _GEN_2286 & _GEN_2238
      & (_GEN_426
           ? _GEN_1132
           : _GEN_430
               ? _GEN_1428 | _GEN_1132
               : _GEN_431 & searcher_is_older_9 & _GEN_1429 | _GEN_1132);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_9_bits_observed <=
      _GEN_426 | ~_GEN_1069
      & (dis_ld_val_1
           ? ~_GEN_948 & ldq_9_bits_observed
           : ~_GEN_864 & ldq_9_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_9_bits_forward_std_val <=
      _GEN_2334 & _GEN_2286 & _GEN_2238
      & (~_GEN_787 & _GEN_2078 | ~_GEN_1069
         & (dis_ld_val_1
              ? ~_GEN_948 & ldq_9_bits_forward_std_val
              : ~_GEN_864 & ldq_9_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2079) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_9_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_10_valid <=
      ~_GEN_2424 & _GEN_2335 & _GEN_2287
      & (_GEN_2205 ? ~_GEN_2142 & _GEN_1072 : ~_GEN_2215 & _GEN_1072);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1071) begin	// lsu.scala:304:5, :305:44
      ldq_10_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_10_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_10_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_10_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_10_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_10_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_10_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_10_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_10_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_987) begin	// lsu.scala:304:5, :306:44
      ldq_10_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_10_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_10_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_10_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_10_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_10_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_10_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_865) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_10_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_10_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_10_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_10_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_10_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_10_valid)	// lsu.scala:210:16
      ldq_10_bits_uop_br_mask <=
        ldq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1071)	// lsu.scala:304:5, :305:44
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_987)	// lsu.scala:304:5, :306:44
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_865)	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1263) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_10_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_10_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_10_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_10_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_10_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_10_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_10_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_10_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_10_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_10_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_10_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1071)	// lsu.scala:304:5, :305:44
      ldq_10_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_987)	// lsu.scala:304:5, :306:44
      ldq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_865)	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1109)	// lsu.scala:210:16, :304:5, :306:44
      ldq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_10_bits_uop_ppred_busy <= ~_GEN_1109 & ldq_10_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_10_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hA
      | (_GEN_1071
           ? io_core_dis_uops_2_bits_exception
           : _GEN_987
               ? io_core_dis_uops_1_bits_exception
               : _GEN_865
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_10_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_10_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2335 & _GEN_2287
      & (_GEN_2205 ? ~_GEN_2142 & _GEN_1264 : ~_GEN_2215 & _GEN_1264);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_10_bits_executed <=
      ~_GEN_2424 & _GEN_2335 & _GEN_2287 & _GEN_2239
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_771))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1398 & _GEN_2043 : ~(_GEN_757 & _GEN_1398) & _GEN_2043)
            : _GEN_2043) | ~_GEN_1071
         & (dis_ld_val_1
              ? ~_GEN_950 & ldq_10_bits_executed
              : ~_GEN_865 & ldq_10_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_10_bits_succeeded <=
      _GEN_2335 & _GEN_2287 & _GEN_2239
      & (_GEN_2081
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'hA
                ? _ldq_bits_succeeded_T
                : ~_GEN_1071
                  & (dis_ld_val_1
                       ? ~_GEN_950 & ldq_10_bits_succeeded
                       : ~_GEN_865 & ldq_10_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_10_bits_order_fail <=
      _GEN_2335 & _GEN_2287 & _GEN_2239
      & (_GEN_437
           ? _GEN_1133
           : _GEN_441
               ? _GEN_1430 | _GEN_1133
               : _GEN_442 & searcher_is_older_10 & _GEN_1431 | _GEN_1133);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_10_bits_observed <=
      _GEN_437 | ~_GEN_1071
      & (dis_ld_val_1
           ? ~_GEN_950 & ldq_10_bits_observed
           : ~_GEN_865 & ldq_10_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_10_bits_forward_std_val <=
      _GEN_2335 & _GEN_2287 & _GEN_2239
      & (~_GEN_787 & _GEN_2080 | ~_GEN_1071
         & (dis_ld_val_1
              ? ~_GEN_950 & ldq_10_bits_forward_std_val
              : ~_GEN_865 & ldq_10_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2081) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_10_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_11_valid <=
      ~_GEN_2424 & _GEN_2336 & _GEN_2288
      & (_GEN_2205 ? ~_GEN_2143 & _GEN_1074 : ~_GEN_2216 & _GEN_1074);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1073) begin	// lsu.scala:304:5, :305:44
      ldq_11_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_11_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_11_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_11_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_11_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_11_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_11_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_11_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_11_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_988) begin	// lsu.scala:304:5, :306:44
      ldq_11_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_11_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_11_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_11_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_11_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_11_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_11_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_866) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_11_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_11_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_11_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_11_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_11_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_11_valid)	// lsu.scala:210:16
      ldq_11_bits_uop_br_mask <=
        ldq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1073)	// lsu.scala:304:5, :305:44
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_988)	// lsu.scala:304:5, :306:44
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_866)	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1265) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_11_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_11_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_11_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_11_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_11_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_11_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_11_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_11_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_11_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_11_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_11_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1073)	// lsu.scala:304:5, :305:44
      ldq_11_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_988)	// lsu.scala:304:5, :306:44
      ldq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_866)	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1110)	// lsu.scala:210:16, :304:5, :306:44
      ldq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_11_bits_uop_ppred_busy <= ~_GEN_1110 & ldq_11_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_11_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hB
      | (_GEN_1073
           ? io_core_dis_uops_2_bits_exception
           : _GEN_988
               ? io_core_dis_uops_1_bits_exception
               : _GEN_866
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_11_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_11_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2336 & _GEN_2288
      & (_GEN_2205 ? ~_GEN_2143 & _GEN_1266 : ~_GEN_2216 & _GEN_1266);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_11_bits_executed <=
      ~_GEN_2424 & _GEN_2336 & _GEN_2288 & _GEN_2240
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_772))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1399 & _GEN_2044 : ~(_GEN_757 & _GEN_1399) & _GEN_2044)
            : _GEN_2044) | ~_GEN_1073
         & (dis_ld_val_1
              ? ~_GEN_952 & ldq_11_bits_executed
              : ~_GEN_866 & ldq_11_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_11_bits_succeeded <=
      _GEN_2336 & _GEN_2288 & _GEN_2240
      & (_GEN_2083
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'hB
                ? _ldq_bits_succeeded_T
                : ~_GEN_1073
                  & (dis_ld_val_1
                       ? ~_GEN_952 & ldq_11_bits_succeeded
                       : ~_GEN_866 & ldq_11_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_11_bits_order_fail <=
      _GEN_2336 & _GEN_2288 & _GEN_2240
      & (_GEN_448
           ? _GEN_1134
           : _GEN_452
               ? _GEN_1432 | _GEN_1134
               : _GEN_453 & searcher_is_older_11 & _GEN_1433 | _GEN_1134);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_11_bits_observed <=
      _GEN_448 | ~_GEN_1073
      & (dis_ld_val_1
           ? ~_GEN_952 & ldq_11_bits_observed
           : ~_GEN_866 & ldq_11_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_11_bits_forward_std_val <=
      _GEN_2336 & _GEN_2288 & _GEN_2240
      & (~_GEN_787 & _GEN_2082 | ~_GEN_1073
         & (dis_ld_val_1
              ? ~_GEN_952 & ldq_11_bits_forward_std_val
              : ~_GEN_866 & ldq_11_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2083) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_11_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_12_valid <=
      ~_GEN_2424 & _GEN_2337 & _GEN_2289
      & (_GEN_2205 ? ~_GEN_2144 & _GEN_1076 : ~_GEN_2217 & _GEN_1076);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1075) begin	// lsu.scala:304:5, :305:44
      ldq_12_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_12_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_12_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_12_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_12_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_12_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_12_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_12_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_12_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_989) begin	// lsu.scala:304:5, :306:44
      ldq_12_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_12_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_12_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_12_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_12_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_12_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_12_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_867) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_12_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_12_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_12_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_12_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_12_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_12_valid)	// lsu.scala:210:16
      ldq_12_bits_uop_br_mask <=
        ldq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1075)	// lsu.scala:304:5, :305:44
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_989)	// lsu.scala:304:5, :306:44
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_867)	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1267) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_12_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_12_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_12_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_12_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_12_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_12_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_12_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_12_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_12_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_12_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_12_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1075)	// lsu.scala:304:5, :305:44
      ldq_12_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_989)	// lsu.scala:304:5, :306:44
      ldq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_867)	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1111)	// lsu.scala:210:16, :304:5, :306:44
      ldq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_12_bits_uop_ppred_busy <= ~_GEN_1111 & ldq_12_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_12_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hC
      | (_GEN_1075
           ? io_core_dis_uops_2_bits_exception
           : _GEN_989
               ? io_core_dis_uops_1_bits_exception
               : _GEN_867
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_12_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_12_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2337 & _GEN_2289
      & (_GEN_2205 ? ~_GEN_2144 & _GEN_1268 : ~_GEN_2217 & _GEN_1268);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_12_bits_executed <=
      ~_GEN_2424 & _GEN_2337 & _GEN_2289 & _GEN_2241
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_773))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1400 & _GEN_2045 : ~(_GEN_757 & _GEN_1400) & _GEN_2045)
            : _GEN_2045) | ~_GEN_1075
         & (dis_ld_val_1
              ? ~_GEN_954 & ldq_12_bits_executed
              : ~_GEN_867 & ldq_12_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_12_bits_succeeded <=
      _GEN_2337 & _GEN_2289 & _GEN_2241
      & (_GEN_2085
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'hC
                ? _ldq_bits_succeeded_T
                : ~_GEN_1075
                  & (dis_ld_val_1
                       ? ~_GEN_954 & ldq_12_bits_succeeded
                       : ~_GEN_867 & ldq_12_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_12_bits_order_fail <=
      _GEN_2337 & _GEN_2289 & _GEN_2241
      & (_GEN_459
           ? _GEN_1135
           : _GEN_463
               ? _GEN_1434 | _GEN_1135
               : _GEN_464 & searcher_is_older_12 & _GEN_1435 | _GEN_1135);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_12_bits_observed <=
      _GEN_459 | ~_GEN_1075
      & (dis_ld_val_1
           ? ~_GEN_954 & ldq_12_bits_observed
           : ~_GEN_867 & ldq_12_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_12_bits_forward_std_val <=
      _GEN_2337 & _GEN_2289 & _GEN_2241
      & (~_GEN_787 & _GEN_2084 | ~_GEN_1075
         & (dis_ld_val_1
              ? ~_GEN_954 & ldq_12_bits_forward_std_val
              : ~_GEN_867 & ldq_12_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2085) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_12_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_13_valid <=
      ~_GEN_2424 & _GEN_2338 & _GEN_2290
      & (_GEN_2205 ? ~_GEN_2145 & _GEN_1078 : ~_GEN_2218 & _GEN_1078);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1077) begin	// lsu.scala:304:5, :305:44
      ldq_13_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_13_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_13_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_13_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_13_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_13_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_13_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_13_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_13_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_990) begin	// lsu.scala:304:5, :306:44
      ldq_13_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_13_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_13_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_13_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_13_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_13_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_13_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_868) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_13_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_13_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_13_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_13_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_13_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_13_valid)	// lsu.scala:210:16
      ldq_13_bits_uop_br_mask <=
        ldq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1077)	// lsu.scala:304:5, :305:44
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_990)	// lsu.scala:304:5, :306:44
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_868)	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1269) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_13_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_13_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_13_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_13_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_13_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_13_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_13_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_13_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_13_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_13_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_13_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1077)	// lsu.scala:304:5, :305:44
      ldq_13_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_990)	// lsu.scala:304:5, :306:44
      ldq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_868)	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1112)	// lsu.scala:210:16, :304:5, :306:44
      ldq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_13_bits_uop_ppred_busy <= ~_GEN_1112 & ldq_13_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_13_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hD
      | (_GEN_1077
           ? io_core_dis_uops_2_bits_exception
           : _GEN_990
               ? io_core_dis_uops_1_bits_exception
               : _GEN_868
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_13_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_13_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2338 & _GEN_2290
      & (_GEN_2205 ? ~_GEN_2145 & _GEN_1270 : ~_GEN_2218 & _GEN_1270);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_13_bits_executed <=
      ~_GEN_2424 & _GEN_2338 & _GEN_2290 & _GEN_2242
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_774))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1401 & _GEN_2046 : ~(_GEN_757 & _GEN_1401) & _GEN_2046)
            : _GEN_2046) | ~_GEN_1077
         & (dis_ld_val_1
              ? ~_GEN_956 & ldq_13_bits_executed
              : ~_GEN_868 & ldq_13_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_13_bits_succeeded <=
      _GEN_2338 & _GEN_2290 & _GEN_2242
      & (_GEN_2087
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'hD
                ? _ldq_bits_succeeded_T
                : ~_GEN_1077
                  & (dis_ld_val_1
                       ? ~_GEN_956 & ldq_13_bits_succeeded
                       : ~_GEN_868 & ldq_13_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_13_bits_order_fail <=
      _GEN_2338 & _GEN_2290 & _GEN_2242
      & (_GEN_470
           ? _GEN_1136
           : _GEN_474
               ? _GEN_1436 | _GEN_1136
               : _GEN_475 & searcher_is_older_13 & _GEN_1437 | _GEN_1136);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_13_bits_observed <=
      _GEN_470 | ~_GEN_1077
      & (dis_ld_val_1
           ? ~_GEN_956 & ldq_13_bits_observed
           : ~_GEN_868 & ldq_13_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_13_bits_forward_std_val <=
      _GEN_2338 & _GEN_2290 & _GEN_2242
      & (~_GEN_787 & _GEN_2086 | ~_GEN_1077
         & (dis_ld_val_1
              ? ~_GEN_956 & ldq_13_bits_forward_std_val
              : ~_GEN_868 & ldq_13_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2087) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_13_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_14_valid <=
      ~_GEN_2424 & _GEN_2339 & _GEN_2291
      & (_GEN_2205 ? ~_GEN_2146 & _GEN_1080 : ~_GEN_2219 & _GEN_1080);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1079) begin	// lsu.scala:304:5, :305:44
      ldq_14_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_14_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_14_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_14_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_14_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_14_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_14_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_14_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_14_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_991) begin	// lsu.scala:304:5, :306:44
      ldq_14_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_14_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_14_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_14_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_14_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_14_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_14_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_869) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_14_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_14_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_14_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_14_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_14_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_14_valid)	// lsu.scala:210:16
      ldq_14_bits_uop_br_mask <=
        ldq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1079)	// lsu.scala:304:5, :305:44
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_991)	// lsu.scala:304:5, :306:44
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_869)	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1271) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_14_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_14_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_14_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_14_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_14_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_14_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_14_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_14_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_14_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_14_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_14_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1079)	// lsu.scala:304:5, :305:44
      ldq_14_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_991)	// lsu.scala:304:5, :306:44
      ldq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_869)	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1113)	// lsu.scala:210:16, :304:5, :306:44
      ldq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_14_bits_uop_ppred_busy <= ~_GEN_1113 & ldq_14_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_14_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hE
      | (_GEN_1079
           ? io_core_dis_uops_2_bits_exception
           : _GEN_991
               ? io_core_dis_uops_1_bits_exception
               : _GEN_869
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_14_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_14_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2339 & _GEN_2291
      & (_GEN_2205 ? ~_GEN_2146 & _GEN_1272 : ~_GEN_2219 & _GEN_1272);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_14_bits_executed <=
      ~_GEN_2424 & _GEN_2339 & _GEN_2291 & _GEN_2243
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_775))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1402 & _GEN_2047 : ~(_GEN_757 & _GEN_1402) & _GEN_2047)
            : _GEN_2047) | ~_GEN_1079
         & (dis_ld_val_1
              ? ~_GEN_958 & ldq_14_bits_executed
              : ~_GEN_869 & ldq_14_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_14_bits_succeeded <=
      _GEN_2339 & _GEN_2291 & _GEN_2243
      & (_GEN_2089
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'hE
                ? _ldq_bits_succeeded_T
                : ~_GEN_1079
                  & (dis_ld_val_1
                       ? ~_GEN_958 & ldq_14_bits_succeeded
                       : ~_GEN_869 & ldq_14_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_14_bits_order_fail <=
      _GEN_2339 & _GEN_2291 & _GEN_2243
      & (_GEN_481
           ? _GEN_1137
           : _GEN_485
               ? _GEN_1438 | _GEN_1137
               : _GEN_486 & searcher_is_older_14 & _GEN_1439 | _GEN_1137);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_14_bits_observed <=
      _GEN_481 | ~_GEN_1079
      & (dis_ld_val_1
           ? ~_GEN_958 & ldq_14_bits_observed
           : ~_GEN_869 & ldq_14_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_14_bits_forward_std_val <=
      _GEN_2339 & _GEN_2291 & _GEN_2243
      & (~_GEN_787 & _GEN_2088 | ~_GEN_1079
         & (dis_ld_val_1
              ? ~_GEN_958 & ldq_14_bits_forward_std_val
              : ~_GEN_869 & ldq_14_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2089) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_14_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_15_valid <=
      ~_GEN_2424 & _GEN_2340 & _GEN_2292
      & (_GEN_2205 ? ~_GEN_2147 & _GEN_1082 : ~_GEN_2220 & _GEN_1082);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1081) begin	// lsu.scala:304:5, :305:44
      ldq_15_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_15_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_15_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_15_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_15_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_15_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_15_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_15_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_15_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_992) begin	// lsu.scala:304:5, :306:44
      ldq_15_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_15_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_15_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_15_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_15_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_15_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_15_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_870) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_15_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_15_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_15_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_15_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_15_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_15_valid)	// lsu.scala:210:16
      ldq_15_bits_uop_br_mask <=
        ldq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1081)	// lsu.scala:304:5, :305:44
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_992)	// lsu.scala:304:5, :306:44
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_870)	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1273) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_15_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_15_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_15_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_15_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_15_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_15_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_15_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_15_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_15_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_15_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_15_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1081)	// lsu.scala:304:5, :305:44
      ldq_15_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_992)	// lsu.scala:304:5, :306:44
      ldq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_870)	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1114)	// lsu.scala:210:16, :304:5, :306:44
      ldq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_15_bits_uop_ppred_busy <= ~_GEN_1114 & ldq_15_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_15_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hF
      | (_GEN_1081
           ? io_core_dis_uops_2_bits_exception
           : _GEN_992
               ? io_core_dis_uops_1_bits_exception
               : _GEN_870
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_15_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_15_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2340 & _GEN_2292
      & (_GEN_2205 ? ~_GEN_2147 & _GEN_1274 : ~_GEN_2220 & _GEN_1274);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_15_bits_executed <=
      ~_GEN_2424 & _GEN_2340 & _GEN_2292 & _GEN_2244
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_776))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1403 & _GEN_2048 : ~(_GEN_757 & _GEN_1403) & _GEN_2048)
            : _GEN_2048) | ~_GEN_1081
         & (dis_ld_val_1
              ? ~_GEN_960 & ldq_15_bits_executed
              : ~_GEN_870 & ldq_15_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_15_bits_succeeded <=
      _GEN_2340 & _GEN_2292 & _GEN_2244
      & (_GEN_2091
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'hF
                ? _ldq_bits_succeeded_T
                : ~_GEN_1081
                  & (dis_ld_val_1
                       ? ~_GEN_960 & ldq_15_bits_succeeded
                       : ~_GEN_870 & ldq_15_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_15_bits_order_fail <=
      _GEN_2340 & _GEN_2292 & _GEN_2244
      & (_GEN_492
           ? _GEN_1138
           : _GEN_496
               ? _GEN_1440 | _GEN_1138
               : _GEN_497 & searcher_is_older_15 & _GEN_1441 | _GEN_1138);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_15_bits_observed <=
      _GEN_492 | ~_GEN_1081
      & (dis_ld_val_1
           ? ~_GEN_960 & ldq_15_bits_observed
           : ~_GEN_870 & ldq_15_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_15_bits_forward_std_val <=
      _GEN_2340 & _GEN_2292 & _GEN_2244
      & (~_GEN_787 & _GEN_2090 | ~_GEN_1081
         & (dis_ld_val_1
              ? ~_GEN_960 & ldq_15_bits_forward_std_val
              : ~_GEN_870 & ldq_15_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2091) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_15_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_16_valid <=
      ~_GEN_2424 & _GEN_2341 & _GEN_2293
      & (_GEN_2205 ? ~_GEN_2148 & _GEN_1084 : ~_GEN_2221 & _GEN_1084);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1083) begin	// lsu.scala:304:5, :305:44
      ldq_16_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_16_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_16_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_16_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_16_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_16_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_16_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_16_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_16_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_16_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_16_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_16_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_16_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_16_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_16_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_16_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_16_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_16_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_16_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_16_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_16_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_16_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_16_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_16_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_16_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_16_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_16_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_16_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_16_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_16_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_16_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_993) begin	// lsu.scala:304:5, :306:44
      ldq_16_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_16_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_16_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_16_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_16_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_16_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_16_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_16_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_16_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_16_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_16_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_16_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_16_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_16_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_16_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_16_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_16_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_16_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_16_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_16_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_16_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_16_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_16_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_16_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_16_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_16_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_16_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_16_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_16_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_871) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_16_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_16_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_16_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_16_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_16_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_16_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_16_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_16_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_16_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_16_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_16_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_16_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_16_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_16_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_16_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_16_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_16_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_16_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_16_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_16_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_16_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_16_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_16_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_16_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_16_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_16_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_16_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_16_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_16_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_16_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_16_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_16_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_16_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_16_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_16_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_16_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_16_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_16_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_16_valid)	// lsu.scala:210:16
      ldq_16_bits_uop_br_mask <=
        ldq_16_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1083)	// lsu.scala:304:5, :305:44
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_993)	// lsu.scala:304:5, :306:44
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_871)	// lsu.scala:210:16, :304:5, :305:44
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1275) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_16_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_16_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_16_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_16_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_16_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_16_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_16_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_16_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_16_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_16_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_16_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_16_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_16_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1083)	// lsu.scala:304:5, :305:44
      ldq_16_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_993)	// lsu.scala:304:5, :306:44
      ldq_16_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_871)	// lsu.scala:210:16, :304:5, :305:44
      ldq_16_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1115)	// lsu.scala:210:16, :304:5, :306:44
      ldq_16_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_16_bits_uop_ppred_busy <= ~_GEN_1115 & ldq_16_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_16_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h10
      | (_GEN_1083
           ? io_core_dis_uops_2_bits_exception
           : _GEN_993
               ? io_core_dis_uops_1_bits_exception
               : _GEN_871
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_16_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_16_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2341 & _GEN_2293
      & (_GEN_2205 ? ~_GEN_2148 & _GEN_1276 : ~_GEN_2221 & _GEN_1276);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_16_bits_executed <=
      ~_GEN_2424 & _GEN_2341 & _GEN_2293 & _GEN_2245
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_777))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1404 & _GEN_2049 : ~(_GEN_757 & _GEN_1404) & _GEN_2049)
            : _GEN_2049) | ~_GEN_1083
         & (dis_ld_val_1
              ? ~_GEN_962 & ldq_16_bits_executed
              : ~_GEN_871 & ldq_16_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_16_bits_succeeded <=
      _GEN_2341 & _GEN_2293 & _GEN_2245
      & (_GEN_2093
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h10
                ? _ldq_bits_succeeded_T
                : ~_GEN_1083
                  & (dis_ld_val_1
                       ? ~_GEN_962 & ldq_16_bits_succeeded
                       : ~_GEN_871 & ldq_16_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_16_bits_order_fail <=
      _GEN_2341 & _GEN_2293 & _GEN_2245
      & (_GEN_503
           ? _GEN_1139
           : _GEN_507
               ? _GEN_1442 | _GEN_1139
               : _GEN_508 & searcher_is_older_16 & _GEN_1443 | _GEN_1139);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_16_bits_observed <=
      _GEN_503 | ~_GEN_1083
      & (dis_ld_val_1
           ? ~_GEN_962 & ldq_16_bits_observed
           : ~_GEN_871 & ldq_16_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_16_bits_forward_std_val <=
      _GEN_2341 & _GEN_2293 & _GEN_2245
      & (~_GEN_787 & _GEN_2092 | ~_GEN_1083
         & (dis_ld_val_1
              ? ~_GEN_962 & ldq_16_bits_forward_std_val
              : ~_GEN_871 & ldq_16_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2093) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_16_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_17_valid <=
      ~_GEN_2424 & _GEN_2342 & _GEN_2294
      & (_GEN_2205 ? ~_GEN_2149 & _GEN_1086 : ~_GEN_2222 & _GEN_1086);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1085) begin	// lsu.scala:304:5, :305:44
      ldq_17_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_17_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_17_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_17_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_17_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_17_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_17_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_17_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_17_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_17_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_17_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_17_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_17_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_17_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_17_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_17_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_17_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_17_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_17_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_17_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_17_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_17_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_17_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_17_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_17_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_17_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_17_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_17_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_17_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_17_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_17_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_994) begin	// lsu.scala:304:5, :306:44
      ldq_17_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_17_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_17_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_17_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_17_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_17_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_17_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_17_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_17_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_17_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_17_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_17_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_17_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_17_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_17_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_17_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_17_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_17_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_17_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_17_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_17_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_17_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_17_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_17_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_17_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_17_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_17_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_17_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_17_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_872) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_17_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_17_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_17_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_17_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_17_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_17_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_17_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_17_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_17_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_17_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_17_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_17_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_17_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_17_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_17_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_17_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_17_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_17_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_17_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_17_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_17_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_17_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_17_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_17_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_17_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_17_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_17_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_17_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_17_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_17_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_17_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_17_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_17_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_17_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_17_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_17_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_17_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_17_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_17_valid)	// lsu.scala:210:16
      ldq_17_bits_uop_br_mask <=
        ldq_17_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1085)	// lsu.scala:304:5, :305:44
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_994)	// lsu.scala:304:5, :306:44
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_872)	// lsu.scala:210:16, :304:5, :305:44
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1277) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_17_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_17_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_17_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_17_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_17_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_17_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_17_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_17_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_17_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_17_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_17_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_17_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_17_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1085)	// lsu.scala:304:5, :305:44
      ldq_17_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_994)	// lsu.scala:304:5, :306:44
      ldq_17_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_872)	// lsu.scala:210:16, :304:5, :305:44
      ldq_17_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1116)	// lsu.scala:210:16, :304:5, :306:44
      ldq_17_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_17_bits_uop_ppred_busy <= ~_GEN_1116 & ldq_17_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_17_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h11
      | (_GEN_1085
           ? io_core_dis_uops_2_bits_exception
           : _GEN_994
               ? io_core_dis_uops_1_bits_exception
               : _GEN_872
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_17_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_17_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2342 & _GEN_2294
      & (_GEN_2205 ? ~_GEN_2149 & _GEN_1278 : ~_GEN_2222 & _GEN_1278);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_17_bits_executed <=
      ~_GEN_2424 & _GEN_2342 & _GEN_2294 & _GEN_2246
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_778))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1405 & _GEN_2050 : ~(_GEN_757 & _GEN_1405) & _GEN_2050)
            : _GEN_2050) | ~_GEN_1085
         & (dis_ld_val_1
              ? ~_GEN_964 & ldq_17_bits_executed
              : ~_GEN_872 & ldq_17_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_17_bits_succeeded <=
      _GEN_2342 & _GEN_2294 & _GEN_2246
      & (_GEN_2095
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h11
                ? _ldq_bits_succeeded_T
                : ~_GEN_1085
                  & (dis_ld_val_1
                       ? ~_GEN_964 & ldq_17_bits_succeeded
                       : ~_GEN_872 & ldq_17_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_17_bits_order_fail <=
      _GEN_2342 & _GEN_2294 & _GEN_2246
      & (_GEN_514
           ? _GEN_1140
           : _GEN_518
               ? _GEN_1444 | _GEN_1140
               : _GEN_519 & searcher_is_older_17 & _GEN_1445 | _GEN_1140);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_17_bits_observed <=
      _GEN_514 | ~_GEN_1085
      & (dis_ld_val_1
           ? ~_GEN_964 & ldq_17_bits_observed
           : ~_GEN_872 & ldq_17_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_17_bits_forward_std_val <=
      _GEN_2342 & _GEN_2294 & _GEN_2246
      & (~_GEN_787 & _GEN_2094 | ~_GEN_1085
         & (dis_ld_val_1
              ? ~_GEN_964 & ldq_17_bits_forward_std_val
              : ~_GEN_872 & ldq_17_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2095) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_17_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_18_valid <=
      ~_GEN_2424 & _GEN_2343 & _GEN_2295
      & (_GEN_2205 ? ~_GEN_2150 & _GEN_1088 : ~_GEN_2223 & _GEN_1088);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1087) begin	// lsu.scala:304:5, :305:44
      ldq_18_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_18_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_18_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_18_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_18_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_18_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_18_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_18_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_18_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_18_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_18_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_18_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_18_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_18_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_18_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_18_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_18_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_18_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_18_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_18_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_18_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_18_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_18_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_18_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_18_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_18_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_18_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_18_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_18_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_18_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_18_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_995) begin	// lsu.scala:304:5, :306:44
      ldq_18_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_18_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_18_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_18_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_18_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_18_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_18_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_18_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_18_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_18_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_18_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_18_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_18_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_18_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_18_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_18_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_18_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_18_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_18_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_18_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_18_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_18_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_18_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_18_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_18_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_18_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_18_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_18_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_18_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_873) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_18_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_18_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_18_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_18_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_18_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_18_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_18_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_18_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_18_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_18_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_18_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_18_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_18_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_18_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_18_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_18_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_18_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_18_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_18_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_18_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_18_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_18_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_18_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_18_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_18_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_18_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_18_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_18_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_18_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_18_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_18_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_18_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_18_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_18_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_18_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_18_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_18_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_18_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_18_valid)	// lsu.scala:210:16
      ldq_18_bits_uop_br_mask <=
        ldq_18_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1087)	// lsu.scala:304:5, :305:44
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_995)	// lsu.scala:304:5, :306:44
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_873)	// lsu.scala:210:16, :304:5, :305:44
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1279) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_18_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_18_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_18_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_18_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_18_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_18_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_18_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_18_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_18_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_18_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_18_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_18_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_18_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1087)	// lsu.scala:304:5, :305:44
      ldq_18_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_995)	// lsu.scala:304:5, :306:44
      ldq_18_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_873)	// lsu.scala:210:16, :304:5, :305:44
      ldq_18_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1117)	// lsu.scala:210:16, :304:5, :306:44
      ldq_18_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_18_bits_uop_ppred_busy <= ~_GEN_1117 & ldq_18_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_18_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h12
      | (_GEN_1087
           ? io_core_dis_uops_2_bits_exception
           : _GEN_995
               ? io_core_dis_uops_1_bits_exception
               : _GEN_873
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_18_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_18_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2343 & _GEN_2295
      & (_GEN_2205 ? ~_GEN_2150 & _GEN_1280 : ~_GEN_2223 & _GEN_1280);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_18_bits_executed <=
      ~_GEN_2424 & _GEN_2343 & _GEN_2295 & _GEN_2247
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_779))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1406 & _GEN_2051 : ~(_GEN_757 & _GEN_1406) & _GEN_2051)
            : _GEN_2051) | ~_GEN_1087
         & (dis_ld_val_1
              ? ~_GEN_966 & ldq_18_bits_executed
              : ~_GEN_873 & ldq_18_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_18_bits_succeeded <=
      _GEN_2343 & _GEN_2295 & _GEN_2247
      & (_GEN_2097
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h12
                ? _ldq_bits_succeeded_T
                : ~_GEN_1087
                  & (dis_ld_val_1
                       ? ~_GEN_966 & ldq_18_bits_succeeded
                       : ~_GEN_873 & ldq_18_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_18_bits_order_fail <=
      _GEN_2343 & _GEN_2295 & _GEN_2247
      & (_GEN_525
           ? _GEN_1141
           : _GEN_529
               ? _GEN_1446 | _GEN_1141
               : _GEN_530 & searcher_is_older_18 & _GEN_1447 | _GEN_1141);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_18_bits_observed <=
      _GEN_525 | ~_GEN_1087
      & (dis_ld_val_1
           ? ~_GEN_966 & ldq_18_bits_observed
           : ~_GEN_873 & ldq_18_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_18_bits_forward_std_val <=
      _GEN_2343 & _GEN_2295 & _GEN_2247
      & (~_GEN_787 & _GEN_2096 | ~_GEN_1087
         & (dis_ld_val_1
              ? ~_GEN_966 & ldq_18_bits_forward_std_val
              : ~_GEN_873 & ldq_18_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2097) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_18_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_19_valid <=
      ~_GEN_2424 & _GEN_2344 & _GEN_2296
      & (_GEN_2205 ? ~_GEN_2151 & _GEN_1090 : ~_GEN_2224 & _GEN_1090);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1089) begin	// lsu.scala:304:5, :305:44
      ldq_19_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_19_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_19_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_19_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_19_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_19_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_19_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_19_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_19_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_19_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_19_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_19_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_19_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_19_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_19_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_19_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_19_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_19_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_19_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_19_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_19_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_19_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_19_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_19_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_19_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_19_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_19_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_19_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_19_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_19_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_19_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_996) begin	// lsu.scala:304:5, :306:44
      ldq_19_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_19_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_19_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_19_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_19_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_19_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_19_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_19_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_19_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_19_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_19_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_19_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_19_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_19_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_19_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_19_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_19_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_19_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_19_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_19_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_19_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_19_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_19_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_19_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_19_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_19_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_19_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_19_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_19_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_874) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_19_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_19_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_19_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_19_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_19_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_19_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_19_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_19_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_19_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_19_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_19_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_19_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_19_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_19_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_19_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_19_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_19_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_19_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_19_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_19_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_19_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_19_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_19_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_19_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_19_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_19_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_19_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_19_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_19_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_19_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_19_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_19_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_19_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_19_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_19_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_19_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_19_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_19_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_19_valid)	// lsu.scala:210:16
      ldq_19_bits_uop_br_mask <=
        ldq_19_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1089)	// lsu.scala:304:5, :305:44
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_996)	// lsu.scala:304:5, :306:44
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_874)	// lsu.scala:210:16, :304:5, :305:44
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1281) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_19_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_19_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_19_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_19_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_19_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_19_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_19_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_19_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_19_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_19_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_19_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_19_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_19_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1089)	// lsu.scala:304:5, :305:44
      ldq_19_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_996)	// lsu.scala:304:5, :306:44
      ldq_19_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_874)	// lsu.scala:210:16, :304:5, :305:44
      ldq_19_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1118)	// lsu.scala:210:16, :304:5, :306:44
      ldq_19_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_19_bits_uop_ppred_busy <= ~_GEN_1118 & ldq_19_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_19_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h13
      | (_GEN_1089
           ? io_core_dis_uops_2_bits_exception
           : _GEN_996
               ? io_core_dis_uops_1_bits_exception
               : _GEN_874
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_19_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_19_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2344 & _GEN_2296
      & (_GEN_2205 ? ~_GEN_2151 & _GEN_1282 : ~_GEN_2224 & _GEN_1282);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_19_bits_executed <=
      ~_GEN_2424 & _GEN_2344 & _GEN_2296 & _GEN_2248
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_780))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1407 & _GEN_2052 : ~(_GEN_757 & _GEN_1407) & _GEN_2052)
            : _GEN_2052) | ~_GEN_1089
         & (dis_ld_val_1
              ? ~_GEN_968 & ldq_19_bits_executed
              : ~_GEN_874 & ldq_19_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_19_bits_succeeded <=
      _GEN_2344 & _GEN_2296 & _GEN_2248
      & (_GEN_2099
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h13
                ? _ldq_bits_succeeded_T
                : ~_GEN_1089
                  & (dis_ld_val_1
                       ? ~_GEN_968 & ldq_19_bits_succeeded
                       : ~_GEN_874 & ldq_19_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_19_bits_order_fail <=
      _GEN_2344 & _GEN_2296 & _GEN_2248
      & (_GEN_536
           ? _GEN_1142
           : _GEN_540
               ? _GEN_1448 | _GEN_1142
               : _GEN_541 & searcher_is_older_19 & _GEN_1449 | _GEN_1142);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_19_bits_observed <=
      _GEN_536 | ~_GEN_1089
      & (dis_ld_val_1
           ? ~_GEN_968 & ldq_19_bits_observed
           : ~_GEN_874 & ldq_19_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_19_bits_forward_std_val <=
      _GEN_2344 & _GEN_2296 & _GEN_2248
      & (~_GEN_787 & _GEN_2098 | ~_GEN_1089
         & (dis_ld_val_1
              ? ~_GEN_968 & ldq_19_bits_forward_std_val
              : ~_GEN_874 & ldq_19_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2099) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_19_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_20_valid <=
      ~_GEN_2424 & _GEN_2345 & _GEN_2297
      & (_GEN_2205 ? ~_GEN_2152 & _GEN_1092 : ~_GEN_2225 & _GEN_1092);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1091) begin	// lsu.scala:304:5, :305:44
      ldq_20_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_20_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_20_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_20_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_20_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_20_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_20_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_20_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_20_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_20_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_20_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_20_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_20_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_20_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_20_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_20_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_20_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_20_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_20_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_20_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_20_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_20_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_20_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_20_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_20_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_20_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_20_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_20_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_20_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_20_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_20_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_997) begin	// lsu.scala:304:5, :306:44
      ldq_20_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_20_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_20_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_20_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_20_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_20_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_20_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_20_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_20_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_20_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_20_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_20_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_20_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_20_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_20_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_20_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_20_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_20_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_20_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_20_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_20_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_20_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_20_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_20_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_20_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_20_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_20_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_20_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_20_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_875) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_20_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_20_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_20_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_20_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_20_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_20_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_20_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_20_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_20_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_20_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_20_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_20_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_20_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_20_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_20_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_20_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_20_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_20_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_20_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_20_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_20_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_20_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_20_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_20_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_20_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_20_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_20_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_20_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_20_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_20_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_20_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_20_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_20_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_20_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_20_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_20_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_20_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_20_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_20_valid)	// lsu.scala:210:16
      ldq_20_bits_uop_br_mask <=
        ldq_20_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1091)	// lsu.scala:304:5, :305:44
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_997)	// lsu.scala:304:5, :306:44
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_875)	// lsu.scala:210:16, :304:5, :305:44
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1283) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_20_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_20_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_20_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_20_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_20_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_20_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_20_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_20_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_20_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_20_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_20_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_20_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_20_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1091)	// lsu.scala:304:5, :305:44
      ldq_20_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_997)	// lsu.scala:304:5, :306:44
      ldq_20_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_875)	// lsu.scala:210:16, :304:5, :305:44
      ldq_20_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1119)	// lsu.scala:210:16, :304:5, :306:44
      ldq_20_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_20_bits_uop_ppred_busy <= ~_GEN_1119 & ldq_20_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_20_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h14
      | (_GEN_1091
           ? io_core_dis_uops_2_bits_exception
           : _GEN_997
               ? io_core_dis_uops_1_bits_exception
               : _GEN_875
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_20_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_20_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2345 & _GEN_2297
      & (_GEN_2205 ? ~_GEN_2152 & _GEN_1284 : ~_GEN_2225 & _GEN_1284);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_20_bits_executed <=
      ~_GEN_2424 & _GEN_2345 & _GEN_2297 & _GEN_2249
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_781))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1408 & _GEN_2053 : ~(_GEN_757 & _GEN_1408) & _GEN_2053)
            : _GEN_2053) | ~_GEN_1091
         & (dis_ld_val_1
              ? ~_GEN_970 & ldq_20_bits_executed
              : ~_GEN_875 & ldq_20_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_20_bits_succeeded <=
      _GEN_2345 & _GEN_2297 & _GEN_2249
      & (_GEN_2101
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h14
                ? _ldq_bits_succeeded_T
                : ~_GEN_1091
                  & (dis_ld_val_1
                       ? ~_GEN_970 & ldq_20_bits_succeeded
                       : ~_GEN_875 & ldq_20_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_20_bits_order_fail <=
      _GEN_2345 & _GEN_2297 & _GEN_2249
      & (_GEN_547
           ? _GEN_1143
           : _GEN_551
               ? _GEN_1450 | _GEN_1143
               : _GEN_552 & searcher_is_older_20 & _GEN_1451 | _GEN_1143);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_20_bits_observed <=
      _GEN_547 | ~_GEN_1091
      & (dis_ld_val_1
           ? ~_GEN_970 & ldq_20_bits_observed
           : ~_GEN_875 & ldq_20_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_20_bits_forward_std_val <=
      _GEN_2345 & _GEN_2297 & _GEN_2249
      & (~_GEN_787 & _GEN_2100 | ~_GEN_1091
         & (dis_ld_val_1
              ? ~_GEN_970 & ldq_20_bits_forward_std_val
              : ~_GEN_875 & ldq_20_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2101) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_20_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_21_valid <=
      ~_GEN_2424 & _GEN_2346 & _GEN_2298
      & (_GEN_2205 ? ~_GEN_2153 & _GEN_1094 : ~_GEN_2226 & _GEN_1094);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1093) begin	// lsu.scala:304:5, :305:44
      ldq_21_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_21_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_21_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_21_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_21_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_21_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_21_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_21_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_21_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_21_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_21_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_21_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_21_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_21_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_21_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_21_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_21_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_21_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_21_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_21_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_21_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_21_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_21_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_21_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_21_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_21_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_21_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_21_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_21_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_21_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_21_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_998) begin	// lsu.scala:304:5, :306:44
      ldq_21_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_21_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_21_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_21_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_21_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_21_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_21_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_21_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_21_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_21_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_21_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_21_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_21_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_21_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_21_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_21_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_21_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_21_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_21_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_21_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_21_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_21_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_21_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_21_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_21_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_21_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_21_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_21_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_21_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_876) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_21_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_21_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_21_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_21_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_21_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_21_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_21_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_21_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_21_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_21_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_21_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_21_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_21_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_21_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_21_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_21_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_21_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_21_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_21_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_21_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_21_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_21_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_21_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_21_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_21_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_21_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_21_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_21_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_21_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_21_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_21_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_21_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_21_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_21_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_21_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_21_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_21_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_21_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_21_valid)	// lsu.scala:210:16
      ldq_21_bits_uop_br_mask <=
        ldq_21_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1093)	// lsu.scala:304:5, :305:44
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_998)	// lsu.scala:304:5, :306:44
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_876)	// lsu.scala:210:16, :304:5, :305:44
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1285) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_21_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_21_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_21_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_21_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_21_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_21_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_21_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_21_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_21_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_21_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_21_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_21_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_21_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1093)	// lsu.scala:304:5, :305:44
      ldq_21_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_998)	// lsu.scala:304:5, :306:44
      ldq_21_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_876)	// lsu.scala:210:16, :304:5, :305:44
      ldq_21_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1120)	// lsu.scala:210:16, :304:5, :306:44
      ldq_21_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_21_bits_uop_ppred_busy <= ~_GEN_1120 & ldq_21_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_21_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h15
      | (_GEN_1093
           ? io_core_dis_uops_2_bits_exception
           : _GEN_998
               ? io_core_dis_uops_1_bits_exception
               : _GEN_876
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_21_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_21_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2346 & _GEN_2298
      & (_GEN_2205 ? ~_GEN_2153 & _GEN_1286 : ~_GEN_2226 & _GEN_1286);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_21_bits_executed <=
      ~_GEN_2424 & _GEN_2346 & _GEN_2298 & _GEN_2250
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_782))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1409 & _GEN_2054 : ~(_GEN_757 & _GEN_1409) & _GEN_2054)
            : _GEN_2054) | ~_GEN_1093
         & (dis_ld_val_1
              ? ~_GEN_972 & ldq_21_bits_executed
              : ~_GEN_876 & ldq_21_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_21_bits_succeeded <=
      _GEN_2346 & _GEN_2298 & _GEN_2250
      & (_GEN_2103
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h15
                ? _ldq_bits_succeeded_T
                : ~_GEN_1093
                  & (dis_ld_val_1
                       ? ~_GEN_972 & ldq_21_bits_succeeded
                       : ~_GEN_876 & ldq_21_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_21_bits_order_fail <=
      _GEN_2346 & _GEN_2298 & _GEN_2250
      & (_GEN_558
           ? _GEN_1144
           : _GEN_562
               ? _GEN_1452 | _GEN_1144
               : _GEN_563 & searcher_is_older_21 & _GEN_1453 | _GEN_1144);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_21_bits_observed <=
      _GEN_558 | ~_GEN_1093
      & (dis_ld_val_1
           ? ~_GEN_972 & ldq_21_bits_observed
           : ~_GEN_876 & ldq_21_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_21_bits_forward_std_val <=
      _GEN_2346 & _GEN_2298 & _GEN_2250
      & (~_GEN_787 & _GEN_2102 | ~_GEN_1093
         & (dis_ld_val_1
              ? ~_GEN_972 & ldq_21_bits_forward_std_val
              : ~_GEN_876 & ldq_21_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2103) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_21_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_22_valid <=
      ~_GEN_2424 & _GEN_2347 & _GEN_2299
      & (_GEN_2205 ? ~_GEN_2154 & _GEN_1096 : ~_GEN_2227 & _GEN_1096);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1095) begin	// lsu.scala:304:5, :305:44
      ldq_22_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_22_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_22_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_22_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_22_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_22_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_22_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_22_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_22_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_22_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_22_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_22_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_22_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_22_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_22_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_22_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_22_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_22_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_22_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_22_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_22_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_22_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_22_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_22_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_22_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_22_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_22_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_22_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_22_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_22_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_22_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_999) begin	// lsu.scala:304:5, :306:44
      ldq_22_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_22_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_22_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_22_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_22_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_22_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_22_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_22_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_22_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_22_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_22_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_22_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_22_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_22_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_22_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_22_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_22_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_22_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_22_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_22_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_22_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_22_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_22_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_22_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_22_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_22_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_22_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_22_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_22_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_877) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_22_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_22_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_22_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_22_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_22_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_22_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_22_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_22_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_22_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_22_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_22_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_22_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_22_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_22_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_22_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_22_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_22_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_22_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_22_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_22_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_22_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_22_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_22_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_22_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_22_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_22_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_22_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_22_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_22_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_22_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_22_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_22_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_22_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_22_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_22_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_22_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_22_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_22_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_22_valid)	// lsu.scala:210:16
      ldq_22_bits_uop_br_mask <=
        ldq_22_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1095)	// lsu.scala:304:5, :305:44
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_999)	// lsu.scala:304:5, :306:44
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_877)	// lsu.scala:210:16, :304:5, :305:44
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1287) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_22_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_22_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_22_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_22_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_22_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_22_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_22_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_22_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_22_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_22_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_22_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_22_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_22_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1095)	// lsu.scala:304:5, :305:44
      ldq_22_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_999)	// lsu.scala:304:5, :306:44
      ldq_22_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_877)	// lsu.scala:210:16, :304:5, :305:44
      ldq_22_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1121)	// lsu.scala:210:16, :304:5, :306:44
      ldq_22_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_22_bits_uop_ppred_busy <= ~_GEN_1121 & ldq_22_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_22_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h16
      | (_GEN_1095
           ? io_core_dis_uops_2_bits_exception
           : _GEN_999
               ? io_core_dis_uops_1_bits_exception
               : _GEN_877
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_22_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_22_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2347 & _GEN_2299
      & (_GEN_2205 ? ~_GEN_2154 & _GEN_1288 : ~_GEN_2227 & _GEN_1288);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_22_bits_executed <=
      ~_GEN_2424 & _GEN_2347 & _GEN_2299 & _GEN_2251
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_783))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1410 & _GEN_2055 : ~(_GEN_757 & _GEN_1410) & _GEN_2055)
            : _GEN_2055) | ~_GEN_1095
         & (dis_ld_val_1
              ? ~_GEN_974 & ldq_22_bits_executed
              : ~_GEN_877 & ldq_22_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_22_bits_succeeded <=
      _GEN_2347 & _GEN_2299 & _GEN_2251
      & (_GEN_2105
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h16
                ? _ldq_bits_succeeded_T
                : ~_GEN_1095
                  & (dis_ld_val_1
                       ? ~_GEN_974 & ldq_22_bits_succeeded
                       : ~_GEN_877 & ldq_22_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_22_bits_order_fail <=
      _GEN_2347 & _GEN_2299 & _GEN_2251
      & (_GEN_569
           ? _GEN_1145
           : _GEN_573
               ? _GEN_1454 | _GEN_1145
               : _GEN_574 & searcher_is_older_22 & _GEN_1455 | _GEN_1145);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_22_bits_observed <=
      _GEN_569 | ~_GEN_1095
      & (dis_ld_val_1
           ? ~_GEN_974 & ldq_22_bits_observed
           : ~_GEN_877 & ldq_22_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_22_bits_forward_std_val <=
      _GEN_2347 & _GEN_2299 & _GEN_2251
      & (~_GEN_787 & _GEN_2104 | ~_GEN_1095
         & (dis_ld_val_1
              ? ~_GEN_974 & ldq_22_bits_forward_std_val
              : ~_GEN_877 & ldq_22_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2105) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_22_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_23_valid <=
      ~_GEN_2424 & _GEN_2348 & _GEN_2300
      & (_GEN_2205 ? ~_GEN_2155 & _GEN_1098 : ~_GEN_2228 & _GEN_1098);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_1097) begin	// lsu.scala:304:5, :305:44
      ldq_23_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:210:16
      ldq_23_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:210:16
      ldq_23_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:210:16
      ldq_23_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_23_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;	// lsu.scala:210:16
      ldq_23_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;	// lsu.scala:210:16
      ldq_23_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;	// lsu.scala:210:16
      ldq_23_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;	// lsu.scala:210:16
      ldq_23_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:210:16
      ldq_23_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:210:16
      ldq_23_bits_uop_taken <= io_core_dis_uops_2_bits_taken;	// lsu.scala:210:16
      ldq_23_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:210:16
      ldq_23_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:210:16
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:210:16
      ldq_23_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:210:16
      ldq_23_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:210:16
      ldq_23_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:210:16
      ldq_23_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:210:16
      ldq_23_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;	// lsu.scala:210:16
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;	// lsu.scala:210:16
      ldq_23_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;	// lsu.scala:210:16
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;	// lsu.scala:210:16
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;	// lsu.scala:210:16
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;	// lsu.scala:210:16
      ldq_23_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_23_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;	// lsu.scala:210:16
      ldq_23_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;	// lsu.scala:210:16
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;	// lsu.scala:210:16
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;	// lsu.scala:210:16
      ldq_23_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_23_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_23_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_23_bits_st_dep_mask <= _GEN_1050;	// lsu.scala:210:16, :336:31
      if (dis_st_val_1) begin	// lsu.scala:302:85
        if (wrap_5)	// util.scala:205:25
          ldq_23_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_23_bits_youngest_stq_idx <= _GEN_104;	// lsu.scala:210:16, util.scala:206:28
      end
      else if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_23_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_23_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_23_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_1000) begin	// lsu.scala:304:5, :306:44
      ldq_23_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_23_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_23_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_23_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_23_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_23_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_23_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_23_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_23_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_23_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_23_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_23_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_23_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_23_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_23_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_23_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_23_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_23_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_23_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_23_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_23_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_23_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_23_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_23_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_23_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_23_bits_st_dep_mask <= _GEN_928;	// lsu.scala:210:16, :336:31
      if (dis_st_val) begin	// lsu.scala:302:85
        if (wrap_1)	// util.scala:205:25
          ldq_23_bits_youngest_stq_idx <= 5'h0;	// lsu.scala:210:16
        else	// util.scala:205:25
          ldq_23_bits_youngest_stq_idx <= _GEN_97;	// lsu.scala:210:16, util.scala:206:28
      end
      else	// lsu.scala:302:85
        ldq_23_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_878) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_23_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_23_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_23_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_23_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_23_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_23_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_23_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_23_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_23_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_23_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_23_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_23_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_23_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_23_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_23_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_23_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_23_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_23_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_23_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_23_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_23_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_23_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_23_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_23_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_23_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_23_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_23_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_23_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_23_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_23_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_23_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_23_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_23_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_23_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_23_bits_st_dep_mask <= _GEN_854;	// lsu.scala:210:16, :260:33
      ldq_23_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_23_bits_st_dep_mask <=
        (_GEN_853 | ~(_ldq_23_bits_st_dep_mask_T[23:0])) & ldq_23_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_23_valid)	// lsu.scala:210:16
      ldq_23_bits_uop_br_mask <=
        ldq_23_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_1097)	// lsu.scala:304:5, :305:44
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_1000)	// lsu.scala:304:5, :306:44
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_878)	// lsu.scala:210:16, :304:5, :305:44
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_1289) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_23_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_23_bits_uop_pdst <= _GEN_154;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_23_bits_uop_pdst <= _GEN_207;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_23_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_23_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_23_bits_addr_bits <= _GEN_312;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_23_bits_addr_bits <= _GEN_199;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_23_bits_addr_bits <= _GEN_208;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_23_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_23_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_23_bits_addr_bits <= _GEN_313;	// lsu.scala:210:16, :768:30
      ldq_23_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_23_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_1097)	// lsu.scala:304:5, :305:44
      ldq_23_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_1000)	// lsu.scala:304:5, :306:44
      ldq_23_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_878)	// lsu.scala:210:16, :304:5, :305:44
      ldq_23_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_1122)	// lsu.scala:210:16, :304:5, :306:44
      ldq_23_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_23_bits_uop_ppred_busy <= ~_GEN_1122 & ldq_23_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_23_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h17
      | (_GEN_1097
           ? io_core_dis_uops_2_bits_exception
           : _GEN_1000
               ? io_core_dis_uops_1_bits_exception
               : _GEN_878
                   ? io_core_dis_uops_0_bits_exception
                   : ldq_23_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58, util.scala:205:25
    ldq_23_bits_addr_valid <=
      ~_GEN_2424 & _GEN_2348 & _GEN_2300
      & (_GEN_2205 ? ~_GEN_2155 & _GEN_1290 : ~_GEN_2228 & _GEN_1290);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_23_bits_executed <=
      ~_GEN_2424 & _GEN_2348 & _GEN_2300 & _GEN_2252
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_784))
      & ((_GEN_753
            ? (_GEN_2057 ? ~_GEN_1411 & _GEN_2056 : ~(_GEN_757 & _GEN_1411) & _GEN_2056)
            : _GEN_2056) | ~_GEN_1097
         & (dis_ld_val_1
              ? ~_GEN_976 & ldq_23_bits_executed
              : ~_GEN_878 & ldq_23_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_23_bits_succeeded <=
      _GEN_2348 & _GEN_2300 & _GEN_2252
      & (_GEN_2107
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 5'h17
                ? _ldq_bits_succeeded_T
                : ~_GEN_1097
                  & (dis_ld_val_1
                       ? ~_GEN_976 & ldq_23_bits_succeeded
                       : ~_GEN_878 & ldq_23_bits_succeeded))
           : _GEN_797);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31, util.scala:205:25
    ldq_23_bits_order_fail <=
      _GEN_2348 & _GEN_2300 & _GEN_2252
      & (_GEN_580
           ? _GEN_1146
           : _GEN_584
               ? _GEN_1456 | _GEN_1146
               : _GEN_585 & searcher_is_older_23 & _GEN_1457 | _GEN_1146);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_23_bits_observed <=
      _GEN_580 | ~_GEN_1097
      & (dis_ld_val_1
           ? ~_GEN_976 & ldq_23_bits_observed
           : ~_GEN_878 & ldq_23_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_23_bits_forward_std_val <=
      _GEN_2348 & _GEN_2300 & _GEN_2252
      & (~_GEN_787 & _GEN_2106 | ~_GEN_1097
         & (dis_ld_val_1
              ? ~_GEN_976 & ldq_23_bits_forward_std_val
              : ~_GEN_878 & ldq_23_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_2107) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_23_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    stq_0_valid <=
      ~_GEN_2427 & (clear_store ? ~_GEN_2350 & _GEN_1148 : ~_GEN_2108 & _GEN_1148);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    if (_GEN_2425) begin	// lsu.scala:1505:3, :1597:3, :1602:5, :1603:16
      stq_0_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_0_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_0_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_0_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_0_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_0_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_0_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_0_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_0_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_0_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_0_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_1_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_1_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_1_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_1_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_1_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_1_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_1_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_1_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_1_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_1_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_2_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_2_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_2_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_2_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_2_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_2_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_2_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_2_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_2_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_2_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_3_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_3_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_3_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_3_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_3_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_3_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_3_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_3_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_3_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_3_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_4_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_4_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_4_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_4_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_4_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_4_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_4_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_4_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_4_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_4_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_5_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_5_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_5_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_5_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_5_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_5_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_5_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_5_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_5_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_5_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_6_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_6_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_6_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_6_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_6_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_6_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_6_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_6_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_6_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_6_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_7_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_7_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_7_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_7_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_7_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_7_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_7_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_7_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_7_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_7_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_8_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_8_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_8_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_8_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_8_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_8_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_8_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_8_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_8_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_8_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_9_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_9_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_9_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_9_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_9_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_9_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_9_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_9_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_9_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_9_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_10_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_10_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_10_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_10_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_10_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_10_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_10_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_10_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_10_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_10_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_11_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_11_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_11_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_11_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_11_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_11_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_11_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_11_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_11_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_11_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_12_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_12_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_12_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_12_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_12_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_12_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_12_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_12_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_12_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_12_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_13_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_13_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_13_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_13_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_13_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_13_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_13_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_13_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_13_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_13_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_14_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_14_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_14_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_14_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_14_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_14_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_14_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_14_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_14_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_14_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_15_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_15_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_15_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_15_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_15_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_15_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_15_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_15_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_15_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_15_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_16_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_16_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_16_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_16_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_16_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_16_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_16_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_16_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_16_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_16_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_16_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_16_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_16_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_16_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_16_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_16_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_16_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_16_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_16_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_16_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_16_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_16_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_16_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_16_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_16_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_16_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_17_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_17_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_17_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_17_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_17_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_17_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_17_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_17_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_17_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_17_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_17_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_17_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_17_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_17_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_17_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_17_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_17_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_17_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_17_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_17_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_17_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_17_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_17_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_17_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_17_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_17_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_18_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_18_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_18_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_18_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_18_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_18_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_18_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_18_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_18_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_18_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_18_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_18_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_18_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_18_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_18_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_18_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_18_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_18_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_18_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_18_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_18_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_18_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_18_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_18_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_18_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_18_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_19_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_19_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_19_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_19_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_19_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_19_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_19_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_19_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_19_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_19_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_19_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_19_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_19_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_19_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_19_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_19_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_19_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_19_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_19_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_19_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_19_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_19_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_19_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_19_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_19_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_19_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_20_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_20_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_20_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_20_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_20_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_20_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_20_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_20_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_20_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_20_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_20_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_20_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_20_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_20_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_20_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_20_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_20_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_20_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_20_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_20_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_20_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_20_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_20_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_20_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_20_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_20_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_21_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_21_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_21_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_21_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_21_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_21_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_21_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_21_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_21_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_21_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_21_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_21_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_21_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_21_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_21_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_21_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_21_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_21_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_21_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_21_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_21_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_21_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_21_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_21_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_21_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_21_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_22_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_22_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_22_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_22_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_22_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_22_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_22_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_22_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_22_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_22_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_22_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_22_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_22_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_22_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_22_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_22_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_22_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_22_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_22_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_22_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_22_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_22_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_22_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_22_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_22_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_22_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_23_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_23_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_23_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_23_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_23_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_23_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_br_mask <= 16'h0;	// lsu.scala:211:16
      stq_23_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_23_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_23_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_23_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_23_bits_uop_rob_idx <= 7'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ldq_idx <= 5'h0;	// lsu.scala:211:16
      stq_23_bits_uop_stq_idx <= 5'h0;	// lsu.scala:211:16
      stq_23_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_23_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_23_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_23_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_23_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_23_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_23_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_23_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_23_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_23_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_23_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_23_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_23_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_23_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_head <= 5'h0;	// lsu.scala:217:29
      stq_commit_head <= 5'h0;	// lsu.scala:219:29
      stq_execute_head <= 5'h0;	// lsu.scala:220:29
    end
    else begin	// lsu.scala:1505:3, :1597:3, :1602:5, :1603:16
      if (_GEN_1195) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1025) begin	// lsu.scala:304:5, :321:5
          if (_GEN_903) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_0_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_0_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_0_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_0_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_0_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_0_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_0_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_0_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_0_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_0_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_0_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_0_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_0_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_0_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_0_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_0_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_0_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_0_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_0_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_0_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_0_valid)	// lsu.scala:211:16
        stq_0_bits_uop_br_mask <=
          stq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1195) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1025) begin	// lsu.scala:304:5, :321:5
          if (_GEN_903) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1195) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1025) begin	// lsu.scala:304:5, :321:5
          if (_GEN_903) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_0_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_0_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_0_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_0_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_0_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_0_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_0_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_0_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_0_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_0_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_0_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_0_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_0_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_0_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_0_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_0_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_0_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_0_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_0_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_0_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1291) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_0_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_0_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_0_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1195) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1025) begin	// lsu.scala:304:5, :321:5
          if (_GEN_903) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1195) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1025) begin	// lsu.scala:304:5, :321:5
          if (_GEN_903) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_0_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_0_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_0_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_0_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_0_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_0_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_0_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_0_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_0_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_0_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_0_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_0_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_0_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_0_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_0_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_0_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_0_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_0_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_0_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_0_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_0_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_0_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_0_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_0_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_0_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_0_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_0_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_0_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_0_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1196) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1026) begin	// lsu.scala:304:5, :321:5
          if (_GEN_904) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_1_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_1_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_1_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_1_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_1_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_1_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_1_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_1_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_1_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_1_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_1_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_1_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_1_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_1_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_1_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_1_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_1_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_1_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_1_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_1_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_1_valid)	// lsu.scala:211:16
        stq_1_bits_uop_br_mask <=
          stq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1196) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1026) begin	// lsu.scala:304:5, :321:5
          if (_GEN_904) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1196) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1026) begin	// lsu.scala:304:5, :321:5
          if (_GEN_904) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_1_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_1_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_1_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_1_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_1_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_1_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_1_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_1_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_1_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_1_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_1_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_1_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_1_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_1_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_1_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_1_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_1_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_1_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_1_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_1_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1293) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_1_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_1_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_1_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1196) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1026) begin	// lsu.scala:304:5, :321:5
          if (_GEN_904) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1196) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1026) begin	// lsu.scala:304:5, :321:5
          if (_GEN_904) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_1_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_1_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_1_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_1_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_1_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_1_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_1_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_1_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_1_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_1_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_1_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_1_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_1_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_1_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_1_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_1_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_1_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_1_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_1_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_1_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_1_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_1_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_1_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_1_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_1_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_1_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_1_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_1_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_1_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1197) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1027) begin	// lsu.scala:304:5, :321:5
          if (_GEN_905) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_2_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_2_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_2_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_2_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_2_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_2_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_2_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_2_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_2_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_2_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_2_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_2_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_2_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_2_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_2_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_2_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_2_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_2_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_2_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_2_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_2_valid)	// lsu.scala:211:16
        stq_2_bits_uop_br_mask <=
          stq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1197) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1027) begin	// lsu.scala:304:5, :321:5
          if (_GEN_905) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1197) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1027) begin	// lsu.scala:304:5, :321:5
          if (_GEN_905) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_2_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_2_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_2_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_2_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_2_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_2_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_2_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_2_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_2_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_2_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_2_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_2_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_2_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_2_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_2_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_2_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_2_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_2_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_2_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_2_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1295) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_2_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_2_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_2_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1197) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1027) begin	// lsu.scala:304:5, :321:5
          if (_GEN_905) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1197) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1027) begin	// lsu.scala:304:5, :321:5
          if (_GEN_905) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_2_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_2_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_2_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_2_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_2_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_2_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_2_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_2_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_2_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_2_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_2_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_2_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_2_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_2_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_2_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_2_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_2_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_2_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_2_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_2_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_2_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_2_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_2_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_2_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_2_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_2_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_2_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_2_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_2_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1198) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1028) begin	// lsu.scala:304:5, :321:5
          if (_GEN_906) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_3_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_3_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_3_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_3_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_3_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_3_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_3_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_3_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_3_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_3_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_3_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_3_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_3_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_3_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_3_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_3_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_3_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_3_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_3_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_3_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_3_valid)	// lsu.scala:211:16
        stq_3_bits_uop_br_mask <=
          stq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1198) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1028) begin	// lsu.scala:304:5, :321:5
          if (_GEN_906) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1198) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1028) begin	// lsu.scala:304:5, :321:5
          if (_GEN_906) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_3_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_3_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_3_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_3_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_3_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_3_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_3_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_3_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_3_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_3_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_3_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_3_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_3_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_3_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_3_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_3_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_3_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_3_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_3_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_3_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1297) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_3_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_3_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_3_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1198) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1028) begin	// lsu.scala:304:5, :321:5
          if (_GEN_906) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1198) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1028) begin	// lsu.scala:304:5, :321:5
          if (_GEN_906) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_3_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_3_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_3_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_3_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_3_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_3_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_3_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_3_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_3_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_3_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_3_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_3_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_3_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_3_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_3_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_3_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_3_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_3_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_3_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_3_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_3_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_3_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_3_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_3_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_3_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_3_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_3_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_3_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_3_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1199) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1029) begin	// lsu.scala:304:5, :321:5
          if (_GEN_907) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_4_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_4_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_4_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_4_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_4_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_4_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_4_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_4_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_4_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_4_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_4_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_4_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_4_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_4_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_4_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_4_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_4_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_4_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_4_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_4_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_4_valid)	// lsu.scala:211:16
        stq_4_bits_uop_br_mask <=
          stq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1199) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1029) begin	// lsu.scala:304:5, :321:5
          if (_GEN_907) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1199) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1029) begin	// lsu.scala:304:5, :321:5
          if (_GEN_907) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_4_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_4_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_4_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_4_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_4_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_4_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_4_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_4_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_4_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_4_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_4_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_4_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_4_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_4_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_4_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_4_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_4_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_4_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_4_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_4_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1299) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_4_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_4_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_4_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1199) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1029) begin	// lsu.scala:304:5, :321:5
          if (_GEN_907) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1199) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1029) begin	// lsu.scala:304:5, :321:5
          if (_GEN_907) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_4_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_4_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_4_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_4_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_4_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_4_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_4_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_4_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_4_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_4_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_4_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_4_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_4_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_4_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_4_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_4_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_4_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_4_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_4_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_4_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_4_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_4_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_4_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_4_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_4_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_4_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_4_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_4_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_4_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1200) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1030) begin	// lsu.scala:304:5, :321:5
          if (_GEN_908) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_5_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_5_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_5_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_5_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_5_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_5_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_5_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_5_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_5_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_5_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_5_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_5_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_5_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_5_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_5_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_5_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_5_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_5_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_5_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_5_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_5_valid)	// lsu.scala:211:16
        stq_5_bits_uop_br_mask <=
          stq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1200) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1030) begin	// lsu.scala:304:5, :321:5
          if (_GEN_908) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1200) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1030) begin	// lsu.scala:304:5, :321:5
          if (_GEN_908) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_5_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_5_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_5_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_5_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_5_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_5_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_5_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_5_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_5_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_5_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_5_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_5_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_5_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_5_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_5_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_5_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_5_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_5_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_5_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_5_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1301) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_5_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_5_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_5_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1200) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1030) begin	// lsu.scala:304:5, :321:5
          if (_GEN_908) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1200) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1030) begin	// lsu.scala:304:5, :321:5
          if (_GEN_908) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_5_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_5_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_5_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_5_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_5_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_5_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_5_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_5_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_5_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_5_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_5_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_5_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_5_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_5_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_5_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_5_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_5_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_5_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_5_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_5_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_5_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_5_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_5_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_5_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_5_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_5_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_5_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_5_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_5_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1201) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1031) begin	// lsu.scala:304:5, :321:5
          if (_GEN_909) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_6_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_6_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_6_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_6_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_6_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_6_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_6_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_6_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_6_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_6_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_6_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_6_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_6_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_6_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_6_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_6_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_6_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_6_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_6_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_6_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_6_valid)	// lsu.scala:211:16
        stq_6_bits_uop_br_mask <=
          stq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1201) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1031) begin	// lsu.scala:304:5, :321:5
          if (_GEN_909) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1201) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1031) begin	// lsu.scala:304:5, :321:5
          if (_GEN_909) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_6_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_6_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_6_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_6_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_6_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_6_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_6_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_6_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_6_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_6_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_6_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_6_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_6_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_6_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_6_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_6_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_6_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_6_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_6_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_6_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1303) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_6_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_6_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_6_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1201) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1031) begin	// lsu.scala:304:5, :321:5
          if (_GEN_909) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1201) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1031) begin	// lsu.scala:304:5, :321:5
          if (_GEN_909) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_6_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_6_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_6_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_6_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_6_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_6_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_6_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_6_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_6_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_6_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_6_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_6_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_6_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_6_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_6_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_6_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_6_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_6_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_6_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_6_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_6_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_6_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_6_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_6_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_6_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_6_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_6_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_6_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_6_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1202) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1032) begin	// lsu.scala:304:5, :321:5
          if (_GEN_910) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_7_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_7_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_7_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_7_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_7_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_7_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_7_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_7_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_7_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_7_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_7_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_7_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_7_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_7_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_7_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_7_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_7_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_7_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_7_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_7_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_7_valid)	// lsu.scala:211:16
        stq_7_bits_uop_br_mask <=
          stq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1202) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1032) begin	// lsu.scala:304:5, :321:5
          if (_GEN_910) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1202) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1032) begin	// lsu.scala:304:5, :321:5
          if (_GEN_910) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_7_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_7_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_7_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_7_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_7_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_7_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_7_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_7_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_7_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_7_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_7_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_7_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_7_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_7_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_7_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_7_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_7_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_7_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_7_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_7_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1305) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_7_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_7_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_7_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1202) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1032) begin	// lsu.scala:304:5, :321:5
          if (_GEN_910) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1202) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1032) begin	// lsu.scala:304:5, :321:5
          if (_GEN_910) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_7_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_7_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_7_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_7_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_7_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_7_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_7_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_7_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_7_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_7_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_7_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_7_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_7_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_7_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_7_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_7_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_7_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_7_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_7_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_7_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_7_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_7_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_7_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_7_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_7_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_7_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_7_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_7_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_7_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1203) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1033) begin	// lsu.scala:304:5, :321:5
          if (_GEN_911) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_8_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_8_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_8_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_8_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_8_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_8_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_8_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_8_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_8_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_8_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_8_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_8_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_8_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_8_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_8_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_8_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_8_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_8_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_8_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_8_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_8_valid)	// lsu.scala:211:16
        stq_8_bits_uop_br_mask <=
          stq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1203) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1033) begin	// lsu.scala:304:5, :321:5
          if (_GEN_911) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1203) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1033) begin	// lsu.scala:304:5, :321:5
          if (_GEN_911) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_8_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_8_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_8_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_8_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_8_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_8_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_8_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_8_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_8_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_8_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_8_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_8_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_8_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_8_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_8_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_8_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_8_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_8_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_8_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_8_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1307) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_8_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_8_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_8_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1203) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1033) begin	// lsu.scala:304:5, :321:5
          if (_GEN_911) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1203) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1033) begin	// lsu.scala:304:5, :321:5
          if (_GEN_911) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_8_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_8_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_8_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_8_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_8_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_8_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_8_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_8_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_8_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_8_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_8_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_8_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_8_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_8_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_8_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_8_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_8_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_8_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_8_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_8_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_8_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_8_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_8_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_8_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_8_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_8_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_8_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_8_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_8_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1204) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1034) begin	// lsu.scala:304:5, :321:5
          if (_GEN_912) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_9_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_9_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_9_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_9_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_9_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_9_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_9_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_9_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_9_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_9_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_9_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_9_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_9_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_9_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_9_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_9_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_9_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_9_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_9_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_9_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_9_valid)	// lsu.scala:211:16
        stq_9_bits_uop_br_mask <=
          stq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1204) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1034) begin	// lsu.scala:304:5, :321:5
          if (_GEN_912) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1204) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1034) begin	// lsu.scala:304:5, :321:5
          if (_GEN_912) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_9_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_9_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_9_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_9_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_9_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_9_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_9_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_9_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_9_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_9_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_9_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_9_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_9_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_9_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_9_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_9_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_9_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_9_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_9_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_9_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1309) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_9_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_9_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_9_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1204) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1034) begin	// lsu.scala:304:5, :321:5
          if (_GEN_912) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1204) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1034) begin	// lsu.scala:304:5, :321:5
          if (_GEN_912) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_9_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_9_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_9_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_9_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_9_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_9_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_9_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_9_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_9_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_9_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_9_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_9_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_9_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_9_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_9_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_9_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_9_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_9_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_9_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_9_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_9_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_9_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_9_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_9_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_9_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_9_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_9_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_9_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_9_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1205) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1035) begin	// lsu.scala:304:5, :321:5
          if (_GEN_913) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_10_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_10_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_10_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_10_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_10_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_10_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_10_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_10_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_10_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_10_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_10_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_10_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_10_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_10_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_10_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_10_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_10_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_10_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_10_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_10_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_10_valid)	// lsu.scala:211:16
        stq_10_bits_uop_br_mask <=
          stq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1205) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1035) begin	// lsu.scala:304:5, :321:5
          if (_GEN_913) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1205) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1035) begin	// lsu.scala:304:5, :321:5
          if (_GEN_913) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_10_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_10_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_10_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_10_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_10_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_10_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_10_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_10_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_10_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_10_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_10_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_10_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_10_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_10_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_10_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_10_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_10_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_10_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_10_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_10_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1311) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_10_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_10_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_10_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1205) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1035) begin	// lsu.scala:304:5, :321:5
          if (_GEN_913) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1205) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1035) begin	// lsu.scala:304:5, :321:5
          if (_GEN_913) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_10_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_10_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_10_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_10_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_10_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_10_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_10_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_10_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_10_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_10_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_10_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_10_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_10_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_10_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_10_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_10_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_10_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_10_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_10_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_10_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_10_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_10_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_10_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_10_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_10_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_10_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_10_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_10_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_10_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1206) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1036) begin	// lsu.scala:304:5, :321:5
          if (_GEN_914) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_11_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_11_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_11_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_11_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_11_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_11_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_11_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_11_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_11_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_11_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_11_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_11_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_11_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_11_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_11_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_11_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_11_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_11_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_11_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_11_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_11_valid)	// lsu.scala:211:16
        stq_11_bits_uop_br_mask <=
          stq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1206) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1036) begin	// lsu.scala:304:5, :321:5
          if (_GEN_914) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1206) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1036) begin	// lsu.scala:304:5, :321:5
          if (_GEN_914) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_11_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_11_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_11_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_11_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_11_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_11_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_11_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_11_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_11_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_11_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_11_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_11_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_11_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_11_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_11_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_11_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_11_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_11_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_11_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_11_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1313) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_11_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_11_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_11_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1206) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1036) begin	// lsu.scala:304:5, :321:5
          if (_GEN_914) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1206) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1036) begin	// lsu.scala:304:5, :321:5
          if (_GEN_914) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_11_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_11_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_11_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_11_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_11_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_11_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_11_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_11_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_11_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_11_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_11_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_11_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_11_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_11_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_11_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_11_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_11_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_11_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_11_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_11_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_11_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_11_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_11_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_11_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_11_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_11_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_11_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_11_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_11_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1207) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1037) begin	// lsu.scala:304:5, :321:5
          if (_GEN_915) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_12_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_12_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_12_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_12_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_12_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_12_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_12_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_12_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_12_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_12_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_12_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_12_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_12_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_12_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_12_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_12_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_12_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_12_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_12_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_12_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_12_valid)	// lsu.scala:211:16
        stq_12_bits_uop_br_mask <=
          stq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1207) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1037) begin	// lsu.scala:304:5, :321:5
          if (_GEN_915) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1207) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1037) begin	// lsu.scala:304:5, :321:5
          if (_GEN_915) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_12_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_12_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_12_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_12_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_12_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_12_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_12_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_12_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_12_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_12_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_12_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_12_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_12_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_12_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_12_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_12_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_12_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_12_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_12_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_12_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1315) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_12_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_12_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_12_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1207) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1037) begin	// lsu.scala:304:5, :321:5
          if (_GEN_915) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1207) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1037) begin	// lsu.scala:304:5, :321:5
          if (_GEN_915) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_12_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_12_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_12_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_12_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_12_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_12_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_12_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_12_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_12_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_12_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_12_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_12_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_12_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_12_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_12_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_12_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_12_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_12_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_12_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_12_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_12_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_12_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_12_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_12_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_12_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_12_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_12_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_12_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_12_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1208) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1038) begin	// lsu.scala:304:5, :321:5
          if (_GEN_916) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_13_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_13_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_13_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_13_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_13_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_13_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_13_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_13_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_13_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_13_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_13_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_13_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_13_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_13_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_13_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_13_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_13_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_13_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_13_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_13_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_13_valid)	// lsu.scala:211:16
        stq_13_bits_uop_br_mask <=
          stq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1208) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1038) begin	// lsu.scala:304:5, :321:5
          if (_GEN_916) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1208) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1038) begin	// lsu.scala:304:5, :321:5
          if (_GEN_916) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_13_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_13_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_13_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_13_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_13_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_13_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_13_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_13_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_13_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_13_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_13_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_13_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_13_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_13_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_13_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_13_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_13_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_13_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_13_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_13_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1317) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_13_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_13_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_13_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1208) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1038) begin	// lsu.scala:304:5, :321:5
          if (_GEN_916) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1208) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1038) begin	// lsu.scala:304:5, :321:5
          if (_GEN_916) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_13_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_13_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_13_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_13_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_13_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_13_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_13_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_13_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_13_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_13_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_13_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_13_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_13_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_13_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_13_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_13_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_13_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_13_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_13_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_13_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_13_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_13_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_13_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_13_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_13_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_13_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_13_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_13_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_13_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1209) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1039) begin	// lsu.scala:304:5, :321:5
          if (_GEN_917) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_14_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_14_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_14_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_14_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_14_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_14_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_14_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_14_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_14_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_14_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_14_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_14_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_14_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_14_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_14_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_14_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_14_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_14_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_14_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_14_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_14_valid)	// lsu.scala:211:16
        stq_14_bits_uop_br_mask <=
          stq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1209) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1039) begin	// lsu.scala:304:5, :321:5
          if (_GEN_917) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1209) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1039) begin	// lsu.scala:304:5, :321:5
          if (_GEN_917) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_14_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_14_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_14_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_14_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_14_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_14_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_14_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_14_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_14_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_14_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_14_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_14_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_14_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_14_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_14_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_14_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_14_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_14_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_14_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_14_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1319) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_14_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_14_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_14_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1209) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1039) begin	// lsu.scala:304:5, :321:5
          if (_GEN_917) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1209) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1039) begin	// lsu.scala:304:5, :321:5
          if (_GEN_917) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_14_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_14_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_14_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_14_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_14_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_14_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_14_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_14_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_14_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_14_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_14_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_14_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_14_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_14_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_14_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_14_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_14_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_14_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_14_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_14_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_14_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_14_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_14_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_14_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_14_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_14_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_14_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_14_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_14_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1210) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1040) begin	// lsu.scala:304:5, :321:5
          if (_GEN_918) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_15_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_15_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_15_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_15_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_15_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_15_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_15_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_15_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_15_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_15_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_15_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_15_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_15_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_15_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_15_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_15_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_15_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_15_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_15_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_15_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_15_valid)	// lsu.scala:211:16
        stq_15_bits_uop_br_mask <=
          stq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1210) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1040) begin	// lsu.scala:304:5, :321:5
          if (_GEN_918) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1210) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1040) begin	// lsu.scala:304:5, :321:5
          if (_GEN_918) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_15_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_15_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_15_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_15_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_15_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_15_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_15_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_15_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_15_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_15_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_15_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_15_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_15_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_15_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_15_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_15_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_15_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_15_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_15_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_15_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1321) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_15_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_15_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_15_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1210) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1040) begin	// lsu.scala:304:5, :321:5
          if (_GEN_918) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1210) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1040) begin	// lsu.scala:304:5, :321:5
          if (_GEN_918) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_15_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_15_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_15_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_15_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_15_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_15_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_15_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_15_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_15_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_15_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_15_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_15_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_15_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_15_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_15_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_15_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_15_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_15_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_15_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_15_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_15_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_15_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_15_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_15_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_15_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_15_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_15_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_15_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_15_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1211) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1041) begin	// lsu.scala:304:5, :321:5
          if (_GEN_919) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_16_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_16_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_16_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_16_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_16_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_16_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_16_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_16_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_16_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_16_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_16_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_16_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_16_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_16_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_16_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_16_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_16_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_16_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_16_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_16_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_16_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_16_valid)	// lsu.scala:211:16
        stq_16_bits_uop_br_mask <=
          stq_16_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1211) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1041) begin	// lsu.scala:304:5, :321:5
          if (_GEN_919) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_16_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_16_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_16_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1211) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1041) begin	// lsu.scala:304:5, :321:5
          if (_GEN_919) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_16_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_16_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_16_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_16_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_16_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_16_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_16_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_16_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_16_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_16_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_16_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_16_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_16_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_16_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_16_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_16_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_16_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_16_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_16_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_16_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_16_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_16_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_16_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_16_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_16_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_16_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_16_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1323) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_16_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_16_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_16_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_16_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1211) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1041) begin	// lsu.scala:304:5, :321:5
          if (_GEN_919) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_16_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_16_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_16_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1211) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1041) begin	// lsu.scala:304:5, :321:5
          if (_GEN_919) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_16_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_16_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_16_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_16_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_16_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_16_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_16_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_16_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_16_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_16_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_16_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_16_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_16_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_16_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_16_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_16_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_16_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_16_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_16_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_16_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_16_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_16_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_16_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_16_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_16_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_16_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_16_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_16_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_16_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_16_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_16_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_16_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_16_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_16_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_16_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_16_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_16_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_16_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_16_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_16_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_16_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_16_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1212) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1042) begin	// lsu.scala:304:5, :321:5
          if (_GEN_920) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_17_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_17_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_17_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_17_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_17_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_17_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_17_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_17_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_17_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_17_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_17_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_17_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_17_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_17_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_17_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_17_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_17_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_17_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_17_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_17_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_17_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_17_valid)	// lsu.scala:211:16
        stq_17_bits_uop_br_mask <=
          stq_17_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1212) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1042) begin	// lsu.scala:304:5, :321:5
          if (_GEN_920) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_17_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_17_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_17_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1212) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1042) begin	// lsu.scala:304:5, :321:5
          if (_GEN_920) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_17_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_17_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_17_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_17_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_17_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_17_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_17_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_17_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_17_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_17_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_17_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_17_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_17_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_17_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_17_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_17_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_17_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_17_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_17_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_17_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_17_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_17_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_17_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_17_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_17_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_17_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_17_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1325) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_17_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_17_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_17_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_17_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1212) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1042) begin	// lsu.scala:304:5, :321:5
          if (_GEN_920) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_17_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_17_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_17_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1212) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1042) begin	// lsu.scala:304:5, :321:5
          if (_GEN_920) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_17_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_17_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_17_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_17_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_17_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_17_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_17_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_17_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_17_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_17_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_17_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_17_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_17_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_17_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_17_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_17_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_17_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_17_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_17_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_17_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_17_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_17_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_17_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_17_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_17_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_17_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_17_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_17_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_17_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_17_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_17_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_17_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_17_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_17_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_17_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_17_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_17_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_17_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_17_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_17_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_17_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_17_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1213) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1043) begin	// lsu.scala:304:5, :321:5
          if (_GEN_921) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_18_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_18_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_18_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_18_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_18_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_18_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_18_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_18_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_18_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_18_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_18_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_18_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_18_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_18_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_18_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_18_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_18_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_18_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_18_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_18_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_18_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_18_valid)	// lsu.scala:211:16
        stq_18_bits_uop_br_mask <=
          stq_18_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1213) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1043) begin	// lsu.scala:304:5, :321:5
          if (_GEN_921) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_18_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_18_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_18_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1213) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1043) begin	// lsu.scala:304:5, :321:5
          if (_GEN_921) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_18_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_18_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_18_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_18_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_18_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_18_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_18_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_18_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_18_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_18_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_18_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_18_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_18_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_18_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_18_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_18_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_18_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_18_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_18_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_18_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_18_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_18_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_18_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_18_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_18_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_18_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_18_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1327) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_18_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_18_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_18_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_18_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1213) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1043) begin	// lsu.scala:304:5, :321:5
          if (_GEN_921) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_18_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_18_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_18_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1213) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1043) begin	// lsu.scala:304:5, :321:5
          if (_GEN_921) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_18_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_18_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_18_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_18_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_18_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_18_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_18_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_18_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_18_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_18_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_18_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_18_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_18_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_18_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_18_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_18_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_18_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_18_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_18_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_18_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_18_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_18_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_18_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_18_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_18_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_18_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_18_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_18_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_18_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_18_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_18_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_18_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_18_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_18_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_18_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_18_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_18_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_18_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_18_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_18_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_18_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_18_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1214) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1044) begin	// lsu.scala:304:5, :321:5
          if (_GEN_922) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_19_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_19_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_19_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_19_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_19_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_19_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_19_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_19_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_19_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_19_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_19_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_19_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_19_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_19_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_19_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_19_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_19_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_19_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_19_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_19_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_19_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_19_valid)	// lsu.scala:211:16
        stq_19_bits_uop_br_mask <=
          stq_19_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1214) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1044) begin	// lsu.scala:304:5, :321:5
          if (_GEN_922) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_19_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_19_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_19_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1214) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1044) begin	// lsu.scala:304:5, :321:5
          if (_GEN_922) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_19_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_19_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_19_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_19_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_19_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_19_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_19_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_19_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_19_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_19_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_19_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_19_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_19_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_19_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_19_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_19_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_19_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_19_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_19_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_19_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_19_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_19_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_19_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_19_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_19_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_19_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_19_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1329) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_19_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_19_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_19_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_19_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1214) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1044) begin	// lsu.scala:304:5, :321:5
          if (_GEN_922) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_19_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_19_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_19_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1214) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1044) begin	// lsu.scala:304:5, :321:5
          if (_GEN_922) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_19_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_19_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_19_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_19_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_19_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_19_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_19_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_19_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_19_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_19_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_19_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_19_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_19_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_19_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_19_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_19_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_19_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_19_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_19_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_19_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_19_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_19_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_19_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_19_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_19_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_19_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_19_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_19_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_19_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_19_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_19_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_19_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_19_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_19_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_19_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_19_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_19_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_19_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_19_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_19_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_19_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_19_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1215) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1045) begin	// lsu.scala:304:5, :321:5
          if (_GEN_923) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_20_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_20_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_20_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_20_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_20_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_20_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_20_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_20_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_20_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_20_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_20_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_20_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_20_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_20_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_20_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_20_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_20_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_20_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_20_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_20_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_20_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_20_valid)	// lsu.scala:211:16
        stq_20_bits_uop_br_mask <=
          stq_20_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1215) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1045) begin	// lsu.scala:304:5, :321:5
          if (_GEN_923) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_20_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_20_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_20_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1215) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1045) begin	// lsu.scala:304:5, :321:5
          if (_GEN_923) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_20_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_20_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_20_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_20_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_20_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_20_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_20_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_20_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_20_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_20_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_20_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_20_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_20_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_20_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_20_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_20_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_20_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_20_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_20_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_20_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_20_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_20_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_20_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_20_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_20_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_20_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_20_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1331) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_20_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_20_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_20_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_20_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1215) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1045) begin	// lsu.scala:304:5, :321:5
          if (_GEN_923) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_20_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_20_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_20_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1215) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1045) begin	// lsu.scala:304:5, :321:5
          if (_GEN_923) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_20_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_20_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_20_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_20_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_20_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_20_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_20_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_20_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_20_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_20_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_20_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_20_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_20_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_20_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_20_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_20_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_20_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_20_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_20_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_20_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_20_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_20_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_20_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_20_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_20_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_20_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_20_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_20_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_20_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_20_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_20_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_20_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_20_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_20_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_20_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_20_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_20_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_20_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_20_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_20_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_20_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_20_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1216) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1046) begin	// lsu.scala:304:5, :321:5
          if (_GEN_924) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_21_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_21_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_21_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_21_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_21_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_21_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_21_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_21_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_21_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_21_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_21_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_21_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_21_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_21_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_21_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_21_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_21_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_21_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_21_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_21_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_21_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_21_valid)	// lsu.scala:211:16
        stq_21_bits_uop_br_mask <=
          stq_21_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1216) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1046) begin	// lsu.scala:304:5, :321:5
          if (_GEN_924) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_21_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_21_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_21_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1216) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1046) begin	// lsu.scala:304:5, :321:5
          if (_GEN_924) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_21_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_21_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_21_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_21_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_21_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_21_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_21_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_21_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_21_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_21_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_21_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_21_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_21_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_21_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_21_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_21_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_21_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_21_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_21_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_21_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_21_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_21_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_21_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_21_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_21_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_21_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_21_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1333) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_21_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_21_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_21_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_21_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1216) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1046) begin	// lsu.scala:304:5, :321:5
          if (_GEN_924) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_21_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_21_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_21_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1216) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1046) begin	// lsu.scala:304:5, :321:5
          if (_GEN_924) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_21_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_21_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_21_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_21_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_21_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_21_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_21_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_21_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_21_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_21_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_21_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_21_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_21_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_21_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_21_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_21_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_21_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_21_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_21_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_21_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_21_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_21_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_21_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_21_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_21_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_21_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_21_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_21_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_21_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_21_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_21_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_21_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_21_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_21_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_21_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_21_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_21_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_21_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_21_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_21_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_21_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_21_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1217) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1047) begin	// lsu.scala:304:5, :321:5
          if (_GEN_925) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_22_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_22_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_22_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_22_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_22_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_22_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_22_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_22_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_22_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_22_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_22_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_22_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_22_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_22_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_22_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_22_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_22_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_22_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_22_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_22_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_22_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_22_valid)	// lsu.scala:211:16
        stq_22_bits_uop_br_mask <=
          stq_22_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1217) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1047) begin	// lsu.scala:304:5, :321:5
          if (_GEN_925) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_22_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_22_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_22_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1217) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1047) begin	// lsu.scala:304:5, :321:5
          if (_GEN_925) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_22_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_22_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_22_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_22_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_22_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_22_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_22_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_22_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_22_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_22_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_22_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_22_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_22_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_22_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_22_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_22_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_22_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_22_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_22_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_22_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_22_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_22_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_22_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_22_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_22_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_22_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_22_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1335) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_22_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_22_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_22_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_22_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1217) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1047) begin	// lsu.scala:304:5, :321:5
          if (_GEN_925) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_22_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_22_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_22_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1217) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1047) begin	// lsu.scala:304:5, :321:5
          if (_GEN_925) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_22_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_22_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_22_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_22_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_22_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_22_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_22_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_22_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_22_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_22_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_22_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_22_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_22_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_22_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_22_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_22_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_22_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_22_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_22_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_22_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_22_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_22_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_22_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_22_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_22_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_22_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_22_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_22_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_22_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_22_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_22_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_22_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_22_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_22_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_22_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_22_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_22_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_22_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_22_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_22_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_22_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_22_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_1218) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1048) begin	// lsu.scala:304:5, :321:5
          if (_GEN_926) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_23_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
            stq_23_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
            stq_23_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
            stq_23_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
            stq_23_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
            stq_23_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
            stq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
            stq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
            stq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
            stq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
            stq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
            stq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
            stq_23_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_23_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
          stq_23_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
          stq_23_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
          stq_23_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
          stq_23_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
          stq_23_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
          stq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_23_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_23_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;	// lsu.scala:211:16
        stq_23_bits_uop_inst <= io_core_dis_uops_2_bits_inst;	// lsu.scala:211:16
        stq_23_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;	// lsu.scala:211:16
        stq_23_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;	// lsu.scala:211:16
        stq_23_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;	// lsu.scala:211:16
        stq_23_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_23_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_23_valid)	// lsu.scala:211:16
        stq_23_bits_uop_br_mask <=
          stq_23_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_1218) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1048) begin	// lsu.scala:304:5, :321:5
          if (_GEN_926) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_23_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_23_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_23_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_1218) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1048) begin	// lsu.scala:304:5, :321:5
          if (_GEN_926) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_23_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
            stq_23_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
            stq_23_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
            stq_23_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
            stq_23_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
            stq_23_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
            stq_23_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
            stq_23_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
            stq_23_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_23_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
          stq_23_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
          stq_23_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
          stq_23_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
          stq_23_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
          stq_23_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
          stq_23_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
          stq_23_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
          stq_23_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_23_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;	// lsu.scala:211:16
        stq_23_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;	// lsu.scala:211:16
        stq_23_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;	// lsu.scala:211:16
        stq_23_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;	// lsu.scala:211:16
        stq_23_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;	// lsu.scala:211:16
        stq_23_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;	// lsu.scala:211:16
        stq_23_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;	// lsu.scala:211:16
        stq_23_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;	// lsu.scala:211:16
        stq_23_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_1337) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_23_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_23_bits_uop_pdst <= _GEN_154;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_23_bits_uop_pdst <= _GEN_207;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_23_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_1218) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1048) begin	// lsu.scala:304:5, :321:5
          if (_GEN_926) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else	// lsu.scala:211:16, :304:5, :321:5
            stq_23_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
        end
        else	// lsu.scala:304:5, :321:5
          stq_23_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_23_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;	// lsu.scala:211:16
      if (_GEN_1218) begin	// lsu.scala:304:5, :321:5
        if (_GEN_1048) begin	// lsu.scala:304:5, :321:5
          if (_GEN_926) begin	// lsu.scala:211:16, :304:5, :321:5
          end
          else begin	// lsu.scala:211:16, :304:5, :321:5
            stq_23_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
            stq_23_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
            stq_23_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
            stq_23_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
            stq_23_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
            stq_23_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
            stq_23_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
            stq_23_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
            stq_23_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
            stq_23_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
            stq_23_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
            stq_23_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
            stq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
            stq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
            stq_23_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
            stq_23_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
          end
        end
        else begin	// lsu.scala:304:5, :321:5
          stq_23_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
          stq_23_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
          stq_23_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
          stq_23_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
          stq_23_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
          stq_23_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
          stq_23_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
          stq_23_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
          stq_23_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
          stq_23_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
          stq_23_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
          stq_23_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
          stq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_23_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
          stq_23_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_23_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;	// lsu.scala:211:16
        stq_23_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;	// lsu.scala:211:16
        stq_23_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;	// lsu.scala:211:16
        stq_23_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;	// lsu.scala:211:16
        stq_23_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;	// lsu.scala:211:16
        stq_23_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;	// lsu.scala:211:16
        stq_23_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;	// lsu.scala:211:16
        stq_23_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;	// lsu.scala:211:16
        stq_23_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;	// lsu.scala:211:16
        stq_23_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;	// lsu.scala:211:16
        stq_23_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;	// lsu.scala:211:16
        stq_23_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;	// lsu.scala:211:16
        stq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_23_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;	// lsu.scala:211:16
        stq_23_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (clear_store) begin	// lsu.scala:1495:3, :1500:17
        if (stq_head == 5'h17)	// lsu.scala:217:29, util.scala:205:25
          stq_head <= 5'h0;	// lsu.scala:217:29
        else	// util.scala:205:25
          stq_head <= stq_head + 5'h1;	// lsu.scala:217:29, :305:44, util.scala:206:28
      end
      if (commit_store_2) begin	// lsu.scala:1451:49
        if (_GEN_831 == 5'h17)	// lsu.scala:1482:31, util.scala:205:25
          stq_commit_head <= 5'h0;	// lsu.scala:219:29
        else	// util.scala:205:25
          stq_commit_head <= _GEN_831 + 5'h1;	// lsu.scala:219:29, :305:44, :1482:31, util.scala:206:28
      end
      else if (commit_store_1) begin	// lsu.scala:1451:49
        if (wrap_14)	// util.scala:205:25
          stq_commit_head <= 5'h0;	// lsu.scala:219:29
        else	// util.scala:205:25
          stq_commit_head <= _GEN_830;	// lsu.scala:219:29, util.scala:206:28
      end
      else if (commit_store) begin	// lsu.scala:1451:49
        if (wrap_12)	// util.scala:205:25
          stq_commit_head <= 5'h0;	// lsu.scala:219:29
        else	// util.scala:205:25
          stq_commit_head <= _GEN_826;	// lsu.scala:219:29, util.scala:206:28
      end
      if (clear_store & _GEN_845) begin	// lsu.scala:1284:5, :1494:29, :1495:3, :1500:17, :1505:3, :1514:5, :1515:24
        if (stq_execute_head == 5'h17)	// lsu.scala:220:29, util.scala:205:25
          stq_execute_head <= 5'h0;	// lsu.scala:220:29
        else	// util.scala:205:25
          stq_execute_head <= stq_execute_head + 5'h1;	// lsu.scala:220:29, :305:44, util.scala:206:28
      end
      else if (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
               | io_dmem_nack_0_bits_uop_uses_ldq
               | io_dmem_nack_0_bits_uop_stq_idx < stq_head ^ stq_execute_head < stq_head
               ^ io_dmem_nack_0_bits_uop_stq_idx >= stq_execute_head) begin	// lsu.scala:217:29, :220:29, :766:39, :1174:30, :1284:5, :1287:7, :1291:7, :1299:86, util.scala:363:{52,64,78}
        if (_GEN_315 | ~(will_fire_store_commit_0 & dmem_req_fire_0)) begin	// lsu.scala:220:29, :535:65, :752:55, :766:39, :773:43, :780:45, :789:{44,50}
        end
        else if (stq_execute_head == 5'h17)	// lsu.scala:220:29, util.scala:205:25
          stq_execute_head <= 5'h0;	// lsu.scala:220:29
        else	// util.scala:205:25
          stq_execute_head <= stq_execute_head + 5'h1;	// lsu.scala:220:29, :305:44, util.scala:206:28
      end
      else	// lsu.scala:766:39, :1284:5, :1287:7
        stq_execute_head <= io_dmem_nack_0_bits_uop_stq_idx;	// lsu.scala:220:29
    end
    stq_0_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1195)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_903) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1001 | ~_GEN_903)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_0_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1195 & _GEN_1025 & _GEN_903 & stq_0_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h0
         | (_GEN_1195
              ? (_GEN_1025
                   ? (_GEN_903
                        ? stq_0_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903 ? stq_0_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1195
           ? (_GEN_1025
                ? (_GEN_903
                     ? stq_0_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_addr_valid <=
      ~_GEN_2427 & (clear_store ? ~_GEN_2350 & _GEN_1292 : ~_GEN_2108 & _GEN_1292);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1291) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_0_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_0_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_0_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_0_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_0_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_0_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_0_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_0_bits_data_valid <=
      ~_GEN_2427 & (clear_store ? ~_GEN_2350 & _GEN_1340 : ~_GEN_2108 & _GEN_1340);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1339) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_0_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_0_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_0_bits_committed <=
      ~_GEN_2397
      & (commit_store_2 & _GEN_2301
         | (commit_store_1 ? _GEN_2253 | _GEN_2157 | _GEN_1219 : _GEN_2157 | _GEN_1219));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_0_bits_succeeded <=
      ~_GEN_2397
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h0
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h0)) & _GEN_1195
         & _GEN_1025 & _GEN_903 & stq_0_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_1_valid <=
      ~_GEN_2429 & (clear_store ? ~_GEN_2352 & _GEN_1150 : ~_GEN_2109 & _GEN_1150);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_1_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1196)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_904) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1002 | ~_GEN_904)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_1_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1196 & _GEN_1026 & _GEN_904 & stq_1_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1
         | (_GEN_1196
              ? (_GEN_1026
                   ? (_GEN_904
                        ? stq_1_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904 ? stq_1_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1196
           ? (_GEN_1026
                ? (_GEN_904
                     ? stq_1_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_addr_valid <=
      ~_GEN_2429 & (clear_store ? ~_GEN_2352 & _GEN_1294 : ~_GEN_2109 & _GEN_1294);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1293) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_1_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_1_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_1_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_1_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_1_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_1_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_1_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_1_bits_data_valid <=
      ~_GEN_2429 & (clear_store ? ~_GEN_2352 & _GEN_1342 : ~_GEN_2109 & _GEN_1342);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1341) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_1_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_1_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_1_bits_committed <=
      ~_GEN_2398
      & (commit_store_2 & _GEN_2302
         | (commit_store_1 ? _GEN_2254 | _GEN_2159 | _GEN_1220 : _GEN_2159 | _GEN_1220));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_1_bits_succeeded <=
      ~_GEN_2398
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h1)) & _GEN_1196
         & _GEN_1026 & _GEN_904 & stq_1_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_2_valid <=
      ~_GEN_2431 & (clear_store ? ~_GEN_2354 & _GEN_1152 : ~_GEN_2110 & _GEN_1152);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_2_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1197)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_905) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1003 | ~_GEN_905)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_2_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1197 & _GEN_1027 & _GEN_905 & stq_2_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h2
         | (_GEN_1197
              ? (_GEN_1027
                   ? (_GEN_905
                        ? stq_2_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905 ? stq_2_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1197
           ? (_GEN_1027
                ? (_GEN_905
                     ? stq_2_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_addr_valid <=
      ~_GEN_2431 & (clear_store ? ~_GEN_2354 & _GEN_1296 : ~_GEN_2110 & _GEN_1296);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1295) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_2_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_2_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_2_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_2_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_2_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_2_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_2_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_2_bits_data_valid <=
      ~_GEN_2431 & (clear_store ? ~_GEN_2354 & _GEN_1344 : ~_GEN_2110 & _GEN_1344);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1343) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_2_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_2_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_2_bits_committed <=
      ~_GEN_2399
      & (commit_store_2 & _GEN_2303
         | (commit_store_1 ? _GEN_2255 | _GEN_2161 | _GEN_1221 : _GEN_2161 | _GEN_1221));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_2_bits_succeeded <=
      ~_GEN_2399
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h2
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h2)) & _GEN_1197
         & _GEN_1027 & _GEN_905 & stq_2_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_3_valid <=
      ~_GEN_2433 & (clear_store ? ~_GEN_2356 & _GEN_1154 : ~_GEN_2111 & _GEN_1154);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_3_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1198)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_906) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1004 | ~_GEN_906)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_3_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1198 & _GEN_1028 & _GEN_906 & stq_3_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h3
         | (_GEN_1198
              ? (_GEN_1028
                   ? (_GEN_906
                        ? stq_3_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906 ? stq_3_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1198
           ? (_GEN_1028
                ? (_GEN_906
                     ? stq_3_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_addr_valid <=
      ~_GEN_2433 & (clear_store ? ~_GEN_2356 & _GEN_1298 : ~_GEN_2111 & _GEN_1298);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1297) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_3_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_3_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_3_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_3_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_3_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_3_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_3_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_3_bits_data_valid <=
      ~_GEN_2433 & (clear_store ? ~_GEN_2356 & _GEN_1346 : ~_GEN_2111 & _GEN_1346);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1345) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_3_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_3_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_3_bits_committed <=
      ~_GEN_2400
      & (commit_store_2 & _GEN_2304
         | (commit_store_1 ? _GEN_2256 | _GEN_2163 | _GEN_1222 : _GEN_2163 | _GEN_1222));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_3_bits_succeeded <=
      ~_GEN_2400
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h3
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h3)) & _GEN_1198
         & _GEN_1028 & _GEN_906 & stq_3_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_4_valid <=
      ~_GEN_2435 & (clear_store ? ~_GEN_2358 & _GEN_1156 : ~_GEN_2112 & _GEN_1156);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_4_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1199)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_907) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1005 | ~_GEN_907)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_4_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1199 & _GEN_1029 & _GEN_907 & stq_4_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h4
         | (_GEN_1199
              ? (_GEN_1029
                   ? (_GEN_907
                        ? stq_4_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907 ? stq_4_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1199
           ? (_GEN_1029
                ? (_GEN_907
                     ? stq_4_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_addr_valid <=
      ~_GEN_2435 & (clear_store ? ~_GEN_2358 & _GEN_1300 : ~_GEN_2112 & _GEN_1300);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1299) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_4_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_4_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_4_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_4_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_4_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_4_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_4_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_4_bits_data_valid <=
      ~_GEN_2435 & (clear_store ? ~_GEN_2358 & _GEN_1348 : ~_GEN_2112 & _GEN_1348);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1347) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_4_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_4_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_4_bits_committed <=
      ~_GEN_2401
      & (commit_store_2 & _GEN_2305
         | (commit_store_1 ? _GEN_2257 | _GEN_2165 | _GEN_1223 : _GEN_2165 | _GEN_1223));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_4_bits_succeeded <=
      ~_GEN_2401
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h4
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h4)) & _GEN_1199
         & _GEN_1029 & _GEN_907 & stq_4_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_5_valid <=
      ~_GEN_2437 & (clear_store ? ~_GEN_2360 & _GEN_1158 : ~_GEN_2113 & _GEN_1158);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_5_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1200)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_908) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1006 | ~_GEN_908)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_5_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1200 & _GEN_1030 & _GEN_908 & stq_5_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h5
         | (_GEN_1200
              ? (_GEN_1030
                   ? (_GEN_908
                        ? stq_5_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908 ? stq_5_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1200
           ? (_GEN_1030
                ? (_GEN_908
                     ? stq_5_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_addr_valid <=
      ~_GEN_2437 & (clear_store ? ~_GEN_2360 & _GEN_1302 : ~_GEN_2113 & _GEN_1302);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1301) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_5_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_5_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_5_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_5_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_5_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_5_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_5_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_5_bits_data_valid <=
      ~_GEN_2437 & (clear_store ? ~_GEN_2360 & _GEN_1350 : ~_GEN_2113 & _GEN_1350);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1349) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_5_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_5_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_5_bits_committed <=
      ~_GEN_2402
      & (commit_store_2 & _GEN_2306
         | (commit_store_1 ? _GEN_2258 | _GEN_2167 | _GEN_1224 : _GEN_2167 | _GEN_1224));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_5_bits_succeeded <=
      ~_GEN_2402
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h5
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h5)) & _GEN_1200
         & _GEN_1030 & _GEN_908 & stq_5_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_6_valid <=
      ~_GEN_2439 & (clear_store ? ~_GEN_2362 & _GEN_1160 : ~_GEN_2114 & _GEN_1160);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_6_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1201)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_909) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1007 | ~_GEN_909)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_6_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1201 & _GEN_1031 & _GEN_909 & stq_6_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h6
         | (_GEN_1201
              ? (_GEN_1031
                   ? (_GEN_909
                        ? stq_6_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909 ? stq_6_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1201
           ? (_GEN_1031
                ? (_GEN_909
                     ? stq_6_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_addr_valid <=
      ~_GEN_2439 & (clear_store ? ~_GEN_2362 & _GEN_1304 : ~_GEN_2114 & _GEN_1304);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1303) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_6_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_6_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_6_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_6_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_6_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_6_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_6_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_6_bits_data_valid <=
      ~_GEN_2439 & (clear_store ? ~_GEN_2362 & _GEN_1352 : ~_GEN_2114 & _GEN_1352);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1351) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_6_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_6_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_6_bits_committed <=
      ~_GEN_2403
      & (commit_store_2 & _GEN_2307
         | (commit_store_1 ? _GEN_2259 | _GEN_2169 | _GEN_1225 : _GEN_2169 | _GEN_1225));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_6_bits_succeeded <=
      ~_GEN_2403
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h6
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h6)) & _GEN_1201
         & _GEN_1031 & _GEN_909 & stq_6_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_7_valid <=
      ~_GEN_2441 & (clear_store ? ~_GEN_2364 & _GEN_1162 : ~_GEN_2115 & _GEN_1162);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_7_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1202)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_910) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1008 | ~_GEN_910)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_7_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1202 & _GEN_1032 & _GEN_910 & stq_7_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h7
         | (_GEN_1202
              ? (_GEN_1032
                   ? (_GEN_910
                        ? stq_7_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910 ? stq_7_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1202
           ? (_GEN_1032
                ? (_GEN_910
                     ? stq_7_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_addr_valid <=
      ~_GEN_2441 & (clear_store ? ~_GEN_2364 & _GEN_1306 : ~_GEN_2115 & _GEN_1306);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1305) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_7_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_7_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_7_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_7_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_7_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_7_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_7_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_7_bits_data_valid <=
      ~_GEN_2441 & (clear_store ? ~_GEN_2364 & _GEN_1354 : ~_GEN_2115 & _GEN_1354);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1353) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_7_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_7_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_7_bits_committed <=
      ~_GEN_2404
      & (commit_store_2 & _GEN_2308
         | (commit_store_1 ? _GEN_2260 | _GEN_2171 | _GEN_1226 : _GEN_2171 | _GEN_1226));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_7_bits_succeeded <=
      ~_GEN_2404
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h7
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h7)) & _GEN_1202
         & _GEN_1032 & _GEN_910 & stq_7_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_8_valid <=
      ~_GEN_2443 & (clear_store ? ~_GEN_2366 & _GEN_1164 : ~_GEN_2116 & _GEN_1164);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_8_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1203)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_911) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1009 | ~_GEN_911)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_8_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1203 & _GEN_1033 & _GEN_911 & stq_8_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h8
         | (_GEN_1203
              ? (_GEN_1033
                   ? (_GEN_911
                        ? stq_8_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911 ? stq_8_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1203
           ? (_GEN_1033
                ? (_GEN_911
                     ? stq_8_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_addr_valid <=
      ~_GEN_2443 & (clear_store ? ~_GEN_2366 & _GEN_1308 : ~_GEN_2116 & _GEN_1308);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1307) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_8_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_8_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_8_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_8_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_8_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_8_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_8_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_8_bits_data_valid <=
      ~_GEN_2443 & (clear_store ? ~_GEN_2366 & _GEN_1356 : ~_GEN_2116 & _GEN_1356);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1355) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_8_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_8_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_8_bits_committed <=
      ~_GEN_2405
      & (commit_store_2 & _GEN_2309
         | (commit_store_1 ? _GEN_2261 | _GEN_2173 | _GEN_1227 : _GEN_2173 | _GEN_1227));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_8_bits_succeeded <=
      ~_GEN_2405
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h8
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h8)) & _GEN_1203
         & _GEN_1033 & _GEN_911 & stq_8_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_9_valid <=
      ~_GEN_2445 & (clear_store ? ~_GEN_2368 & _GEN_1166 : ~_GEN_2117 & _GEN_1166);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_9_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1204)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_912) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1010 | ~_GEN_912)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_9_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1204 & _GEN_1034 & _GEN_912 & stq_9_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h9
         | (_GEN_1204
              ? (_GEN_1034
                   ? (_GEN_912
                        ? stq_9_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912 ? stq_9_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1204
           ? (_GEN_1034
                ? (_GEN_912
                     ? stq_9_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_addr_valid <=
      ~_GEN_2445 & (clear_store ? ~_GEN_2368 & _GEN_1310 : ~_GEN_2117 & _GEN_1310);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1309) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_9_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_9_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_9_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_9_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_9_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_9_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_9_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_9_bits_data_valid <=
      ~_GEN_2445 & (clear_store ? ~_GEN_2368 & _GEN_1358 : ~_GEN_2117 & _GEN_1358);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1357) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_9_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_9_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_9_bits_committed <=
      ~_GEN_2406
      & (commit_store_2 & _GEN_2310
         | (commit_store_1 ? _GEN_2262 | _GEN_2175 | _GEN_1228 : _GEN_2175 | _GEN_1228));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_9_bits_succeeded <=
      ~_GEN_2406
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h9
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h9)) & _GEN_1204
         & _GEN_1034 & _GEN_912 & stq_9_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_10_valid <=
      ~_GEN_2447 & (clear_store ? ~_GEN_2370 & _GEN_1168 : ~_GEN_2118 & _GEN_1168);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_10_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1205)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_913) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1011 | ~_GEN_913)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_10_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1205 & _GEN_1035 & _GEN_913 & stq_10_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hA
         | (_GEN_1205
              ? (_GEN_1035
                   ? (_GEN_913
                        ? stq_10_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913 ? stq_10_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1205
           ? (_GEN_1035
                ? (_GEN_913
                     ? stq_10_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_addr_valid <=
      ~_GEN_2447 & (clear_store ? ~_GEN_2370 & _GEN_1312 : ~_GEN_2118 & _GEN_1312);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1311) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_10_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_10_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_10_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_10_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_10_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_10_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_10_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_10_bits_data_valid <=
      ~_GEN_2447 & (clear_store ? ~_GEN_2370 & _GEN_1360 : ~_GEN_2118 & _GEN_1360);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1359) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_10_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_10_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_10_bits_committed <=
      ~_GEN_2407
      & (commit_store_2 & _GEN_2311
         | (commit_store_1 ? _GEN_2263 | _GEN_2177 | _GEN_1229 : _GEN_2177 | _GEN_1229));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_10_bits_succeeded <=
      ~_GEN_2407
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hA
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hA)) & _GEN_1205
         & _GEN_1035 & _GEN_913 & stq_10_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_11_valid <=
      ~_GEN_2449 & (clear_store ? ~_GEN_2372 & _GEN_1170 : ~_GEN_2119 & _GEN_1170);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_11_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1206)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_914) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1012 | ~_GEN_914)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_11_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1206 & _GEN_1036 & _GEN_914 & stq_11_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hB
         | (_GEN_1206
              ? (_GEN_1036
                   ? (_GEN_914
                        ? stq_11_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914 ? stq_11_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1206
           ? (_GEN_1036
                ? (_GEN_914
                     ? stq_11_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_addr_valid <=
      ~_GEN_2449 & (clear_store ? ~_GEN_2372 & _GEN_1314 : ~_GEN_2119 & _GEN_1314);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1313) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_11_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_11_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_11_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_11_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_11_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_11_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_11_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_11_bits_data_valid <=
      ~_GEN_2449 & (clear_store ? ~_GEN_2372 & _GEN_1362 : ~_GEN_2119 & _GEN_1362);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1361) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_11_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_11_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_11_bits_committed <=
      ~_GEN_2408
      & (commit_store_2 & _GEN_2312
         | (commit_store_1 ? _GEN_2264 | _GEN_2179 | _GEN_1230 : _GEN_2179 | _GEN_1230));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_11_bits_succeeded <=
      ~_GEN_2408
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hB
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hB)) & _GEN_1206
         & _GEN_1036 & _GEN_914 & stq_11_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_12_valid <=
      ~_GEN_2451 & (clear_store ? ~_GEN_2374 & _GEN_1172 : ~_GEN_2120 & _GEN_1172);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_12_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1207)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_915) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1013 | ~_GEN_915)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_12_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1207 & _GEN_1037 & _GEN_915 & stq_12_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hC
         | (_GEN_1207
              ? (_GEN_1037
                   ? (_GEN_915
                        ? stq_12_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915 ? stq_12_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1207
           ? (_GEN_1037
                ? (_GEN_915
                     ? stq_12_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_addr_valid <=
      ~_GEN_2451 & (clear_store ? ~_GEN_2374 & _GEN_1316 : ~_GEN_2120 & _GEN_1316);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1315) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_12_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_12_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_12_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_12_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_12_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_12_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_12_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_12_bits_data_valid <=
      ~_GEN_2451 & (clear_store ? ~_GEN_2374 & _GEN_1364 : ~_GEN_2120 & _GEN_1364);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1363) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_12_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_12_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_12_bits_committed <=
      ~_GEN_2409
      & (commit_store_2 & _GEN_2313
         | (commit_store_1 ? _GEN_2265 | _GEN_2181 | _GEN_1231 : _GEN_2181 | _GEN_1231));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_12_bits_succeeded <=
      ~_GEN_2409
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hC
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hC)) & _GEN_1207
         & _GEN_1037 & _GEN_915 & stq_12_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_13_valid <=
      ~_GEN_2453 & (clear_store ? ~_GEN_2376 & _GEN_1174 : ~_GEN_2121 & _GEN_1174);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_13_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1208)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_916) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1014 | ~_GEN_916)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_13_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1208 & _GEN_1038 & _GEN_916 & stq_13_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hD
         | (_GEN_1208
              ? (_GEN_1038
                   ? (_GEN_916
                        ? stq_13_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916 ? stq_13_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1208
           ? (_GEN_1038
                ? (_GEN_916
                     ? stq_13_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_addr_valid <=
      ~_GEN_2453 & (clear_store ? ~_GEN_2376 & _GEN_1318 : ~_GEN_2121 & _GEN_1318);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1317) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_13_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_13_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_13_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_13_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_13_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_13_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_13_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_13_bits_data_valid <=
      ~_GEN_2453 & (clear_store ? ~_GEN_2376 & _GEN_1366 : ~_GEN_2121 & _GEN_1366);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1365) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_13_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_13_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_13_bits_committed <=
      ~_GEN_2410
      & (commit_store_2 & _GEN_2314
         | (commit_store_1 ? _GEN_2266 | _GEN_2183 | _GEN_1232 : _GEN_2183 | _GEN_1232));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_13_bits_succeeded <=
      ~_GEN_2410
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hD
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hD)) & _GEN_1208
         & _GEN_1038 & _GEN_916 & stq_13_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_14_valid <=
      ~_GEN_2455 & (clear_store ? ~_GEN_2378 & _GEN_1176 : ~_GEN_2122 & _GEN_1176);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_14_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1209)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_917) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1015 | ~_GEN_917)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_14_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1209 & _GEN_1039 & _GEN_917 & stq_14_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hE
         | (_GEN_1209
              ? (_GEN_1039
                   ? (_GEN_917
                        ? stq_14_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917 ? stq_14_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1209
           ? (_GEN_1039
                ? (_GEN_917
                     ? stq_14_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_addr_valid <=
      ~_GEN_2455 & (clear_store ? ~_GEN_2378 & _GEN_1320 : ~_GEN_2122 & _GEN_1320);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1319) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_14_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_14_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_14_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_14_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_14_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_14_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_14_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_14_bits_data_valid <=
      ~_GEN_2455 & (clear_store ? ~_GEN_2378 & _GEN_1368 : ~_GEN_2122 & _GEN_1368);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1367) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_14_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_14_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_14_bits_committed <=
      ~_GEN_2411
      & (commit_store_2 & _GEN_2315
         | (commit_store_1 ? _GEN_2267 | _GEN_2185 | _GEN_1233 : _GEN_2185 | _GEN_1233));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_14_bits_succeeded <=
      ~_GEN_2411
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hE
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hE)) & _GEN_1209
         & _GEN_1039 & _GEN_917 & stq_14_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_15_valid <=
      ~_GEN_2457 & (clear_store ? ~_GEN_2380 & _GEN_1178 : ~_GEN_2123 & _GEN_1178);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_15_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1210)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_918) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1016 | ~_GEN_918)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_15_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1210 & _GEN_1040 & _GEN_918 & stq_15_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hF
         | (_GEN_1210
              ? (_GEN_1040
                   ? (_GEN_918
                        ? stq_15_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918 ? stq_15_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1210
           ? (_GEN_1040
                ? (_GEN_918
                     ? stq_15_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_addr_valid <=
      ~_GEN_2457 & (clear_store ? ~_GEN_2380 & _GEN_1322 : ~_GEN_2123 & _GEN_1322);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1321) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_15_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_15_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_15_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_15_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_15_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_15_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_15_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_15_bits_data_valid <=
      ~_GEN_2457 & (clear_store ? ~_GEN_2380 & _GEN_1370 : ~_GEN_2123 & _GEN_1370);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1369) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_15_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_15_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_15_bits_committed <=
      ~_GEN_2412
      & (commit_store_2 & _GEN_2316
         | (commit_store_1 ? _GEN_2268 | _GEN_2187 | _GEN_1234 : _GEN_2187 | _GEN_1234));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_15_bits_succeeded <=
      ~_GEN_2412
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hF
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hF)) & _GEN_1210
         & _GEN_1040 & _GEN_918 & stq_15_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_16_valid <=
      ~_GEN_2459 & (clear_store ? ~_GEN_2382 & _GEN_1180 : ~_GEN_2124 & _GEN_1180);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_16_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1211)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_16_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_919) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_16_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1017 | ~_GEN_919)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_16_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_16_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1211 & _GEN_1041 & _GEN_919 & stq_16_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h10
         | (_GEN_1211
              ? (_GEN_1041
                   ? (_GEN_919
                        ? stq_16_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919 ? stq_16_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1211
           ? (_GEN_1041
                ? (_GEN_919
                     ? stq_16_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_16_bits_addr_valid <=
      ~_GEN_2459 & (clear_store ? ~_GEN_2382 & _GEN_1324 : ~_GEN_2124 & _GEN_1324);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1323) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_16_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_16_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_16_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_16_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_16_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_16_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_16_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_16_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_16_bits_data_valid <=
      ~_GEN_2459 & (clear_store ? ~_GEN_2382 & _GEN_1372 : ~_GEN_2124 & _GEN_1372);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1371) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_16_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_16_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_16_bits_committed <=
      ~_GEN_2413
      & (commit_store_2 & _GEN_2317
         | (commit_store_1 ? _GEN_2269 | _GEN_2189 | _GEN_1235 : _GEN_2189 | _GEN_1235));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_16_bits_succeeded <=
      ~_GEN_2413
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h10
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h10))
         & _GEN_1211 & _GEN_1041 & _GEN_919 & stq_16_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_17_valid <=
      ~_GEN_2461 & (clear_store ? ~_GEN_2384 & _GEN_1182 : ~_GEN_2125 & _GEN_1182);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_17_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1212)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_17_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_920) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_17_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1018 | ~_GEN_920)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_17_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_17_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1212 & _GEN_1042 & _GEN_920 & stq_17_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h11
         | (_GEN_1212
              ? (_GEN_1042
                   ? (_GEN_920
                        ? stq_17_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920 ? stq_17_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1212
           ? (_GEN_1042
                ? (_GEN_920
                     ? stq_17_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_17_bits_addr_valid <=
      ~_GEN_2461 & (clear_store ? ~_GEN_2384 & _GEN_1326 : ~_GEN_2125 & _GEN_1326);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1325) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_17_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_17_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_17_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_17_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_17_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_17_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_17_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_17_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_17_bits_data_valid <=
      ~_GEN_2461 & (clear_store ? ~_GEN_2384 & _GEN_1374 : ~_GEN_2125 & _GEN_1374);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1373) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_17_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_17_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_17_bits_committed <=
      ~_GEN_2414
      & (commit_store_2 & _GEN_2318
         | (commit_store_1 ? _GEN_2270 | _GEN_2191 | _GEN_1236 : _GEN_2191 | _GEN_1236));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_17_bits_succeeded <=
      ~_GEN_2414
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h11
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h11))
         & _GEN_1212 & _GEN_1042 & _GEN_920 & stq_17_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_18_valid <=
      ~_GEN_2463 & (clear_store ? ~_GEN_2386 & _GEN_1184 : ~_GEN_2126 & _GEN_1184);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_18_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1213)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_18_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_921) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_18_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1019 | ~_GEN_921)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_18_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_18_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1213 & _GEN_1043 & _GEN_921 & stq_18_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h12
         | (_GEN_1213
              ? (_GEN_1043
                   ? (_GEN_921
                        ? stq_18_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921 ? stq_18_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1213
           ? (_GEN_1043
                ? (_GEN_921
                     ? stq_18_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_18_bits_addr_valid <=
      ~_GEN_2463 & (clear_store ? ~_GEN_2386 & _GEN_1328 : ~_GEN_2126 & _GEN_1328);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1327) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_18_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_18_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_18_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_18_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_18_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_18_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_18_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_18_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_18_bits_data_valid <=
      ~_GEN_2463 & (clear_store ? ~_GEN_2386 & _GEN_1376 : ~_GEN_2126 & _GEN_1376);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1375) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_18_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_18_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_18_bits_committed <=
      ~_GEN_2415
      & (commit_store_2 & _GEN_2319
         | (commit_store_1 ? _GEN_2271 | _GEN_2193 | _GEN_1237 : _GEN_2193 | _GEN_1237));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_18_bits_succeeded <=
      ~_GEN_2415
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h12
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h12))
         & _GEN_1213 & _GEN_1043 & _GEN_921 & stq_18_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_19_valid <=
      ~_GEN_2465 & (clear_store ? ~_GEN_2388 & _GEN_1186 : ~_GEN_2127 & _GEN_1186);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_19_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1214)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_19_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_922) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_19_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1020 | ~_GEN_922)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_19_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_19_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1214 & _GEN_1044 & _GEN_922 & stq_19_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h13
         | (_GEN_1214
              ? (_GEN_1044
                   ? (_GEN_922
                        ? stq_19_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922 ? stq_19_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1214
           ? (_GEN_1044
                ? (_GEN_922
                     ? stq_19_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_19_bits_addr_valid <=
      ~_GEN_2465 & (clear_store ? ~_GEN_2388 & _GEN_1330 : ~_GEN_2127 & _GEN_1330);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1329) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_19_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_19_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_19_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_19_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_19_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_19_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_19_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_19_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_19_bits_data_valid <=
      ~_GEN_2465 & (clear_store ? ~_GEN_2388 & _GEN_1378 : ~_GEN_2127 & _GEN_1378);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1377) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_19_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_19_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_19_bits_committed <=
      ~_GEN_2416
      & (commit_store_2 & _GEN_2320
         | (commit_store_1 ? _GEN_2272 | _GEN_2195 | _GEN_1238 : _GEN_2195 | _GEN_1238));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_19_bits_succeeded <=
      ~_GEN_2416
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h13
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h13))
         & _GEN_1214 & _GEN_1044 & _GEN_922 & stq_19_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_20_valid <=
      ~_GEN_2467 & (clear_store ? ~_GEN_2390 & _GEN_1188 : ~_GEN_2128 & _GEN_1188);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_20_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1215)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_20_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_923) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_20_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1021 | ~_GEN_923)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_20_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_20_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1215 & _GEN_1045 & _GEN_923 & stq_20_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h14
         | (_GEN_1215
              ? (_GEN_1045
                   ? (_GEN_923
                        ? stq_20_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923 ? stq_20_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1215
           ? (_GEN_1045
                ? (_GEN_923
                     ? stq_20_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_20_bits_addr_valid <=
      ~_GEN_2467 & (clear_store ? ~_GEN_2390 & _GEN_1332 : ~_GEN_2128 & _GEN_1332);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1331) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_20_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_20_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_20_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_20_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_20_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_20_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_20_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_20_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_20_bits_data_valid <=
      ~_GEN_2467 & (clear_store ? ~_GEN_2390 & _GEN_1380 : ~_GEN_2128 & _GEN_1380);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1379) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_20_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_20_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_20_bits_committed <=
      ~_GEN_2417
      & (commit_store_2 & _GEN_2321
         | (commit_store_1 ? _GEN_2273 | _GEN_2197 | _GEN_1239 : _GEN_2197 | _GEN_1239));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_20_bits_succeeded <=
      ~_GEN_2417
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h14
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h14))
         & _GEN_1215 & _GEN_1045 & _GEN_923 & stq_20_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_21_valid <=
      ~_GEN_2469 & (clear_store ? ~_GEN_2392 & _GEN_1190 : ~_GEN_2129 & _GEN_1190);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_21_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1216)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_21_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_924) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_21_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1022 | ~_GEN_924)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_21_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_21_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1216 & _GEN_1046 & _GEN_924 & stq_21_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h15
         | (_GEN_1216
              ? (_GEN_1046
                   ? (_GEN_924
                        ? stq_21_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924 ? stq_21_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1216
           ? (_GEN_1046
                ? (_GEN_924
                     ? stq_21_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_21_bits_addr_valid <=
      ~_GEN_2469 & (clear_store ? ~_GEN_2392 & _GEN_1334 : ~_GEN_2129 & _GEN_1334);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1333) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_21_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_21_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_21_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_21_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_21_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_21_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_21_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_21_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_21_bits_data_valid <=
      ~_GEN_2469 & (clear_store ? ~_GEN_2392 & _GEN_1382 : ~_GEN_2129 & _GEN_1382);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1381) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_21_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_21_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_21_bits_committed <=
      ~_GEN_2418
      & (commit_store_2 & _GEN_2322
         | (commit_store_1 ? _GEN_2274 | _GEN_2199 | _GEN_1240 : _GEN_2199 | _GEN_1240));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_21_bits_succeeded <=
      ~_GEN_2418
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h15
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h15))
         & _GEN_1216 & _GEN_1046 & _GEN_924 & stq_21_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_22_valid <=
      ~_GEN_2471 & (clear_store ? ~_GEN_2394 & _GEN_1192 : ~_GEN_2130 & _GEN_1192);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_22_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1217)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_22_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_925) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_22_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1023 | ~_GEN_925)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_22_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_22_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1217 & _GEN_1047 & _GEN_925 & stq_22_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h16
         | (_GEN_1217
              ? (_GEN_1047
                   ? (_GEN_925
                        ? stq_22_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925 ? stq_22_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1217
           ? (_GEN_1047
                ? (_GEN_925
                     ? stq_22_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_22_bits_addr_valid <=
      ~_GEN_2471 & (clear_store ? ~_GEN_2394 & _GEN_1336 : ~_GEN_2130 & _GEN_1336);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1335) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_22_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_22_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_22_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_22_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_22_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_22_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_22_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_22_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_22_bits_data_valid <=
      ~_GEN_2471 & (clear_store ? ~_GEN_2394 & _GEN_1384 : ~_GEN_2130 & _GEN_1384);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1383) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_22_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_22_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_22_bits_committed <=
      ~_GEN_2419
      & (commit_store_2 & _GEN_2323
         | (commit_store_1 ? _GEN_2275 | _GEN_2201 | _GEN_1241 : _GEN_2201 | _GEN_1241));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_22_bits_succeeded <=
      ~_GEN_2419
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h16
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h16))
         & _GEN_1217 & _GEN_1047 & _GEN_925 & stq_22_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_23_valid <=
      ~_GEN_2473 & (clear_store ? ~_GEN_2396 & _GEN_1194 : ~_GEN_2131 & _GEN_1194);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_23_bits_uop_is_rvc <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
                : io_core_dis_uops_1_bits_is_rvc)
           : io_core_dis_uops_2_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_ctrl_fcn_dw <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_ctrl_fcn_dw
                     : io_core_dis_uops_0_bits_ctrl_fcn_dw)
                : io_core_dis_uops_1_bits_ctrl_fcn_dw)
           : io_core_dis_uops_2_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_ctrl_is_load <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_ctrl_is_load
                     : io_core_dis_uops_0_bits_ctrl_is_load)
                : io_core_dis_uops_1_bits_ctrl_is_load)
           : io_core_dis_uops_2_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_ctrl_is_sta <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_ctrl_is_sta
                     : io_core_dis_uops_0_bits_ctrl_is_sta)
                : io_core_dis_uops_1_bits_ctrl_is_sta)
           : io_core_dis_uops_2_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_ctrl_is_std <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_ctrl_is_std
                     : io_core_dis_uops_0_bits_ctrl_is_std)
                : io_core_dis_uops_1_bits_ctrl_is_std)
           : io_core_dis_uops_2_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_iw_p1_poisoned <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_iw_p1_poisoned
                     : io_core_dis_uops_0_bits_iw_p1_poisoned)
                : io_core_dis_uops_1_bits_iw_p1_poisoned)
           : io_core_dis_uops_2_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_iw_p2_poisoned <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_iw_p2_poisoned
                     : io_core_dis_uops_0_bits_iw_p2_poisoned)
                : io_core_dis_uops_1_bits_iw_p2_poisoned)
           : io_core_dis_uops_2_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_br <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
                : io_core_dis_uops_1_bits_is_br)
           : io_core_dis_uops_2_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_jalr <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
                : io_core_dis_uops_1_bits_is_jalr)
           : io_core_dis_uops_2_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_jal <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
                : io_core_dis_uops_1_bits_is_jal)
           : io_core_dis_uops_2_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_sfb <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
                : io_core_dis_uops_1_bits_is_sfb)
           : io_core_dis_uops_2_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_edge_inst <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_edge_inst
                     : io_core_dis_uops_0_bits_edge_inst)
                : io_core_dis_uops_1_bits_edge_inst)
           : io_core_dis_uops_2_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_taken <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_taken : io_core_dis_uops_0_bits_taken)
                : io_core_dis_uops_1_bits_taken)
           : io_core_dis_uops_2_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    if (_GEN_2425 | ~_GEN_1218)	// lsu.scala:304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
      stq_23_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    else if (dis_ld_val_1) begin	// lsu.scala:301:85
      if (_GEN_926) begin	// lsu.scala:211:16, :304:5, :321:5
      end
      else	// lsu.scala:211:16, :304:5, :321:5
        stq_23_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    end
    else if (_GEN_1024 | ~_GEN_926)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
      stq_23_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
    stq_23_bits_uop_prs1_busy <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_prs1_busy
                     : io_core_dis_uops_0_bits_prs1_busy)
                : io_core_dis_uops_1_bits_prs1_busy)
           : io_core_dis_uops_2_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_prs2_busy <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_prs2_busy
                     : io_core_dis_uops_0_bits_prs2_busy)
                : io_core_dis_uops_1_bits_prs2_busy)
           : io_core_dis_uops_2_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_prs3_busy <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_prs3_busy
                     : io_core_dis_uops_0_bits_prs3_busy)
                : io_core_dis_uops_1_bits_prs3_busy)
           : io_core_dis_uops_2_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_ppred_busy <=
      ~_GEN_2425 & _GEN_1218 & _GEN_1048 & _GEN_926 & stq_23_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_exception <=
      ~_GEN_2425
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h17
         | (_GEN_1218
              ? (_GEN_1048
                   ? (_GEN_926
                        ? stq_23_bits_uop_exception
                        : io_core_dis_uops_0_bits_exception)
                   : io_core_dis_uops_1_bits_exception)
              : io_core_dis_uops_2_bits_exception));	// lsu.scala:211:16, :304:5, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32, util.scala:205:25
    stq_23_bits_uop_bypassable <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_bypassable
                     : io_core_dis_uops_0_bits_bypassable)
                : io_core_dis_uops_1_bits_bypassable)
           : io_core_dis_uops_2_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_mem_signed <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_mem_signed
                     : io_core_dis_uops_0_bits_mem_signed)
                : io_core_dis_uops_1_bits_mem_signed)
           : io_core_dis_uops_2_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_fence <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
                : io_core_dis_uops_1_bits_is_fence)
           : io_core_dis_uops_2_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_fencei <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_is_fencei
                     : io_core_dis_uops_0_bits_is_fencei)
                : io_core_dis_uops_1_bits_is_fencei)
           : io_core_dis_uops_2_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_amo <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
                : io_core_dis_uops_1_bits_is_amo)
           : io_core_dis_uops_2_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_uses_ldq <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
                : io_core_dis_uops_1_bits_uses_ldq)
           : io_core_dis_uops_2_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_uses_stq <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
                : io_core_dis_uops_1_bits_uses_stq)
           : io_core_dis_uops_2_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_sys_pc2epc <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_is_sys_pc2epc
                     : io_core_dis_uops_0_bits_is_sys_pc2epc)
                : io_core_dis_uops_1_bits_is_sys_pc2epc)
           : io_core_dis_uops_2_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_is_unique <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_is_unique
                     : io_core_dis_uops_0_bits_is_unique)
                : io_core_dis_uops_1_bits_is_unique)
           : io_core_dis_uops_2_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_flush_on_commit <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_flush_on_commit
                     : io_core_dis_uops_0_bits_flush_on_commit)
                : io_core_dis_uops_1_bits_flush_on_commit)
           : io_core_dis_uops_2_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_ldst_is_rs1 <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_ldst_is_rs1
                     : io_core_dis_uops_0_bits_ldst_is_rs1)
                : io_core_dis_uops_1_bits_ldst_is_rs1)
           : io_core_dis_uops_2_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_ldst_val <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
                : io_core_dis_uops_1_bits_ldst_val)
           : io_core_dis_uops_2_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_frs3_en <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
                : io_core_dis_uops_1_bits_frs3_en)
           : io_core_dis_uops_2_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_fp_val <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926 ? stq_23_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
                : io_core_dis_uops_1_bits_fp_val)
           : io_core_dis_uops_2_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_fp_single <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_fp_single
                     : io_core_dis_uops_0_bits_fp_single)
                : io_core_dis_uops_1_bits_fp_single)
           : io_core_dis_uops_2_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_xcpt_pf_if <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_xcpt_pf_if
                     : io_core_dis_uops_0_bits_xcpt_pf_if)
                : io_core_dis_uops_1_bits_xcpt_pf_if)
           : io_core_dis_uops_2_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_xcpt_ae_if <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_xcpt_ae_if
                     : io_core_dis_uops_0_bits_xcpt_ae_if)
                : io_core_dis_uops_1_bits_xcpt_ae_if)
           : io_core_dis_uops_2_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_xcpt_ma_if <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_xcpt_ma_if
                     : io_core_dis_uops_0_bits_xcpt_ma_if)
                : io_core_dis_uops_1_bits_xcpt_ma_if)
           : io_core_dis_uops_2_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_bp_debug_if <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_bp_debug_if
                     : io_core_dis_uops_0_bits_bp_debug_if)
                : io_core_dis_uops_1_bits_bp_debug_if)
           : io_core_dis_uops_2_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_uop_bp_xcpt_if <=
      ~_GEN_2425
      & (_GEN_1218
           ? (_GEN_1048
                ? (_GEN_926
                     ? stq_23_bits_uop_bp_xcpt_if
                     : io_core_dis_uops_0_bits_bp_xcpt_if)
                : io_core_dis_uops_1_bits_bp_xcpt_if)
           : io_core_dis_uops_2_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_23_bits_addr_valid <=
      ~_GEN_2473 & (clear_store ? ~_GEN_2396 & _GEN_1338 : ~_GEN_2131 & _GEN_1338);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_1337) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_23_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_23_bits_addr_bits <= _GEN_312;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_23_bits_addr_bits <= _GEN_199;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_23_bits_addr_bits <= _GEN_208;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_23_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_23_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_23_bits_addr_bits <= _GEN_313;	// lsu.scala:211:16, :768:30
      stq_23_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_23_bits_data_valid <=
      ~_GEN_2473 & (clear_store ? ~_GEN_2396 & _GEN_1386 : ~_GEN_2131 & _GEN_1386);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_1385) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_23_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_23_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_23_bits_committed <=
      ~_GEN_2420
      & (commit_store_2 & _GEN_2324
         | (commit_store_1 ? _GEN_2276 | _GEN_2203 | _GEN_1242 : _GEN_2203 | _GEN_1242));	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_23_bits_succeeded <=
      ~_GEN_2420
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h17
         | (_GEN_315 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h17))
         & _GEN_1218 & _GEN_1048 & _GEN_926 & stq_23_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35, util.scala:205:25
    if (_GEN_2424) begin	// lsu.scala:1596:22
      ldq_head <= 5'h0;	// lsu.scala:215:29
      ldq_tail <= 5'h0;	// lsu.scala:216:29
      if (reset)
        stq_tail <= 5'h0;	// lsu.scala:218:29
      else
        stq_tail <= stq_commit_head;	// lsu.scala:218:29, :219:29
    end
    else begin	// lsu.scala:1596:22
      if (commit_load_2) begin	// lsu.scala:1452:49
        if (_GEN_833 == 5'h17)	// lsu.scala:1486:31, util.scala:205:25
          ldq_head <= 5'h0;	// lsu.scala:215:29
        else	// util.scala:205:25
          ldq_head <= _GEN_833 + 5'h1;	// lsu.scala:215:29, :305:44, :1486:31, util.scala:206:28
      end
      else if (commit_load_1) begin	// lsu.scala:1452:49
        if (wrap_15)	// util.scala:205:25
          ldq_head <= 5'h0;	// lsu.scala:215:29
        else	// util.scala:205:25
          ldq_head <= _GEN_832;	// lsu.scala:215:29, util.scala:206:28
      end
      else if (commit_load) begin	// lsu.scala:1452:49
        if (wrap_13)	// util.scala:205:25
          ldq_head <= 5'h0;	// lsu.scala:215:29
        else	// util.scala:205:25
          ldq_head <= _GEN_828;	// lsu.scala:215:29, util.scala:206:28
      end
      if (io_core_brupdate_b2_mispredict & ~io_core_exception) begin	// lsu.scala:669:22, :1435:40
        ldq_tail <= io_core_brupdate_b2_uop_ldq_idx;	// lsu.scala:216:29
        stq_tail <= io_core_brupdate_b2_uop_stq_idx;	// lsu.scala:218:29
      end
      else begin	// lsu.scala:1435:40
        if (dis_ld_val_2) begin	// lsu.scala:301:85
          if (wrap_8)	// util.scala:205:25
            ldq_tail <= 5'h0;	// lsu.scala:216:29
          else	// util.scala:205:25
            ldq_tail <= _GEN_108;	// lsu.scala:216:29, util.scala:206:28
        end
        else if (dis_ld_val_1) begin	// lsu.scala:301:85
          if (wrap_4)	// util.scala:205:25
            ldq_tail <= 5'h0;	// lsu.scala:216:29
          else	// util.scala:205:25
            ldq_tail <= _GEN_102;	// lsu.scala:216:29, util.scala:206:28
        end
        else if (dis_ld_val) begin	// lsu.scala:301:85
          if (wrap)	// util.scala:205:25
            ldq_tail <= 5'h0;	// lsu.scala:216:29
          else	// util.scala:205:25
            ldq_tail <= _GEN_95;	// lsu.scala:216:29, util.scala:206:28
        end
        if (dis_st_val_2) begin	// lsu.scala:302:85
          if (wrap_9)	// util.scala:205:25
            stq_tail <= 5'h0;	// lsu.scala:218:29
          else	// util.scala:205:25
            stq_tail <= _GEN_109;	// lsu.scala:218:29, util.scala:206:28
        end
        else if (dis_st_val_1) begin	// lsu.scala:302:85
          if (wrap_5)	// util.scala:205:25
            stq_tail <= 5'h0;	// lsu.scala:218:29
          else	// util.scala:205:25
            stq_tail <= _GEN_104;	// lsu.scala:218:29, util.scala:206:28
        end
        else if (dis_st_val) begin	// lsu.scala:302:85
          if (wrap_1)	// util.scala:205:25
            stq_tail <= 5'h0;	// lsu.scala:218:29
          else	// util.scala:205:25
            stq_tail <= _GEN_97;	// lsu.scala:218:29, util.scala:206:28
        end
      end
    end
    if (_GEN_2422) begin	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
      hella_req_addr <= io_hellacache_req_bits_addr;	// lsu.scala:243:34
      hella_req_cmd <= 5'h0;	// lsu.scala:243:34
      hella_req_size <= 2'h3;	// lsu.scala:243:34
    end
    hella_req_signed <= ~_GEN_2422 & hella_req_signed;	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
    hella_req_phys <= _GEN_2422 | hella_req_phys;	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
    if (_GEN_2423)	// lsu.scala:244:34, :1527:34, :1533:38
      hella_data_data <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:244:34, :249:20
    if (can_fire_load_incoming_0 | will_fire_load_retry_0 | _GEN_316
        | ~will_fire_hella_incoming_0) begin	// lsu.scala:245:34, :441:63, :535:65, :766:39, :773:43, :780:45, :794:44, :802:47
    end
    else	// lsu.scala:245:34, :766:39, :773:43, :780:45, :794:44, :802:47
      hella_paddr <= exe_tlb_paddr_0;	// Cat.scala:30:58, lsu.scala:245:34
    if (_GEN_2423) begin	// lsu.scala:244:34, :246:34, :1527:34, :1533:38
      hella_xcpt_ma_ld <= _dtlb_io_resp_0_ma_ld;	// lsu.scala:246:34, :249:20
      hella_xcpt_ma_st <= _dtlb_io_resp_0_ma_st;	// lsu.scala:246:34, :249:20
      hella_xcpt_pf_ld <= _dtlb_io_resp_0_pf_ld;	// lsu.scala:246:34, :249:20
      hella_xcpt_pf_st <= _dtlb_io_resp_0_pf_st;	// lsu.scala:246:34, :249:20
      hella_xcpt_ae_ld <= _dtlb_io_resp_0_ae_ld;	// lsu.scala:246:34, :249:20
      hella_xcpt_ae_st <= _dtlb_io_resp_0_ae_st;	// lsu.scala:246:34, :249:20
    end
    if (will_fire_load_wakeup_0) begin	// lsu.scala:535:65
      p1_block_load_mask_0 <= _GEN_216;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_1 <= _GEN_217;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_2 <= _GEN_218;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_3 <= _GEN_219;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_4 <= _GEN_220;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_5 <= _GEN_221;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_6 <= _GEN_222;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_7 <= _GEN_223;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_8 <= _GEN_224;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_9 <= _GEN_225;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_10 <= _GEN_226;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_11 <= _GEN_227;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_12 <= _GEN_228;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_13 <= _GEN_229;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_14 <= _GEN_230;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_15 <= _GEN_231;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_16 <= _GEN_232;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_17 <= _GEN_233;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_18 <= _GEN_234;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_19 <= _GEN_235;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_20 <= _GEN_236;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_21 <= _GEN_237;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_22 <= _GEN_238;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_23 <= _GEN_239;	// lsu.scala:398:35, :570:49
    end
    else if (can_fire_load_incoming_0) begin	// lsu.scala:441:63
      p1_block_load_mask_0 <= _GEN_240;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_1 <= _GEN_241;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_2 <= _GEN_242;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_3 <= _GEN_243;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_4 <= _GEN_244;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_5 <= _GEN_245;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_6 <= _GEN_246;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_7 <= _GEN_247;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_8 <= _GEN_248;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_9 <= _GEN_249;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_10 <= _GEN_250;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_11 <= _GEN_251;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_12 <= _GEN_252;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_13 <= _GEN_253;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_14 <= _GEN_254;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_15 <= _GEN_255;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_16 <= _GEN_256;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_17 <= _GEN_257;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_18 <= _GEN_258;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_19 <= _GEN_259;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_20 <= _GEN_260;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_21 <= _GEN_261;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_22 <= _GEN_262;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_23 <= _GEN_263;	// lsu.scala:398:35, :572:52
    end
    else begin	// lsu.scala:441:63
      p1_block_load_mask_0 <= _GEN_265;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_1 <= _GEN_267;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_2 <= _GEN_269;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_3 <= _GEN_271;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_4 <= _GEN_273;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_5 <= _GEN_275;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_6 <= _GEN_277;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_7 <= _GEN_279;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_8 <= _GEN_281;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_9 <= _GEN_283;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_10 <= _GEN_285;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_11 <= _GEN_287;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_12 <= _GEN_289;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_13 <= _GEN_291;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_14 <= _GEN_293;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_15 <= _GEN_295;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_16 <= _GEN_297;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_17 <= _GEN_299;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_18 <= _GEN_301;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_19 <= _GEN_303;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_20 <= _GEN_305;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_21 <= _GEN_307;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_22 <= _GEN_309;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_23 <= _GEN_311;	// lsu.scala:398:35, :573:43, :574:49
    end
    p2_block_load_mask_0 <= p1_block_load_mask_0;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_1 <= p1_block_load_mask_1;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_2 <= p1_block_load_mask_2;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_3 <= p1_block_load_mask_3;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_4 <= p1_block_load_mask_4;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_5 <= p1_block_load_mask_5;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_6 <= p1_block_load_mask_6;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_7 <= p1_block_load_mask_7;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_8 <= p1_block_load_mask_8;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_9 <= p1_block_load_mask_9;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_10 <= p1_block_load_mask_10;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_11 <= p1_block_load_mask_11;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_12 <= p1_block_load_mask_12;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_13 <= p1_block_load_mask_13;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_14 <= p1_block_load_mask_14;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_15 <= p1_block_load_mask_15;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_16 <= p1_block_load_mask_16;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_17 <= p1_block_load_mask_17;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_18 <= p1_block_load_mask_18;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_19 <= p1_block_load_mask_19;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_20 <= p1_block_load_mask_20;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_21 <= p1_block_load_mask_21;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_22 <= p1_block_load_mask_22;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_23 <= p1_block_load_mask_23;	// lsu.scala:398:35, :399:35
    _ldq_retry_idx_idx_T_34 =
      _ldq_retry_idx_T_62 & _temp_bits_T_40
        ? 6'h14
        : _ldq_retry_idx_T_65 & _temp_bits_T_42
            ? 6'h15
            : _ldq_retry_idx_T_68 & _temp_bits_T_44
                ? 6'h16
                : ldq_23_bits_addr_valid & ldq_23_bits_addr_is_virtual
                  & ~ldq_retry_idx_block_23 & _temp_bits_T_46
                    ? 6'h17
                    : _ldq_retry_idx_T_2
                        ? 6'h20
                        : _ldq_retry_idx_T_5
                            ? 6'h21
                            : _ldq_retry_idx_T_8
                                ? 6'h22
                                : _ldq_retry_idx_T_11
                                    ? 6'h23
                                    : _ldq_retry_idx_T_14
                                        ? 6'h24
                                        : _ldq_retry_idx_T_17
                                            ? 6'h25
                                            : _ldq_retry_idx_T_20
                                                ? 6'h26
                                                : _ldq_retry_idx_T_23
                                                    ? 6'h27
                                                    : _ldq_retry_idx_T_26
                                                        ? 6'h28
                                                        : _ldq_retry_idx_T_29
                                                            ? 6'h29
                                                            : _ldq_retry_idx_T_32
                                                                ? 6'h2A
                                                                : _ldq_retry_idx_T_35
                                                                    ? 6'h2B
                                                                    : _ldq_retry_idx_T_38
                                                                        ? 6'h2C
                                                                        : _ldq_retry_idx_T_41
                                                                            ? 6'h2D
                                                                            : _ldq_retry_idx_T_44
                                                                                ? 6'h2E
                                                                                : _ldq_retry_idx_T_47
                                                                                    ? 6'h2F
                                                                                    : _ldq_retry_idx_T_50
                                                                                        ? 6'h30
                                                                                        : _ldq_retry_idx_T_53
                                                                                            ? 6'h31
                                                                                            : _ldq_retry_idx_T_56
                                                                                                ? 6'h32
                                                                                                : _ldq_retry_idx_T_59
                                                                                                    ? 6'h33
                                                                                                    : _ldq_retry_idx_T_62
                                                                                                        ? 6'h34
                                                                                                        : _ldq_retry_idx_T_65
                                                                                                            ? 6'h35
                                                                                                            : {5'h1B,
                                                                                                               ~_ldq_retry_idx_T_68};	// Mux.scala:47:69, lsu.scala:210:16, :417:36, :418:{39,42}, util.scala:351:{65,72}
    ldq_retry_idx <=
      _ldq_retry_idx_T_2 & _temp_bits_T
        ? 5'h0
        : _ldq_retry_idx_T_5 & _temp_bits_T_2
            ? 5'h1
            : _ldq_retry_idx_T_8 & _temp_bits_T_4
                ? 5'h2
                : _ldq_retry_idx_T_11 & _temp_bits_T_6
                    ? 5'h3
                    : _ldq_retry_idx_T_14 & _temp_bits_T_8
                        ? 5'h4
                        : _ldq_retry_idx_T_17 & _temp_bits_T_10
                            ? 5'h5
                            : _ldq_retry_idx_T_20 & _temp_bits_T_12
                                ? 5'h6
                                : _ldq_retry_idx_T_23 & _temp_bits_T_14
                                    ? 5'h7
                                    : _ldq_retry_idx_T_26 & _temp_bits_T_16
                                        ? 5'h8
                                        : _ldq_retry_idx_T_29 & _temp_bits_T_18
                                            ? 5'h9
                                            : _ldq_retry_idx_T_32 & _temp_bits_T_20
                                                ? 5'hA
                                                : _ldq_retry_idx_T_35 & _temp_bits_T_22
                                                    ? 5'hB
                                                    : _ldq_retry_idx_T_38
                                                      & _temp_bits_T_24
                                                        ? 5'hC
                                                        : _ldq_retry_idx_T_41
                                                          & _temp_bits_T_26
                                                            ? 5'hD
                                                            : _ldq_retry_idx_T_44
                                                              & _temp_bits_T_28
                                                                ? 5'hE
                                                                : _ldq_retry_idx_T_47
                                                                  & ~(ldq_head[4])
                                                                    ? 5'hF
                                                                    : _ldq_retry_idx_T_50
                                                                      & _temp_bits_T_32
                                                                        ? 5'h10
                                                                        : _ldq_retry_idx_T_53
                                                                          & _temp_bits_T_34
                                                                            ? 5'h11
                                                                            : _ldq_retry_idx_T_56
                                                                              & _temp_bits_T_36
                                                                                ? 5'h12
                                                                                : _ldq_retry_idx_T_59
                                                                                  & _temp_bits_T_38
                                                                                    ? 5'h13
                                                                                    : _ldq_retry_idx_idx_T_34[4:0];	// Mux.scala:47:69, lsu.scala:215:29, :305:44, :415:30, :418:39, util.scala:351:{65,72}
    _stq_retry_idx_idx_T_34 =
      _stq_retry_idx_T_20 & stq_commit_head < 5'h15
        ? 6'h14
        : _stq_retry_idx_T_21 & stq_commit_head < 5'h16
            ? 6'h15
            : _stq_retry_idx_T_22 & stq_commit_head < 5'h17
                ? 6'h16
                : stq_23_bits_addr_valid & stq_23_bits_addr_is_virtual
                  & stq_commit_head[4:3] != 2'h3
                    ? 6'h17
                    : _stq_retry_idx_T
                        ? 6'h20
                        : _stq_retry_idx_T_1
                            ? 6'h21
                            : _stq_retry_idx_T_2
                                ? 6'h22
                                : _stq_retry_idx_T_3
                                    ? 6'h23
                                    : _stq_retry_idx_T_4
                                        ? 6'h24
                                        : _stq_retry_idx_T_5
                                            ? 6'h25
                                            : _stq_retry_idx_T_6
                                                ? 6'h26
                                                : _stq_retry_idx_T_7
                                                    ? 6'h27
                                                    : _stq_retry_idx_T_8
                                                        ? 6'h28
                                                        : _stq_retry_idx_T_9
                                                            ? 6'h29
                                                            : _stq_retry_idx_T_10
                                                                ? 6'h2A
                                                                : _stq_retry_idx_T_11
                                                                    ? 6'h2B
                                                                    : _stq_retry_idx_T_12
                                                                        ? 6'h2C
                                                                        : _stq_retry_idx_T_13
                                                                            ? 6'h2D
                                                                            : _stq_retry_idx_T_14
                                                                                ? 6'h2E
                                                                                : _stq_retry_idx_T_15
                                                                                    ? 6'h2F
                                                                                    : _stq_retry_idx_T_16
                                                                                        ? 6'h30
                                                                                        : _stq_retry_idx_T_17
                                                                                            ? 6'h31
                                                                                            : _stq_retry_idx_T_18
                                                                                                ? 6'h32
                                                                                                : _stq_retry_idx_T_19
                                                                                                    ? 6'h33
                                                                                                    : _stq_retry_idx_T_20
                                                                                                        ? 6'h34
                                                                                                        : _stq_retry_idx_T_21
                                                                                                            ? 6'h35
                                                                                                            : {5'h1B,
                                                                                                               ~_stq_retry_idx_T_22};	// Mux.scala:47:69, lsu.scala:211:16, :219:29, :305:44, :424:18, util.scala:205:25, :351:{65,72}
    stq_retry_idx <=
      _stq_retry_idx_T & stq_commit_head == 5'h0
        ? 5'h0
        : _stq_retry_idx_T_1 & stq_commit_head < 5'h2
            ? 5'h1
            : _stq_retry_idx_T_2 & stq_commit_head < 5'h3
                ? 5'h2
                : _stq_retry_idx_T_3 & stq_commit_head < 5'h4
                    ? 5'h3
                    : _stq_retry_idx_T_4 & stq_commit_head < 5'h5
                        ? 5'h4
                        : _stq_retry_idx_T_5 & stq_commit_head < 5'h6
                            ? 5'h5
                            : _stq_retry_idx_T_6 & stq_commit_head < 5'h7
                                ? 5'h6
                                : _stq_retry_idx_T_7 & stq_commit_head < 5'h8
                                    ? 5'h7
                                    : _stq_retry_idx_T_8 & stq_commit_head < 5'h9
                                        ? 5'h8
                                        : _stq_retry_idx_T_9 & stq_commit_head < 5'hA
                                            ? 5'h9
                                            : _stq_retry_idx_T_10 & stq_commit_head < 5'hB
                                                ? 5'hA
                                                : _stq_retry_idx_T_11
                                                  & stq_commit_head < 5'hC
                                                    ? 5'hB
                                                    : _stq_retry_idx_T_12
                                                      & stq_commit_head < 5'hD
                                                        ? 5'hC
                                                        : _stq_retry_idx_T_13
                                                          & stq_commit_head < 5'hE
                                                            ? 5'hD
                                                            : _stq_retry_idx_T_14
                                                              & stq_commit_head < 5'hF
                                                                ? 5'hE
                                                                : _stq_retry_idx_T_15
                                                                  & ~(stq_commit_head[4])
                                                                    ? 5'hF
                                                                    : _stq_retry_idx_T_16
                                                                      & stq_commit_head < 5'h11
                                                                        ? 5'h10
                                                                        : _stq_retry_idx_T_17
                                                                          & stq_commit_head < 5'h12
                                                                            ? 5'h11
                                                                            : _stq_retry_idx_T_18
                                                                              & stq_commit_head < 5'h13
                                                                                ? 5'h12
                                                                                : _stq_retry_idx_T_19
                                                                                  & stq_commit_head < 5'h14
                                                                                    ? 5'h13
                                                                                    : _stq_retry_idx_idx_T_34[4:0];	// Mux.scala:47:69, lsu.scala:219:29, :305:44, :422:30, :424:18, util.scala:351:{65,72}
    _ldq_wakeup_idx_idx_T_34 =
      _ldq_wakeup_idx_T_167 & _temp_bits_T_40
        ? 6'h14
        : _ldq_wakeup_idx_T_175 & _temp_bits_T_42
            ? 6'h15
            : _ldq_wakeup_idx_T_183 & _temp_bits_T_44
                ? 6'h16
                : ldq_23_bits_addr_valid & ~ldq_23_bits_executed & ~ldq_23_bits_succeeded
                  & ~ldq_23_bits_addr_is_virtual & ~ldq_retry_idx_block_23
                  & _temp_bits_T_46
                    ? 6'h17
                    : _ldq_wakeup_idx_T_7
                        ? 6'h20
                        : _ldq_wakeup_idx_T_15
                            ? 6'h21
                            : _ldq_wakeup_idx_T_23
                                ? 6'h22
                                : _ldq_wakeup_idx_T_31
                                    ? 6'h23
                                    : _ldq_wakeup_idx_T_39
                                        ? 6'h24
                                        : _ldq_wakeup_idx_T_47
                                            ? 6'h25
                                            : _ldq_wakeup_idx_T_55
                                                ? 6'h26
                                                : _ldq_wakeup_idx_T_63
                                                    ? 6'h27
                                                    : _ldq_wakeup_idx_T_71
                                                        ? 6'h28
                                                        : _ldq_wakeup_idx_T_79
                                                            ? 6'h29
                                                            : _ldq_wakeup_idx_T_87
                                                                ? 6'h2A
                                                                : _ldq_wakeup_idx_T_95
                                                                    ? 6'h2B
                                                                    : _ldq_wakeup_idx_T_103
                                                                        ? 6'h2C
                                                                        : _ldq_wakeup_idx_T_111
                                                                            ? 6'h2D
                                                                            : _ldq_wakeup_idx_T_119
                                                                                ? 6'h2E
                                                                                : _ldq_wakeup_idx_T_127
                                                                                    ? 6'h2F
                                                                                    : _ldq_wakeup_idx_T_135
                                                                                        ? 6'h30
                                                                                        : _ldq_wakeup_idx_T_143
                                                                                            ? 6'h31
                                                                                            : _ldq_wakeup_idx_T_151
                                                                                                ? 6'h32
                                                                                                : _ldq_wakeup_idx_T_159
                                                                                                    ? 6'h33
                                                                                                    : _ldq_wakeup_idx_T_167
                                                                                                        ? 6'h34
                                                                                                        : _ldq_wakeup_idx_T_175
                                                                                                            ? 6'h35
                                                                                                            : {5'h1B,
                                                                                                               ~_ldq_wakeup_idx_T_183};	// Mux.scala:47:69, lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}, util.scala:351:{65,72}
    ldq_wakeup_idx <=
      _ldq_wakeup_idx_T_7 & _temp_bits_T
        ? 5'h0
        : _ldq_wakeup_idx_T_15 & _temp_bits_T_2
            ? 5'h1
            : _ldq_wakeup_idx_T_23 & _temp_bits_T_4
                ? 5'h2
                : _ldq_wakeup_idx_T_31 & _temp_bits_T_6
                    ? 5'h3
                    : _ldq_wakeup_idx_T_39 & _temp_bits_T_8
                        ? 5'h4
                        : _ldq_wakeup_idx_T_47 & _temp_bits_T_10
                            ? 5'h5
                            : _ldq_wakeup_idx_T_55 & _temp_bits_T_12
                                ? 5'h6
                                : _ldq_wakeup_idx_T_63 & _temp_bits_T_14
                                    ? 5'h7
                                    : _ldq_wakeup_idx_T_71 & _temp_bits_T_16
                                        ? 5'h8
                                        : _ldq_wakeup_idx_T_79 & _temp_bits_T_18
                                            ? 5'h9
                                            : _ldq_wakeup_idx_T_87 & _temp_bits_T_20
                                                ? 5'hA
                                                : _ldq_wakeup_idx_T_95 & _temp_bits_T_22
                                                    ? 5'hB
                                                    : _ldq_wakeup_idx_T_103
                                                      & _temp_bits_T_24
                                                        ? 5'hC
                                                        : _ldq_wakeup_idx_T_111
                                                          & _temp_bits_T_26
                                                            ? 5'hD
                                                            : _ldq_wakeup_idx_T_119
                                                              & _temp_bits_T_28
                                                                ? 5'hE
                                                                : _ldq_wakeup_idx_T_127
                                                                  & ~(ldq_head[4])
                                                                    ? 5'hF
                                                                    : _ldq_wakeup_idx_T_135
                                                                      & _temp_bits_T_32
                                                                        ? 5'h10
                                                                        : _ldq_wakeup_idx_T_143
                                                                          & _temp_bits_T_34
                                                                            ? 5'h11
                                                                            : _ldq_wakeup_idx_T_151
                                                                              & _temp_bits_T_36
                                                                                ? 5'h12
                                                                                : _ldq_wakeup_idx_T_159
                                                                                  & _temp_bits_T_38
                                                                                    ? 5'h13
                                                                                    : _ldq_wakeup_idx_idx_T_34[4:0];	// Mux.scala:47:69, lsu.scala:215:29, :305:44, :430:31, :433:71, util.scala:351:{65,72}
    can_fire_load_retry_REG <= _dtlb_io_miss_rdy;	// lsu.scala:249:20, :470:40
    can_fire_sta_retry_REG <= _dtlb_io_miss_rdy;	// lsu.scala:249:20, :482:41
    mem_xcpt_valids_0 <=
      (pf_ld_0 | pf_st_0 | ae_ld_0 | ~_will_fire_store_commit_0_T_2
       & _dtlb_io_resp_0_ae_st & _mem_xcpt_uops_WIRE_0_uses_stq | ma_ld_0 | ma_st_0)
      & ~io_core_exception
      & (io_core_brupdate_b1_mispredict_mask & exe_tlb_uop_0_br_mask) == 16'h0;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :659:56, :660:87, :661:75, :662:75, :663:75, :664:75, :667:32, :668:80, :669:{22,41}, util.scala:118:{51,59}
    mem_xcpt_uops_0_br_mask <= exe_tlb_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:597:24, :671:32, util.scala:85:{25,27}
    if (_exe_tlb_uop_T_2) begin	// lsu.scala:599:53
      mem_xcpt_uops_0_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;	// lsu.scala:671:32
      mem_xcpt_uops_0_ldq_idx <= io_core_exe_0_req_bits_uop_ldq_idx;	// lsu.scala:671:32
      mem_xcpt_uops_0_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;	// lsu.scala:671:32
      mem_xcpt_uops_0_uses_ldq <= io_core_exe_0_req_bits_uop_uses_ldq;	// lsu.scala:671:32
      mem_xcpt_uops_0_uses_stq <= io_core_exe_0_req_bits_uop_uses_stq;	// lsu.scala:671:32
    end
    else if (will_fire_load_retry_0) begin	// lsu.scala:535:65
      mem_xcpt_uops_0_rob_idx <= _GEN_149;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_ldq_idx <= _GEN_151;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_stq_idx <= mem_ldq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_uses_ldq <= _GEN_173;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_uses_stq <= _GEN_175;	// lsu.scala:465:79, :671:32
    end
    else begin	// lsu.scala:535:65
      if (will_fire_sta_retry_0) begin	// lsu.scala:536:61
        mem_xcpt_uops_0_rob_idx <= mem_stq_retry_e_out_bits_uop_rob_idx;	// lsu.scala:478:79, :671:32
        mem_xcpt_uops_0_ldq_idx <= _GEN_206;	// lsu.scala:478:79, :671:32
        mem_xcpt_uops_0_stq_idx <= mem_stq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:478:79, :671:32
      end
      else begin	// lsu.scala:536:61
        mem_xcpt_uops_0_rob_idx <= 7'h0;	// lsu.scala:671:32
        mem_xcpt_uops_0_ldq_idx <= 5'h0;	// lsu.scala:671:32
        mem_xcpt_uops_0_stq_idx <= 5'h0;	// lsu.scala:671:32
      end
      mem_xcpt_uops_0_uses_ldq <= _exe_tlb_uop_T_4_uses_ldq;	// lsu.scala:602:24, :671:32
      mem_xcpt_uops_0_uses_stq <= _exe_tlb_uop_T_4_uses_stq;	// lsu.scala:602:24, :671:32
    end
    if (ma_ld_0)	// lsu.scala:659:56
      mem_xcpt_causes_0 <= 4'h4;	// lsu.scala:672:32, :673:8
    else if (ma_st_0)	// lsu.scala:660:87
      mem_xcpt_causes_0 <= 4'h6;	// lsu.scala:672:32, :674:8
    else if (pf_ld_0)	// lsu.scala:661:75
      mem_xcpt_causes_0 <= 4'hD;	// lsu.scala:672:32, util.scala:351:72
    else if (pf_st_0)	// lsu.scala:662:75
      mem_xcpt_causes_0 <= 4'hF;	// lsu.scala:672:32, util.scala:351:72
    else	// lsu.scala:662:75
      mem_xcpt_causes_0 <= {2'h1, ~ae_ld_0, 1'h1};	// lsu.scala:249:20, :663:75, :672:32, :676:8, :677:8, :1312:58
    if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
      mem_xcpt_vaddrs_0 <= io_core_exe_0_req_bits_addr;	// lsu.scala:679:32
    else if (will_fire_sfence_0)	// lsu.scala:536:61
      mem_xcpt_vaddrs_0 <= _GEN_312;	// lsu.scala:610:24, :679:32
    else if (will_fire_load_retry_0)	// lsu.scala:535:65
      mem_xcpt_vaddrs_0 <= _GEN_199;	// lsu.scala:465:79, :679:32
    else if (will_fire_sta_retry_0)	// lsu.scala:536:61
      mem_xcpt_vaddrs_0 <= _GEN_208;	// lsu.scala:478:79, :679:32
    else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
      mem_xcpt_vaddrs_0 <= hella_req_addr;	// lsu.scala:243:34, :679:32
    else	// lsu.scala:535:65
      mem_xcpt_vaddrs_0 <= 40'h0;	// lsu.scala:679:32
    REG <= _GEN_215 | will_fire_load_retry_0 | will_fire_sta_retry_0;	// lsu.scala:535:65, :536:61, :567:93, :718:21, :719:33
    fired_load_incoming_REG <= can_fire_load_incoming_0 & _fired_std_incoming_T;	// lsu.scala:441:63, :894:{51,79}, util.scala:118:59
    fired_stad_incoming_REG <= will_fire_stad_incoming_0 & _fired_std_incoming_T;	// lsu.scala:534:63, :895:{51,79}, util.scala:118:59
    fired_sta_incoming_REG <= will_fire_sta_incoming_0 & _fired_std_incoming_T;	// lsu.scala:536:61, :896:{51,79}, util.scala:118:59
    fired_std_incoming_REG <= will_fire_std_incoming_0 & _fired_std_incoming_T;	// lsu.scala:536:61, :897:{51,79}, util.scala:118:59
    fired_stdf_incoming <=
      fp_stdata_fire
      & (io_core_brupdate_b1_mispredict_mask
         & io_core_fp_stdata_bits_uop_br_mask) == 16'h0;	// Decoupled.scala:40:37, lsu.scala:898:{37,62}, util.scala:118:{51,59}
    fired_sfence_0 <= will_fire_sfence_0;	// lsu.scala:536:61, :899:37
    fired_release_0 <= will_fire_release_0;	// lsu.scala:534:63, :900:37
    fired_load_retry_REG <=
      will_fire_load_retry_0 & (io_core_brupdate_b1_mispredict_mask & _GEN_140) == 16'h0;	// lsu.scala:465:79, :535:65, :901:{51,79}, util.scala:118:{51,59}
    fired_sta_retry_REG <= will_fire_sta_retry_0 & _mem_stq_retry_e_out_valid_T == 16'h0;	// lsu.scala:536:61, :902:{51,79}, util.scala:118:{51,59}
    fired_load_wakeup_REG <=
      will_fire_load_wakeup_0 & (io_core_brupdate_b1_mispredict_mask & _GEN_209) == 16'h0;	// lsu.scala:502:88, :535:65, :904:{51,79}, util.scala:118:{51,59}
    mem_incoming_uop_0_br_mask <=
      io_core_exe_0_req_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:908:37, util.scala:85:{25,27}
    mem_incoming_uop_0_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;	// lsu.scala:908:37
    mem_incoming_uop_0_ldq_idx <= io_core_exe_0_req_bits_uop_ldq_idx;	// lsu.scala:908:37
    mem_incoming_uop_0_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;	// lsu.scala:908:37
    mem_incoming_uop_0_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:908:37
    mem_incoming_uop_0_fp_val <= io_core_exe_0_req_bits_uop_fp_val;	// lsu.scala:908:37
    mem_ldq_incoming_e_0_bits_uop_br_mask <=
      _GEN_110[io_core_exe_0_req_bits_uop_ldq_idx] & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:264:49, :909:37, util.scala:85:27, :89:21
    mem_ldq_incoming_e_0_bits_uop_stq_idx <= _GEN_111[io_core_exe_0_req_bits_uop_ldq_idx];	// lsu.scala:264:49, :909:37
    mem_ldq_incoming_e_0_bits_uop_mem_size <=
      _GEN_112[io_core_exe_0_req_bits_uop_ldq_idx];	// lsu.scala:264:49, :909:37
    mem_ldq_incoming_e_0_bits_st_dep_mask <= _GEN_115[io_core_exe_0_req_bits_uop_ldq_idx];	// lsu.scala:264:49, :909:37
    mem_stq_incoming_e_0_valid <=
      _GEN_2[io_core_exe_0_req_bits_uop_stq_idx]
      & (io_core_brupdate_b1_mispredict_mask
         & _GEN_28[io_core_exe_0_req_bits_uop_stq_idx]) == 16'h0;	// lsu.scala:224:42, :264:49, :910:37, util.scala:108:31, :118:{51,59}
    mem_stq_incoming_e_0_bits_uop_br_mask <=
      _GEN_28[io_core_exe_0_req_bits_uop_stq_idx] & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:224:42, :264:49, :910:37, util.scala:85:27, :89:21
    mem_stq_incoming_e_0_bits_uop_rob_idx <= _GEN_36[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_uop_stq_idx <= _GEN_38[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_uop_mem_size <= _GEN_55[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_uop_is_amo <= _GEN_61[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_addr_valid <= _GEN_87[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_addr_is_virtual <=
      _GEN_90[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_data_valid <= _GEN_91[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_ldq_wakeup_e_bits_uop_br_mask <= _GEN_209 & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:502:88, :911:37, util.scala:85:27, :89:21
    mem_ldq_wakeup_e_bits_uop_stq_idx <= mem_ldq_wakeup_e_out_bits_uop_stq_idx;	// lsu.scala:502:88, :911:37
    mem_ldq_wakeup_e_bits_uop_mem_size <= mem_ldq_wakeup_e_out_bits_uop_mem_size;	// lsu.scala:502:88, :911:37
    mem_ldq_wakeup_e_bits_st_dep_mask <= mem_ldq_wakeup_e_out_bits_st_dep_mask;	// lsu.scala:502:88, :911:37
    mem_ldq_retry_e_bits_uop_br_mask <= _GEN_140 & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:465:79, :912:37, util.scala:85:27, :89:21
    mem_ldq_retry_e_bits_uop_stq_idx <= mem_ldq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:465:79, :912:37
    mem_ldq_retry_e_bits_uop_mem_size <= mem_ldq_retry_e_out_bits_uop_mem_size;	// lsu.scala:465:79, :912:37
    mem_ldq_retry_e_bits_st_dep_mask <= _GEN_115[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79, :912:37
    mem_stq_retry_e_valid <= _GEN_204 & _mem_stq_retry_e_out_valid_T == 16'h0;	// lsu.scala:478:79, :913:37, util.scala:108:31, :118:{51,59}
    mem_stq_retry_e_bits_uop_br_mask <= _GEN_205 & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:478:79, :913:37, util.scala:85:27, :89:21
    mem_stq_retry_e_bits_uop_rob_idx <= mem_stq_retry_e_out_bits_uop_rob_idx;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_uop_stq_idx <= mem_stq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_uop_mem_size <= mem_stq_retry_e_out_bits_uop_mem_size;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_uop_is_amo <= mem_stq_retry_e_out_bits_uop_is_amo;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_data_valid <= _GEN_91[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79, :913:37
    mem_stdf_uop_br_mask <=
      io_core_fp_stdata_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:922:37, util.scala:85:{25,27}
    mem_stdf_uop_rob_idx <= io_core_fp_stdata_bits_uop_rob_idx;	// lsu.scala:922:37
    mem_stdf_uop_stq_idx <= io_core_fp_stdata_bits_uop_stq_idx;	// lsu.scala:922:37
    mem_tlb_miss_0 <= exe_tlb_miss_0;	// lsu.scala:708:58, :925:41
    mem_tlb_uncacheable_0 <= ~_dtlb_io_resp_0_cacheable;	// lsu.scala:249:20, :711:43, :926:41
    if (_GEN_318)	// lsu.scala:766:39, :768:30, :773:43
      mem_paddr_0 <= _GEN_313;	// lsu.scala:768:30, :927:41
    else if (will_fire_store_commit_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_89;	// lsu.scala:224:42, :927:41
    else if (will_fire_load_wakeup_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_210;	// lsu.scala:502:88, :927:41
    else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_313;	// lsu.scala:768:30, :927:41
    else if (will_fire_hella_wakeup_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_317;	// lsu.scala:822:39, :927:41
    else	// lsu.scala:535:65
      mem_paddr_0 <= 40'h0;	// lsu.scala:927:41
    if (fired_stad_incoming_REG | fired_sta_incoming_REG | fired_std_incoming_REG)	// lsu.scala:895:51, :896:51, :897:51, :940:35, :945:27, :947:41, :953:27, :955:41, :961:27, :963:35
      clr_bsy_rob_idx_0 <= mem_stq_incoming_e_0_bits_uop_rob_idx;	// lsu.scala:910:37, :931:28
    else if (fired_sfence_0)	// lsu.scala:899:37
      clr_bsy_rob_idx_0 <= mem_incoming_uop_0_rob_idx;	// lsu.scala:908:37, :931:28
    else if (fired_sta_retry_REG)	// lsu.scala:902:51
      clr_bsy_rob_idx_0 <= mem_stq_retry_e_bits_uop_rob_idx;	// lsu.scala:913:37, :931:28
    else	// lsu.scala:902:51
      clr_bsy_rob_idx_0 <= 7'h0;	// lsu.scala:931:28
    if (fired_stad_incoming_REG)	// lsu.scala:895:51
      clr_bsy_brmask_0 <=
        mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:910:37, :932:28, util.scala:85:{25,27}
    else if (fired_sta_incoming_REG)	// lsu.scala:896:51
      clr_bsy_brmask_0 <=
        mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:910:37, :932:28, util.scala:85:{25,27}
    else if (fired_std_incoming_REG)	// lsu.scala:897:51
      clr_bsy_brmask_0 <=
        mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:910:37, :932:28, util.scala:85:{25,27}
    else if (fired_sfence_0)	// lsu.scala:899:37
      clr_bsy_brmask_0 <= mem_incoming_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:908:37, :932:28, util.scala:85:{25,27}
    else if (fired_sta_retry_REG)	// lsu.scala:902:51
      clr_bsy_brmask_0 <=
        mem_stq_retry_e_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:913:37, :932:28, util.scala:85:{25,27}
    else	// lsu.scala:902:51
      clr_bsy_brmask_0 <= 16'h0;	// lsu.scala:932:28
    io_core_clr_bsy_0_valid_REG <= io_core_exception;	// lsu.scala:979:62
    io_core_clr_bsy_0_valid_REG_1 <= io_core_exception;	// lsu.scala:979:101
    io_core_clr_bsy_0_valid_REG_2 <= io_core_clr_bsy_0_valid_REG_1;	// lsu.scala:979:{93,101}
    if (fired_stdf_incoming) begin	// lsu.scala:898:37
      stdf_clr_bsy_rob_idx <= mem_stdf_uop_rob_idx;	// lsu.scala:922:37, :984:33
      stdf_clr_bsy_brmask <= mem_stdf_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:922:37, :985:33, util.scala:85:{25,27}
    end
    else begin	// lsu.scala:898:37
      stdf_clr_bsy_rob_idx <= 7'h0;	// lsu.scala:984:33
      stdf_clr_bsy_brmask <= 16'h0;	// lsu.scala:985:33
    end
    io_core_clr_bsy_1_valid_REG <= io_core_exception;	// lsu.scala:1004:67
    io_core_clr_bsy_1_valid_REG_1 <= io_core_exception;	// lsu.scala:1004:106
    io_core_clr_bsy_1_valid_REG_2 <= io_core_clr_bsy_1_valid_REG_1;	// lsu.scala:1004:{98,106}
    lcam_addr_REG <= exe_tlb_paddr_0;	// Cat.scala:30:58, lsu.scala:1026:45
    lcam_addr_REG_1 <= io_dmem_release_bits_address;	// lsu.scala:1027:67
    lcam_ldq_idx_REG <= ldq_wakeup_idx;	// lsu.scala:430:31, :1037:58
    lcam_ldq_idx_REG_1 <= ldq_retry_idx;	// lsu.scala:415:30, :1038:58
    lcam_stq_idx_REG <= stq_retry_idx;	// lsu.scala:422:30, :1042:58
    if (can_fire_load_incoming_0) begin	// lsu.scala:441:63
      s1_executing_loads_0 <= _GEN_240 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_1 <= _GEN_241 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_2 <= _GEN_242 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_3 <= _GEN_243 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_4 <= _GEN_244 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_5 <= _GEN_245 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_6 <= _GEN_246 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_7 <= _GEN_247 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_8 <= _GEN_248 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_9 <= _GEN_249 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_10 <= _GEN_250 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_11 <= _GEN_251 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_12 <= _GEN_252 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_13 <= _GEN_253 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_14 <= _GEN_254 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_15 <= _GEN_255 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_16 <= _GEN_256 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_17 <= _GEN_257 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_18 <= _GEN_258 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_19 <= _GEN_259 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_20 <= _GEN_260 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_21 <= _GEN_261 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_22 <= _GEN_262 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_23 <= _GEN_263 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
    end
    else if (will_fire_load_retry_0) begin	// lsu.scala:535:65
      s1_executing_loads_0 <= _GEN_264 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_1 <= _GEN_266 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_2 <= _GEN_268 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_3 <= _GEN_270 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_4 <= _GEN_272 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_5 <= _GEN_274 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_6 <= _GEN_276 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_7 <= _GEN_278 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_8 <= _GEN_280 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_9 <= _GEN_282 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_10 <= _GEN_284 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_11 <= _GEN_286 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_12 <= _GEN_288 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_13 <= _GEN_290 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_14 <= _GEN_292 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_15 <= _GEN_294 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_16 <= _GEN_296 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_17 <= _GEN_298 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_18 <= _GEN_300 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_19 <= _GEN_302 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_20 <= _GEN_304 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_21 <= _GEN_306 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_22 <= _GEN_308 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_23 <= _GEN_310 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
    end
    else begin	// lsu.scala:535:65
      s1_executing_loads_0 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_216 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_1 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_217 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_2 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_218 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_3 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_219 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_4 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_220 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_5 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_221 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_6 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_222 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_7 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_223 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_8 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_224 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_9 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_225 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_10 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_226 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_11 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_227 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_12 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_228 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_13 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_229 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_14 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_230 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_15 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_231 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_16 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_232 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_17 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_233 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_18 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_234 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_19 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_235 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_20 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_236 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_21 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_237 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_22 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_238 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_23 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_239 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
    end
    wb_forward_valid_0 <= mem_forward_valid_0;	// lsu.scala:1064:36, :1189:53
    if (fired_load_incoming_REG)	// lsu.scala:894:51
      wb_forward_ldq_idx_0 <= mem_incoming_uop_0_ldq_idx;	// lsu.scala:908:37, :1065:36
    else if (fired_load_wakeup_REG)	// lsu.scala:904:51
      wb_forward_ldq_idx_0 <= lcam_ldq_idx_REG;	// lsu.scala:1037:58, :1065:36
    else if (fired_load_retry_REG)	// lsu.scala:901:51
      wb_forward_ldq_idx_0 <= lcam_ldq_idx_REG_1;	// lsu.scala:1038:58, :1065:36
    else	// lsu.scala:901:51
      wb_forward_ldq_idx_0 <= 5'h0;	// lsu.scala:1065:36
    if (_lcam_addr_T_1)	// lsu.scala:1025:86
      wb_forward_ld_addr_0 <= _GEN_324;	// lsu.scala:1025:37, :1066:36
    else if (fired_release_0)	// lsu.scala:900:37
      wb_forward_ld_addr_0 <= _GEN_323;	// lsu.scala:1027:41, :1066:36
    else	// lsu.scala:900:37
      wb_forward_ld_addr_0 <= mem_paddr_0;	// lsu.scala:927:41, :1066:36
    wb_forward_stq_idx_0 <= _forwarding_age_logic_0_io_forwarding_idx;	// lsu.scala:1067:36, :1178:57
    older_nacked_REG <= nacking_loads_0;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_1 <= nacking_loads_1;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_1 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_2 <= nacking_loads_2;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_2 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_3 <= nacking_loads_3;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_3 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_4 <= nacking_loads_4;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_4 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_5 <= nacking_loads_5;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_5 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_6 <= nacking_loads_6;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_6 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_7 <= nacking_loads_7;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_7 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_8 <= nacking_loads_8;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_8 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_9 <= nacking_loads_9;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_9 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_10 <= nacking_loads_10;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_10 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_11 <= nacking_loads_11;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_11 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_12 <= nacking_loads_12;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_12 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_13 <= nacking_loads_13;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_13 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_14 <= nacking_loads_14;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_14 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_15 <= nacking_loads_15;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_15 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_16 <= nacking_loads_16;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_16 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_17 <= nacking_loads_17;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_17 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_18 <= nacking_loads_18;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_18 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_19 <= nacking_loads_19;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_19 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_20 <= nacking_loads_20;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_20 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_21 <= nacking_loads_21;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_21 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_22 <= nacking_loads_22;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_22 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_23 <= nacking_loads_23;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_23 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    io_dmem_s1_kill_0_REG_24 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_25 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_26 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_27 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_28 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_29 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_30 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_31 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_32 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_33 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_34 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_35 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_36 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_37 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_38 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_39 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_40 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_41 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_42 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_43 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_44 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_45 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_46 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_47 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_48 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_49 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_50 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_51 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_52 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_53 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_54 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_55 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_56 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_57 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_58 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_59 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_60 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_61 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_62 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_63 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_64 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_65 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_66 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_67 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_68 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_69 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_70 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_71 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_72 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_73 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_74 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_75 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_76 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_77 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_78 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_79 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_80 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_81 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_82 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_83 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_84 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_85 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_86 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_87 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_88 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_89 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_90 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_91 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_92 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_93 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_94 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_95 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    REG_1 <= io_core_exception;	// lsu.scala:1189:64
    REG_2 <=
      (ldst_addr_matches_0_0 | ldst_addr_matches_0_1 | ldst_addr_matches_0_2
       | ldst_addr_matches_0_3 | ldst_addr_matches_0_4 | ldst_addr_matches_0_5
       | ldst_addr_matches_0_6 | ldst_addr_matches_0_7 | ldst_addr_matches_0_8
       | ldst_addr_matches_0_9 | ldst_addr_matches_0_10 | ldst_addr_matches_0_11
       | ldst_addr_matches_0_12 | ldst_addr_matches_0_13 | ldst_addr_matches_0_14
       | ldst_addr_matches_0_15 | ldst_addr_matches_0_16 | ldst_addr_matches_0_17
       | ldst_addr_matches_0_18 | ldst_addr_matches_0_19 | ldst_addr_matches_0_20
       | ldst_addr_matches_0_21 | ldst_addr_matches_0_22 | ldst_addr_matches_0_23)
      & ~mem_forward_valid_0;	// lsu.scala:1148:72, :1150:9, :1189:53, :1199:{18,48,53,56}
    if (will_fire_store_commit_0 | ~can_fire_store_commit_0)	// lsu.scala:493:79, :535:65, :1205:{37,40}
      store_blocked_counter <= 4'h0;	// lsu.scala:1204:36
    else if (can_fire_store_commit_0 & ~will_fire_store_commit_0) begin	// lsu.scala:493:79, :535:65, :584:6, :1207:43
      if (&store_blocked_counter)	// lsu.scala:1204:36, :1208:58
        store_blocked_counter <= store_blocked_counter + 4'h1;	// lsu.scala:305:44, :1204:36, :1208:90
      else	// lsu.scala:1208:58
        store_blocked_counter <= 4'hF;	// lsu.scala:1204:36, util.scala:351:72
    end
    r_xcpt_uop_br_mask <= xcpt_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:1236:25, :1243:21, util.scala:85:{25,27}
    if (use_mem_xcpt) begin	// lsu.scala:1241:115
      r_xcpt_uop_rob_idx <= mem_xcpt_uops_0_rob_idx;	// lsu.scala:671:32, :1236:25
      r_xcpt_cause <= {1'h0, mem_xcpt_causes_0};	// lsu.scala:249:20, :672:32, :708:86, :1236:25, :1250:28
    end
    else begin	// lsu.scala:1241:115
      r_xcpt_uop_rob_idx <= _GEN_148[_ld_xcpt_uop_T_3];	// lsu.scala:465:79, :1236:25, :1239:30, util.scala:363:52
      r_xcpt_cause <= 5'h10;	// lsu.scala:305:44, :1236:25
    end
    r_xcpt_badvaddr <= mem_xcpt_vaddrs_0;	// lsu.scala:679:32, :1236:25
    io_core_ld_miss_REG <= _io_core_spec_ld_wakeup_0_valid_output;	// lsu.scala:1260:69, :1380:37
    spec_ld_succeed_REG <= _io_core_spec_ld_wakeup_0_valid_output;	// lsu.scala:1260:69, :1382:13
    spec_ld_succeed_REG_1 <= mem_incoming_uop_0_ldq_idx;	// lsu.scala:908:37, :1384:56
    if (reset) begin
      hella_state <= 3'h0;	// lsu.scala:242:38
      live_store_mask <= 24'h0;	// lsu.scala:259:32
      clr_bsy_valid_0 <= 1'h0;	// lsu.scala:249:20, :708:86, :930:32
      stdf_clr_bsy_valid <= 1'h0;	// lsu.scala:249:20, :708:86, :983:37
      r_xcpt_valid <= 1'h0;	// lsu.scala:249:20, :708:86, :1235:29
    end
    else begin
      automatic logic [31:0] _GEN_2474 = 32'h1 << _GEN_107;	// lsu.scala:260:71, :336:72, :338:21
      if (|hella_state) begin	// lsu.scala:242:38, :593:24
        automatic logic            _GEN_2475;	// lsu.scala:1540:50
        automatic logic [2:0]      _GEN_2476;	// lsu.scala:242:38, :1582:40, :1584:69, :1585:21
        automatic logic [7:0][2:0] _GEN_2477;	// lsu.scala:803:26, :820:26, :1288:28, :1533:38, :1539:34, :1550:{28,43}, :1552:17, :1553:{28,38}, :1555:63, :1560:40, :1562:69, :1576:42, :1579:76, :1582:40
        _GEN_2475 = will_fire_hella_incoming_0 & dmem_req_fire_0;	// lsu.scala:535:65, :752:55, :1540:50
        _GEN_2476 = _GEN_760 & _GEN_852 ? 3'h0 : hella_state;	// lsu.scala:242:38, :1288:54, :1562:35, :1582:40, :1584:69, :1585:21
        _GEN_2477 =
          {{_GEN_2476},
           {_GEN_2476},
           {will_fire_hella_wakeup_0 & dmem_req_fire_0 ? 3'h4 : hella_state},
           {_GEN_852 ? 3'h0 : _GEN_758 ? 3'h5 : hella_state},
           {3'h0},
           {{1'h1,
             |{hella_xcpt_ma_ld,
               hella_xcpt_ma_st,
               hella_xcpt_pf_ld,
               hella_xcpt_pf_st,
               hella_xcpt_ae_ld,
               hella_xcpt_ae_st},
             1'h0}},
           {io_hellacache_s1_kill ? (_GEN_2475 ? 3'h6 : 3'h0) : {2'h1, ~_GEN_2475}},
           {_GEN_2476}};	// lsu.scala:242:38, :246:34, :249:20, :535:65, :708:86, :752:55, :803:26, :820:26, :1287:7, :1288:28, :1312:58, :1533:38, :1539:34, :1540:{50,80}, :1541:21, :1543:21, :1545:85, :1546:19, :1548:19, :1550:{28,43}, :1552:17, :1553:{28,38}, :1555:{47,54,63}, :1556:19, :1558:19, :1560:40, :1562:{35,69}, :1563:21, :1572:76, :1573:21, :1576:42, :1579:{46,76}, :1580:19, :1582:40, :1584:69, :1585:21, util.scala:351:72
        hella_state <= _GEN_2477[hella_state];	// lsu.scala:242:38, :803:26, :820:26, :1288:28, :1533:38, :1539:34, :1550:{28,43}, :1552:17, :1553:{28,38}, :1555:63, :1560:40, :1562:69, :1576:42, :1579:76, :1582:40
      end
      else if (_GEN_2421)	// Decoupled.scala:40:37
        hella_state <= 3'h1;	// lsu.scala:242:38, :803:26
      live_store_mask <=
        ({24{dis_st_val_2}} & _GEN_2474[23:0] | _GEN_1050)
        & ~{stq_23_valid & (|_GEN_825),
            stq_22_valid & (|_GEN_824),
            stq_21_valid & (|_GEN_823),
            stq_20_valid & (|_GEN_822),
            stq_19_valid & (|_GEN_821),
            stq_18_valid & (|_GEN_820),
            stq_17_valid & (|_GEN_819),
            stq_16_valid & (|_GEN_818),
            stq_15_valid & (|_GEN_817),
            stq_14_valid & (|_GEN_816),
            stq_13_valid & (|_GEN_815),
            stq_12_valid & (|_GEN_814),
            stq_11_valid & (|_GEN_813),
            stq_10_valid & (|_GEN_812),
            stq_9_valid & (|_GEN_811),
            stq_8_valid & (|_GEN_810),
            stq_7_valid & (|_GEN_809),
            stq_6_valid & (|_GEN_808),
            stq_5_valid & (|_GEN_807),
            stq_4_valid & (|_GEN_806),
            stq_3_valid & (|_GEN_805),
            stq_2_valid & (|_GEN_804),
            stq_1_valid & (|_GEN_803),
            stq_0_valid & (|_GEN_802)}
        & ~{_GEN_2424 & ~reset & _GEN_2472,
            _GEN_2424 & ~reset & _GEN_2470,
            _GEN_2424 & ~reset & _GEN_2468,
            _GEN_2424 & ~reset & _GEN_2466,
            _GEN_2424 & ~reset & _GEN_2464,
            _GEN_2424 & ~reset & _GEN_2462,
            _GEN_2424 & ~reset & _GEN_2460,
            _GEN_2424 & ~reset & _GEN_2458,
            _GEN_2424 & ~reset & _GEN_2456,
            _GEN_2424 & ~reset & _GEN_2454,
            _GEN_2424 & ~reset & _GEN_2452,
            _GEN_2424 & ~reset & _GEN_2450,
            _GEN_2424 & ~reset & _GEN_2448,
            _GEN_2424 & ~reset & _GEN_2446,
            _GEN_2424 & ~reset & _GEN_2444,
            _GEN_2424 & ~reset & _GEN_2442,
            _GEN_2424 & ~reset & _GEN_2440,
            _GEN_2424 & ~reset & _GEN_2438,
            _GEN_2424 & ~reset & _GEN_2436,
            _GEN_2424 & ~reset & _GEN_2434,
            _GEN_2424 & ~reset & _GEN_2432,
            _GEN_2424 & ~reset & _GEN_2430,
            _GEN_2424 & ~reset & _GEN_2428,
            _GEN_2424 & ~reset & _GEN_2426};	// lsu.scala:211:16, :259:32, :302:85, :336:{31,72}, :1401:25, :1404:5, :1408:7, :1596:22, :1597:3, :1602:5, :1622:38, :1623:9, :1647:{21,40,48}, :1648:{21,42}, util.scala:118:{51,59}
      if (fired_stad_incoming_REG)	// lsu.scala:895:51
        clr_bsy_valid_0 <=
          mem_stq_incoming_e_0_valid & ~mem_tlb_miss_0
          & ~mem_stq_incoming_e_0_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_incoming_e_0_bits_uop_br_mask) == 16'h0;	// lsu.scala:910:37, :925:41, :930:32, :942:29, :943:{29,68}, util.scala:118:{51,59}
      else if (fired_sta_incoming_REG)	// lsu.scala:896:51
        clr_bsy_valid_0 <=
          mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_data_valid
          & ~mem_tlb_miss_0 & ~mem_stq_incoming_e_0_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_incoming_e_0_bits_uop_br_mask) == 16'h0;	// lsu.scala:910:37, :925:41, :930:32, :950:29, :951:{29,69}, util.scala:118:{51,59}
      else if (fired_std_incoming_REG)	// lsu.scala:897:51
        clr_bsy_valid_0 <=
          mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_addr_valid
          & ~mem_stq_incoming_e_0_bits_addr_is_virtual
          & ~mem_stq_incoming_e_0_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_incoming_e_0_bits_uop_br_mask) == 16'h0;	// lsu.scala:910:37, :930:32, :958:29, :959:{29,74}, util.scala:118:{51,59}
      else	// lsu.scala:897:51
        clr_bsy_valid_0 <=
          fired_sfence_0 | fired_sta_retry_REG & mem_stq_retry_e_valid
          & mem_stq_retry_e_bits_data_valid & ~mem_tlb_miss_0
          & ~mem_stq_retry_e_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_retry_e_bits_uop_br_mask) == 16'h0;	// lsu.scala:899:37, :902:51, :913:37, :925:41, :930:32, :935:25, :963:35, :964:27, :967:38, :968:27, :970:29, :971:29, util.scala:118:{51,59}
      stdf_clr_bsy_valid <=
        fired_stdf_incoming & _GEN_2[mem_stdf_uop_stq_idx] & _GEN_87[mem_stdf_uop_stq_idx]
        & ~_GEN_90[mem_stdf_uop_stq_idx] & ~_GEN_61[mem_stdf_uop_stq_idx]
        & (io_core_brupdate_b1_mispredict_mask & mem_stdf_uop_br_mask) == 16'h0;	// lsu.scala:224:42, :898:37, :922:37, :983:37, :986:24, :989:30, :991:{26,62}, :993:29, :994:29, util.scala:118:{51,59}
      r_xcpt_valid <=
        (ld_xcpt_valid | mem_xcpt_valids_0) & ~io_core_exception
        & (io_core_brupdate_b1_mispredict_mask & xcpt_uop_br_mask) == 16'h0;	// lsu.scala:667:32, :669:22, :1235:29, :1238:44, :1243:21, :1245:34, :1246:39, util.scala:118:{51,59}
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:1022];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [9:0] i = 10'h0; i < 10'h3FF; i += 10'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        ldq_0_valid = _RANDOM[10'h0][0];	// lsu.scala:210:16
        ldq_0_bits_uop_uopc = _RANDOM[10'h0][7:1];	// lsu.scala:210:16
        ldq_0_bits_uop_inst = {_RANDOM[10'h0][31:8], _RANDOM[10'h1][7:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_debug_inst = {_RANDOM[10'h1][31:8], _RANDOM[10'h2][7:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_is_rvc = _RANDOM[10'h2][8];	// lsu.scala:210:16
        ldq_0_bits_uop_debug_pc = {_RANDOM[10'h2][31:9], _RANDOM[10'h3][16:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_iq_type = _RANDOM[10'h3][19:17];	// lsu.scala:210:16
        ldq_0_bits_uop_fu_code = _RANDOM[10'h3][29:20];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_br_type = {_RANDOM[10'h3][31:30], _RANDOM[10'h4][1:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_op1_sel = _RANDOM[10'h4][3:2];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_op2_sel = _RANDOM[10'h4][6:4];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_imm_sel = _RANDOM[10'h4][9:7];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_op_fcn = _RANDOM[10'h4][13:10];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_fcn_dw = _RANDOM[10'h4][14];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_csr_cmd = _RANDOM[10'h4][17:15];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_is_load = _RANDOM[10'h4][18];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_is_sta = _RANDOM[10'h4][19];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_is_std = _RANDOM[10'h4][20];	// lsu.scala:210:16
        ldq_0_bits_uop_iw_state = _RANDOM[10'h4][22:21];	// lsu.scala:210:16
        ldq_0_bits_uop_iw_p1_poisoned = _RANDOM[10'h4][23];	// lsu.scala:210:16
        ldq_0_bits_uop_iw_p2_poisoned = _RANDOM[10'h4][24];	// lsu.scala:210:16
        ldq_0_bits_uop_is_br = _RANDOM[10'h4][25];	// lsu.scala:210:16
        ldq_0_bits_uop_is_jalr = _RANDOM[10'h4][26];	// lsu.scala:210:16
        ldq_0_bits_uop_is_jal = _RANDOM[10'h4][27];	// lsu.scala:210:16
        ldq_0_bits_uop_is_sfb = _RANDOM[10'h4][28];	// lsu.scala:210:16
        ldq_0_bits_uop_br_mask = {_RANDOM[10'h4][31:29], _RANDOM[10'h5][12:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_br_tag = _RANDOM[10'h5][16:13];	// lsu.scala:210:16
        ldq_0_bits_uop_ftq_idx = _RANDOM[10'h5][21:17];	// lsu.scala:210:16
        ldq_0_bits_uop_edge_inst = _RANDOM[10'h5][22];	// lsu.scala:210:16
        ldq_0_bits_uop_pc_lob = _RANDOM[10'h5][28:23];	// lsu.scala:210:16
        ldq_0_bits_uop_taken = _RANDOM[10'h5][29];	// lsu.scala:210:16
        ldq_0_bits_uop_imm_packed = {_RANDOM[10'h5][31:30], _RANDOM[10'h6][17:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_csr_addr = _RANDOM[10'h6][29:18];	// lsu.scala:210:16
        ldq_0_bits_uop_rob_idx = {_RANDOM[10'h6][31:30], _RANDOM[10'h7][4:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_ldq_idx = _RANDOM[10'h7][9:5];	// lsu.scala:210:16
        ldq_0_bits_uop_stq_idx = _RANDOM[10'h7][14:10];	// lsu.scala:210:16
        ldq_0_bits_uop_rxq_idx = _RANDOM[10'h7][16:15];	// lsu.scala:210:16
        ldq_0_bits_uop_pdst = _RANDOM[10'h7][23:17];	// lsu.scala:210:16
        ldq_0_bits_uop_prs1 = _RANDOM[10'h7][30:24];	// lsu.scala:210:16
        ldq_0_bits_uop_prs2 = {_RANDOM[10'h7][31], _RANDOM[10'h8][5:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_prs3 = _RANDOM[10'h8][12:6];	// lsu.scala:210:16
        ldq_0_bits_uop_ppred = _RANDOM[10'h8][17:13];	// lsu.scala:210:16
        ldq_0_bits_uop_prs1_busy = _RANDOM[10'h8][18];	// lsu.scala:210:16
        ldq_0_bits_uop_prs2_busy = _RANDOM[10'h8][19];	// lsu.scala:210:16
        ldq_0_bits_uop_prs3_busy = _RANDOM[10'h8][20];	// lsu.scala:210:16
        ldq_0_bits_uop_ppred_busy = _RANDOM[10'h8][21];	// lsu.scala:210:16
        ldq_0_bits_uop_stale_pdst = _RANDOM[10'h8][28:22];	// lsu.scala:210:16
        ldq_0_bits_uop_exception = _RANDOM[10'h8][29];	// lsu.scala:210:16
        ldq_0_bits_uop_exc_cause =
          {_RANDOM[10'h8][31:30], _RANDOM[10'h9], _RANDOM[10'hA][29:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_bypassable = _RANDOM[10'hA][30];	// lsu.scala:210:16
        ldq_0_bits_uop_mem_cmd = {_RANDOM[10'hA][31], _RANDOM[10'hB][3:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_mem_size = _RANDOM[10'hB][5:4];	// lsu.scala:210:16
        ldq_0_bits_uop_mem_signed = _RANDOM[10'hB][6];	// lsu.scala:210:16
        ldq_0_bits_uop_is_fence = _RANDOM[10'hB][7];	// lsu.scala:210:16
        ldq_0_bits_uop_is_fencei = _RANDOM[10'hB][8];	// lsu.scala:210:16
        ldq_0_bits_uop_is_amo = _RANDOM[10'hB][9];	// lsu.scala:210:16
        ldq_0_bits_uop_uses_ldq = _RANDOM[10'hB][10];	// lsu.scala:210:16
        ldq_0_bits_uop_uses_stq = _RANDOM[10'hB][11];	// lsu.scala:210:16
        ldq_0_bits_uop_is_sys_pc2epc = _RANDOM[10'hB][12];	// lsu.scala:210:16
        ldq_0_bits_uop_is_unique = _RANDOM[10'hB][13];	// lsu.scala:210:16
        ldq_0_bits_uop_flush_on_commit = _RANDOM[10'hB][14];	// lsu.scala:210:16
        ldq_0_bits_uop_ldst_is_rs1 = _RANDOM[10'hB][15];	// lsu.scala:210:16
        ldq_0_bits_uop_ldst = _RANDOM[10'hB][21:16];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs1 = _RANDOM[10'hB][27:22];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs2 = {_RANDOM[10'hB][31:28], _RANDOM[10'hC][1:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_lrs3 = _RANDOM[10'hC][7:2];	// lsu.scala:210:16
        ldq_0_bits_uop_ldst_val = _RANDOM[10'hC][8];	// lsu.scala:210:16
        ldq_0_bits_uop_dst_rtype = _RANDOM[10'hC][10:9];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs1_rtype = _RANDOM[10'hC][12:11];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs2_rtype = _RANDOM[10'hC][14:13];	// lsu.scala:210:16
        ldq_0_bits_uop_frs3_en = _RANDOM[10'hC][15];	// lsu.scala:210:16
        ldq_0_bits_uop_fp_val = _RANDOM[10'hC][16];	// lsu.scala:210:16
        ldq_0_bits_uop_fp_single = _RANDOM[10'hC][17];	// lsu.scala:210:16
        ldq_0_bits_uop_xcpt_pf_if = _RANDOM[10'hC][18];	// lsu.scala:210:16
        ldq_0_bits_uop_xcpt_ae_if = _RANDOM[10'hC][19];	// lsu.scala:210:16
        ldq_0_bits_uop_xcpt_ma_if = _RANDOM[10'hC][20];	// lsu.scala:210:16
        ldq_0_bits_uop_bp_debug_if = _RANDOM[10'hC][21];	// lsu.scala:210:16
        ldq_0_bits_uop_bp_xcpt_if = _RANDOM[10'hC][22];	// lsu.scala:210:16
        ldq_0_bits_uop_debug_fsrc = _RANDOM[10'hC][24:23];	// lsu.scala:210:16
        ldq_0_bits_uop_debug_tsrc = _RANDOM[10'hC][26:25];	// lsu.scala:210:16
        ldq_0_bits_addr_valid = _RANDOM[10'hC][27];	// lsu.scala:210:16
        ldq_0_bits_addr_bits =
          {_RANDOM[10'hC][31:28], _RANDOM[10'hD], _RANDOM[10'hE][3:0]};	// lsu.scala:210:16
        ldq_0_bits_addr_is_virtual = _RANDOM[10'hE][4];	// lsu.scala:210:16
        ldq_0_bits_addr_is_uncacheable = _RANDOM[10'hE][5];	// lsu.scala:210:16
        ldq_0_bits_executed = _RANDOM[10'hE][6];	// lsu.scala:210:16
        ldq_0_bits_succeeded = _RANDOM[10'hE][7];	// lsu.scala:210:16
        ldq_0_bits_order_fail = _RANDOM[10'hE][8];	// lsu.scala:210:16
        ldq_0_bits_observed = _RANDOM[10'hE][9];	// lsu.scala:210:16
        ldq_0_bits_st_dep_mask = {_RANDOM[10'hE][31:10], _RANDOM[10'hF][1:0]};	// lsu.scala:210:16
        ldq_0_bits_youngest_stq_idx = _RANDOM[10'hF][6:2];	// lsu.scala:210:16
        ldq_0_bits_forward_std_val = _RANDOM[10'hF][7];	// lsu.scala:210:16
        ldq_0_bits_forward_stq_idx = _RANDOM[10'hF][12:8];	// lsu.scala:210:16
        ldq_1_valid = _RANDOM[10'h11][13];	// lsu.scala:210:16
        ldq_1_bits_uop_uopc = _RANDOM[10'h11][20:14];	// lsu.scala:210:16
        ldq_1_bits_uop_inst = {_RANDOM[10'h11][31:21], _RANDOM[10'h12][20:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_debug_inst = {_RANDOM[10'h12][31:21], _RANDOM[10'h13][20:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_is_rvc = _RANDOM[10'h13][21];	// lsu.scala:210:16
        ldq_1_bits_uop_debug_pc = {_RANDOM[10'h13][31:22], _RANDOM[10'h14][29:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_iq_type = {_RANDOM[10'h14][31:30], _RANDOM[10'h15][0]};	// lsu.scala:210:16
        ldq_1_bits_uop_fu_code = _RANDOM[10'h15][10:1];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_br_type = _RANDOM[10'h15][14:11];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_op1_sel = _RANDOM[10'h15][16:15];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_op2_sel = _RANDOM[10'h15][19:17];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_imm_sel = _RANDOM[10'h15][22:20];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_op_fcn = _RANDOM[10'h15][26:23];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_fcn_dw = _RANDOM[10'h15][27];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_csr_cmd = _RANDOM[10'h15][30:28];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_is_load = _RANDOM[10'h15][31];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_is_sta = _RANDOM[10'h16][0];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_is_std = _RANDOM[10'h16][1];	// lsu.scala:210:16
        ldq_1_bits_uop_iw_state = _RANDOM[10'h16][3:2];	// lsu.scala:210:16
        ldq_1_bits_uop_iw_p1_poisoned = _RANDOM[10'h16][4];	// lsu.scala:210:16
        ldq_1_bits_uop_iw_p2_poisoned = _RANDOM[10'h16][5];	// lsu.scala:210:16
        ldq_1_bits_uop_is_br = _RANDOM[10'h16][6];	// lsu.scala:210:16
        ldq_1_bits_uop_is_jalr = _RANDOM[10'h16][7];	// lsu.scala:210:16
        ldq_1_bits_uop_is_jal = _RANDOM[10'h16][8];	// lsu.scala:210:16
        ldq_1_bits_uop_is_sfb = _RANDOM[10'h16][9];	// lsu.scala:210:16
        ldq_1_bits_uop_br_mask = _RANDOM[10'h16][25:10];	// lsu.scala:210:16
        ldq_1_bits_uop_br_tag = _RANDOM[10'h16][29:26];	// lsu.scala:210:16
        ldq_1_bits_uop_ftq_idx = {_RANDOM[10'h16][31:30], _RANDOM[10'h17][2:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_edge_inst = _RANDOM[10'h17][3];	// lsu.scala:210:16
        ldq_1_bits_uop_pc_lob = _RANDOM[10'h17][9:4];	// lsu.scala:210:16
        ldq_1_bits_uop_taken = _RANDOM[10'h17][10];	// lsu.scala:210:16
        ldq_1_bits_uop_imm_packed = _RANDOM[10'h17][30:11];	// lsu.scala:210:16
        ldq_1_bits_uop_csr_addr = {_RANDOM[10'h17][31], _RANDOM[10'h18][10:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_rob_idx = _RANDOM[10'h18][17:11];	// lsu.scala:210:16
        ldq_1_bits_uop_ldq_idx = _RANDOM[10'h18][22:18];	// lsu.scala:210:16
        ldq_1_bits_uop_stq_idx = _RANDOM[10'h18][27:23];	// lsu.scala:210:16
        ldq_1_bits_uop_rxq_idx = _RANDOM[10'h18][29:28];	// lsu.scala:210:16
        ldq_1_bits_uop_pdst = {_RANDOM[10'h18][31:30], _RANDOM[10'h19][4:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_prs1 = _RANDOM[10'h19][11:5];	// lsu.scala:210:16
        ldq_1_bits_uop_prs2 = _RANDOM[10'h19][18:12];	// lsu.scala:210:16
        ldq_1_bits_uop_prs3 = _RANDOM[10'h19][25:19];	// lsu.scala:210:16
        ldq_1_bits_uop_ppred = _RANDOM[10'h19][30:26];	// lsu.scala:210:16
        ldq_1_bits_uop_prs1_busy = _RANDOM[10'h19][31];	// lsu.scala:210:16
        ldq_1_bits_uop_prs2_busy = _RANDOM[10'h1A][0];	// lsu.scala:210:16
        ldq_1_bits_uop_prs3_busy = _RANDOM[10'h1A][1];	// lsu.scala:210:16
        ldq_1_bits_uop_ppred_busy = _RANDOM[10'h1A][2];	// lsu.scala:210:16
        ldq_1_bits_uop_stale_pdst = _RANDOM[10'h1A][9:3];	// lsu.scala:210:16
        ldq_1_bits_uop_exception = _RANDOM[10'h1A][10];	// lsu.scala:210:16
        ldq_1_bits_uop_exc_cause =
          {_RANDOM[10'h1A][31:11], _RANDOM[10'h1B], _RANDOM[10'h1C][10:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_bypassable = _RANDOM[10'h1C][11];	// lsu.scala:210:16
        ldq_1_bits_uop_mem_cmd = _RANDOM[10'h1C][16:12];	// lsu.scala:210:16
        ldq_1_bits_uop_mem_size = _RANDOM[10'h1C][18:17];	// lsu.scala:210:16
        ldq_1_bits_uop_mem_signed = _RANDOM[10'h1C][19];	// lsu.scala:210:16
        ldq_1_bits_uop_is_fence = _RANDOM[10'h1C][20];	// lsu.scala:210:16
        ldq_1_bits_uop_is_fencei = _RANDOM[10'h1C][21];	// lsu.scala:210:16
        ldq_1_bits_uop_is_amo = _RANDOM[10'h1C][22];	// lsu.scala:210:16
        ldq_1_bits_uop_uses_ldq = _RANDOM[10'h1C][23];	// lsu.scala:210:16
        ldq_1_bits_uop_uses_stq = _RANDOM[10'h1C][24];	// lsu.scala:210:16
        ldq_1_bits_uop_is_sys_pc2epc = _RANDOM[10'h1C][25];	// lsu.scala:210:16
        ldq_1_bits_uop_is_unique = _RANDOM[10'h1C][26];	// lsu.scala:210:16
        ldq_1_bits_uop_flush_on_commit = _RANDOM[10'h1C][27];	// lsu.scala:210:16
        ldq_1_bits_uop_ldst_is_rs1 = _RANDOM[10'h1C][28];	// lsu.scala:210:16
        ldq_1_bits_uop_ldst = {_RANDOM[10'h1C][31:29], _RANDOM[10'h1D][2:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_lrs1 = _RANDOM[10'h1D][8:3];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs2 = _RANDOM[10'h1D][14:9];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs3 = _RANDOM[10'h1D][20:15];	// lsu.scala:210:16
        ldq_1_bits_uop_ldst_val = _RANDOM[10'h1D][21];	// lsu.scala:210:16
        ldq_1_bits_uop_dst_rtype = _RANDOM[10'h1D][23:22];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs1_rtype = _RANDOM[10'h1D][25:24];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs2_rtype = _RANDOM[10'h1D][27:26];	// lsu.scala:210:16
        ldq_1_bits_uop_frs3_en = _RANDOM[10'h1D][28];	// lsu.scala:210:16
        ldq_1_bits_uop_fp_val = _RANDOM[10'h1D][29];	// lsu.scala:210:16
        ldq_1_bits_uop_fp_single = _RANDOM[10'h1D][30];	// lsu.scala:210:16
        ldq_1_bits_uop_xcpt_pf_if = _RANDOM[10'h1D][31];	// lsu.scala:210:16
        ldq_1_bits_uop_xcpt_ae_if = _RANDOM[10'h1E][0];	// lsu.scala:210:16
        ldq_1_bits_uop_xcpt_ma_if = _RANDOM[10'h1E][1];	// lsu.scala:210:16
        ldq_1_bits_uop_bp_debug_if = _RANDOM[10'h1E][2];	// lsu.scala:210:16
        ldq_1_bits_uop_bp_xcpt_if = _RANDOM[10'h1E][3];	// lsu.scala:210:16
        ldq_1_bits_uop_debug_fsrc = _RANDOM[10'h1E][5:4];	// lsu.scala:210:16
        ldq_1_bits_uop_debug_tsrc = _RANDOM[10'h1E][7:6];	// lsu.scala:210:16
        ldq_1_bits_addr_valid = _RANDOM[10'h1E][8];	// lsu.scala:210:16
        ldq_1_bits_addr_bits = {_RANDOM[10'h1E][31:9], _RANDOM[10'h1F][16:0]};	// lsu.scala:210:16
        ldq_1_bits_addr_is_virtual = _RANDOM[10'h1F][17];	// lsu.scala:210:16
        ldq_1_bits_addr_is_uncacheable = _RANDOM[10'h1F][18];	// lsu.scala:210:16
        ldq_1_bits_executed = _RANDOM[10'h1F][19];	// lsu.scala:210:16
        ldq_1_bits_succeeded = _RANDOM[10'h1F][20];	// lsu.scala:210:16
        ldq_1_bits_order_fail = _RANDOM[10'h1F][21];	// lsu.scala:210:16
        ldq_1_bits_observed = _RANDOM[10'h1F][22];	// lsu.scala:210:16
        ldq_1_bits_st_dep_mask = {_RANDOM[10'h1F][31:23], _RANDOM[10'h20][14:0]};	// lsu.scala:210:16
        ldq_1_bits_youngest_stq_idx = _RANDOM[10'h20][19:15];	// lsu.scala:210:16
        ldq_1_bits_forward_std_val = _RANDOM[10'h20][20];	// lsu.scala:210:16
        ldq_1_bits_forward_stq_idx = _RANDOM[10'h20][25:21];	// lsu.scala:210:16
        ldq_2_valid = _RANDOM[10'h22][26];	// lsu.scala:210:16
        ldq_2_bits_uop_uopc = {_RANDOM[10'h22][31:27], _RANDOM[10'h23][1:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_inst = {_RANDOM[10'h23][31:2], _RANDOM[10'h24][1:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_debug_inst = {_RANDOM[10'h24][31:2], _RANDOM[10'h25][1:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_is_rvc = _RANDOM[10'h25][2];	// lsu.scala:210:16
        ldq_2_bits_uop_debug_pc = {_RANDOM[10'h25][31:3], _RANDOM[10'h26][10:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_iq_type = _RANDOM[10'h26][13:11];	// lsu.scala:210:16
        ldq_2_bits_uop_fu_code = _RANDOM[10'h26][23:14];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_br_type = _RANDOM[10'h26][27:24];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_op1_sel = _RANDOM[10'h26][29:28];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_op2_sel = {_RANDOM[10'h26][31:30], _RANDOM[10'h27][0]};	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_imm_sel = _RANDOM[10'h27][3:1];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_op_fcn = _RANDOM[10'h27][7:4];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_fcn_dw = _RANDOM[10'h27][8];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_csr_cmd = _RANDOM[10'h27][11:9];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_is_load = _RANDOM[10'h27][12];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_is_sta = _RANDOM[10'h27][13];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_is_std = _RANDOM[10'h27][14];	// lsu.scala:210:16
        ldq_2_bits_uop_iw_state = _RANDOM[10'h27][16:15];	// lsu.scala:210:16
        ldq_2_bits_uop_iw_p1_poisoned = _RANDOM[10'h27][17];	// lsu.scala:210:16
        ldq_2_bits_uop_iw_p2_poisoned = _RANDOM[10'h27][18];	// lsu.scala:210:16
        ldq_2_bits_uop_is_br = _RANDOM[10'h27][19];	// lsu.scala:210:16
        ldq_2_bits_uop_is_jalr = _RANDOM[10'h27][20];	// lsu.scala:210:16
        ldq_2_bits_uop_is_jal = _RANDOM[10'h27][21];	// lsu.scala:210:16
        ldq_2_bits_uop_is_sfb = _RANDOM[10'h27][22];	// lsu.scala:210:16
        ldq_2_bits_uop_br_mask = {_RANDOM[10'h27][31:23], _RANDOM[10'h28][6:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_br_tag = _RANDOM[10'h28][10:7];	// lsu.scala:210:16
        ldq_2_bits_uop_ftq_idx = _RANDOM[10'h28][15:11];	// lsu.scala:210:16
        ldq_2_bits_uop_edge_inst = _RANDOM[10'h28][16];	// lsu.scala:210:16
        ldq_2_bits_uop_pc_lob = _RANDOM[10'h28][22:17];	// lsu.scala:210:16
        ldq_2_bits_uop_taken = _RANDOM[10'h28][23];	// lsu.scala:210:16
        ldq_2_bits_uop_imm_packed = {_RANDOM[10'h28][31:24], _RANDOM[10'h29][11:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_csr_addr = _RANDOM[10'h29][23:12];	// lsu.scala:210:16
        ldq_2_bits_uop_rob_idx = _RANDOM[10'h29][30:24];	// lsu.scala:210:16
        ldq_2_bits_uop_ldq_idx = {_RANDOM[10'h29][31], _RANDOM[10'h2A][3:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_stq_idx = _RANDOM[10'h2A][8:4];	// lsu.scala:210:16
        ldq_2_bits_uop_rxq_idx = _RANDOM[10'h2A][10:9];	// lsu.scala:210:16
        ldq_2_bits_uop_pdst = _RANDOM[10'h2A][17:11];	// lsu.scala:210:16
        ldq_2_bits_uop_prs1 = _RANDOM[10'h2A][24:18];	// lsu.scala:210:16
        ldq_2_bits_uop_prs2 = _RANDOM[10'h2A][31:25];	// lsu.scala:210:16
        ldq_2_bits_uop_prs3 = _RANDOM[10'h2B][6:0];	// lsu.scala:210:16
        ldq_2_bits_uop_ppred = _RANDOM[10'h2B][11:7];	// lsu.scala:210:16
        ldq_2_bits_uop_prs1_busy = _RANDOM[10'h2B][12];	// lsu.scala:210:16
        ldq_2_bits_uop_prs2_busy = _RANDOM[10'h2B][13];	// lsu.scala:210:16
        ldq_2_bits_uop_prs3_busy = _RANDOM[10'h2B][14];	// lsu.scala:210:16
        ldq_2_bits_uop_ppred_busy = _RANDOM[10'h2B][15];	// lsu.scala:210:16
        ldq_2_bits_uop_stale_pdst = _RANDOM[10'h2B][22:16];	// lsu.scala:210:16
        ldq_2_bits_uop_exception = _RANDOM[10'h2B][23];	// lsu.scala:210:16
        ldq_2_bits_uop_exc_cause =
          {_RANDOM[10'h2B][31:24], _RANDOM[10'h2C], _RANDOM[10'h2D][23:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_bypassable = _RANDOM[10'h2D][24];	// lsu.scala:210:16
        ldq_2_bits_uop_mem_cmd = _RANDOM[10'h2D][29:25];	// lsu.scala:210:16
        ldq_2_bits_uop_mem_size = _RANDOM[10'h2D][31:30];	// lsu.scala:210:16
        ldq_2_bits_uop_mem_signed = _RANDOM[10'h2E][0];	// lsu.scala:210:16
        ldq_2_bits_uop_is_fence = _RANDOM[10'h2E][1];	// lsu.scala:210:16
        ldq_2_bits_uop_is_fencei = _RANDOM[10'h2E][2];	// lsu.scala:210:16
        ldq_2_bits_uop_is_amo = _RANDOM[10'h2E][3];	// lsu.scala:210:16
        ldq_2_bits_uop_uses_ldq = _RANDOM[10'h2E][4];	// lsu.scala:210:16
        ldq_2_bits_uop_uses_stq = _RANDOM[10'h2E][5];	// lsu.scala:210:16
        ldq_2_bits_uop_is_sys_pc2epc = _RANDOM[10'h2E][6];	// lsu.scala:210:16
        ldq_2_bits_uop_is_unique = _RANDOM[10'h2E][7];	// lsu.scala:210:16
        ldq_2_bits_uop_flush_on_commit = _RANDOM[10'h2E][8];	// lsu.scala:210:16
        ldq_2_bits_uop_ldst_is_rs1 = _RANDOM[10'h2E][9];	// lsu.scala:210:16
        ldq_2_bits_uop_ldst = _RANDOM[10'h2E][15:10];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs1 = _RANDOM[10'h2E][21:16];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs2 = _RANDOM[10'h2E][27:22];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs3 = {_RANDOM[10'h2E][31:28], _RANDOM[10'h2F][1:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_ldst_val = _RANDOM[10'h2F][2];	// lsu.scala:210:16
        ldq_2_bits_uop_dst_rtype = _RANDOM[10'h2F][4:3];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs1_rtype = _RANDOM[10'h2F][6:5];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs2_rtype = _RANDOM[10'h2F][8:7];	// lsu.scala:210:16
        ldq_2_bits_uop_frs3_en = _RANDOM[10'h2F][9];	// lsu.scala:210:16
        ldq_2_bits_uop_fp_val = _RANDOM[10'h2F][10];	// lsu.scala:210:16
        ldq_2_bits_uop_fp_single = _RANDOM[10'h2F][11];	// lsu.scala:210:16
        ldq_2_bits_uop_xcpt_pf_if = _RANDOM[10'h2F][12];	// lsu.scala:210:16
        ldq_2_bits_uop_xcpt_ae_if = _RANDOM[10'h2F][13];	// lsu.scala:210:16
        ldq_2_bits_uop_xcpt_ma_if = _RANDOM[10'h2F][14];	// lsu.scala:210:16
        ldq_2_bits_uop_bp_debug_if = _RANDOM[10'h2F][15];	// lsu.scala:210:16
        ldq_2_bits_uop_bp_xcpt_if = _RANDOM[10'h2F][16];	// lsu.scala:210:16
        ldq_2_bits_uop_debug_fsrc = _RANDOM[10'h2F][18:17];	// lsu.scala:210:16
        ldq_2_bits_uop_debug_tsrc = _RANDOM[10'h2F][20:19];	// lsu.scala:210:16
        ldq_2_bits_addr_valid = _RANDOM[10'h2F][21];	// lsu.scala:210:16
        ldq_2_bits_addr_bits = {_RANDOM[10'h2F][31:22], _RANDOM[10'h30][29:0]};	// lsu.scala:210:16
        ldq_2_bits_addr_is_virtual = _RANDOM[10'h30][30];	// lsu.scala:210:16
        ldq_2_bits_addr_is_uncacheable = _RANDOM[10'h30][31];	// lsu.scala:210:16
        ldq_2_bits_executed = _RANDOM[10'h31][0];	// lsu.scala:210:16
        ldq_2_bits_succeeded = _RANDOM[10'h31][1];	// lsu.scala:210:16
        ldq_2_bits_order_fail = _RANDOM[10'h31][2];	// lsu.scala:210:16
        ldq_2_bits_observed = _RANDOM[10'h31][3];	// lsu.scala:210:16
        ldq_2_bits_st_dep_mask = _RANDOM[10'h31][27:4];	// lsu.scala:210:16
        ldq_2_bits_youngest_stq_idx = {_RANDOM[10'h31][31:28], _RANDOM[10'h32][0]};	// lsu.scala:210:16
        ldq_2_bits_forward_std_val = _RANDOM[10'h32][1];	// lsu.scala:210:16
        ldq_2_bits_forward_stq_idx = _RANDOM[10'h32][6:2];	// lsu.scala:210:16
        ldq_3_valid = _RANDOM[10'h34][7];	// lsu.scala:210:16
        ldq_3_bits_uop_uopc = _RANDOM[10'h34][14:8];	// lsu.scala:210:16
        ldq_3_bits_uop_inst = {_RANDOM[10'h34][31:15], _RANDOM[10'h35][14:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_debug_inst = {_RANDOM[10'h35][31:15], _RANDOM[10'h36][14:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_is_rvc = _RANDOM[10'h36][15];	// lsu.scala:210:16
        ldq_3_bits_uop_debug_pc = {_RANDOM[10'h36][31:16], _RANDOM[10'h37][23:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_iq_type = _RANDOM[10'h37][26:24];	// lsu.scala:210:16
        ldq_3_bits_uop_fu_code = {_RANDOM[10'h37][31:27], _RANDOM[10'h38][4:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_br_type = _RANDOM[10'h38][8:5];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_op1_sel = _RANDOM[10'h38][10:9];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_op2_sel = _RANDOM[10'h38][13:11];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_imm_sel = _RANDOM[10'h38][16:14];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_op_fcn = _RANDOM[10'h38][20:17];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_fcn_dw = _RANDOM[10'h38][21];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_csr_cmd = _RANDOM[10'h38][24:22];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_is_load = _RANDOM[10'h38][25];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_is_sta = _RANDOM[10'h38][26];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_is_std = _RANDOM[10'h38][27];	// lsu.scala:210:16
        ldq_3_bits_uop_iw_state = _RANDOM[10'h38][29:28];	// lsu.scala:210:16
        ldq_3_bits_uop_iw_p1_poisoned = _RANDOM[10'h38][30];	// lsu.scala:210:16
        ldq_3_bits_uop_iw_p2_poisoned = _RANDOM[10'h38][31];	// lsu.scala:210:16
        ldq_3_bits_uop_is_br = _RANDOM[10'h39][0];	// lsu.scala:210:16
        ldq_3_bits_uop_is_jalr = _RANDOM[10'h39][1];	// lsu.scala:210:16
        ldq_3_bits_uop_is_jal = _RANDOM[10'h39][2];	// lsu.scala:210:16
        ldq_3_bits_uop_is_sfb = _RANDOM[10'h39][3];	// lsu.scala:210:16
        ldq_3_bits_uop_br_mask = _RANDOM[10'h39][19:4];	// lsu.scala:210:16
        ldq_3_bits_uop_br_tag = _RANDOM[10'h39][23:20];	// lsu.scala:210:16
        ldq_3_bits_uop_ftq_idx = _RANDOM[10'h39][28:24];	// lsu.scala:210:16
        ldq_3_bits_uop_edge_inst = _RANDOM[10'h39][29];	// lsu.scala:210:16
        ldq_3_bits_uop_pc_lob = {_RANDOM[10'h39][31:30], _RANDOM[10'h3A][3:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_taken = _RANDOM[10'h3A][4];	// lsu.scala:210:16
        ldq_3_bits_uop_imm_packed = _RANDOM[10'h3A][24:5];	// lsu.scala:210:16
        ldq_3_bits_uop_csr_addr = {_RANDOM[10'h3A][31:25], _RANDOM[10'h3B][4:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_rob_idx = _RANDOM[10'h3B][11:5];	// lsu.scala:210:16
        ldq_3_bits_uop_ldq_idx = _RANDOM[10'h3B][16:12];	// lsu.scala:210:16
        ldq_3_bits_uop_stq_idx = _RANDOM[10'h3B][21:17];	// lsu.scala:210:16
        ldq_3_bits_uop_rxq_idx = _RANDOM[10'h3B][23:22];	// lsu.scala:210:16
        ldq_3_bits_uop_pdst = _RANDOM[10'h3B][30:24];	// lsu.scala:210:16
        ldq_3_bits_uop_prs1 = {_RANDOM[10'h3B][31], _RANDOM[10'h3C][5:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_prs2 = _RANDOM[10'h3C][12:6];	// lsu.scala:210:16
        ldq_3_bits_uop_prs3 = _RANDOM[10'h3C][19:13];	// lsu.scala:210:16
        ldq_3_bits_uop_ppred = _RANDOM[10'h3C][24:20];	// lsu.scala:210:16
        ldq_3_bits_uop_prs1_busy = _RANDOM[10'h3C][25];	// lsu.scala:210:16
        ldq_3_bits_uop_prs2_busy = _RANDOM[10'h3C][26];	// lsu.scala:210:16
        ldq_3_bits_uop_prs3_busy = _RANDOM[10'h3C][27];	// lsu.scala:210:16
        ldq_3_bits_uop_ppred_busy = _RANDOM[10'h3C][28];	// lsu.scala:210:16
        ldq_3_bits_uop_stale_pdst = {_RANDOM[10'h3C][31:29], _RANDOM[10'h3D][3:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_exception = _RANDOM[10'h3D][4];	// lsu.scala:210:16
        ldq_3_bits_uop_exc_cause =
          {_RANDOM[10'h3D][31:5], _RANDOM[10'h3E], _RANDOM[10'h3F][4:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_bypassable = _RANDOM[10'h3F][5];	// lsu.scala:210:16
        ldq_3_bits_uop_mem_cmd = _RANDOM[10'h3F][10:6];	// lsu.scala:210:16
        ldq_3_bits_uop_mem_size = _RANDOM[10'h3F][12:11];	// lsu.scala:210:16
        ldq_3_bits_uop_mem_signed = _RANDOM[10'h3F][13];	// lsu.scala:210:16
        ldq_3_bits_uop_is_fence = _RANDOM[10'h3F][14];	// lsu.scala:210:16
        ldq_3_bits_uop_is_fencei = _RANDOM[10'h3F][15];	// lsu.scala:210:16
        ldq_3_bits_uop_is_amo = _RANDOM[10'h3F][16];	// lsu.scala:210:16
        ldq_3_bits_uop_uses_ldq = _RANDOM[10'h3F][17];	// lsu.scala:210:16
        ldq_3_bits_uop_uses_stq = _RANDOM[10'h3F][18];	// lsu.scala:210:16
        ldq_3_bits_uop_is_sys_pc2epc = _RANDOM[10'h3F][19];	// lsu.scala:210:16
        ldq_3_bits_uop_is_unique = _RANDOM[10'h3F][20];	// lsu.scala:210:16
        ldq_3_bits_uop_flush_on_commit = _RANDOM[10'h3F][21];	// lsu.scala:210:16
        ldq_3_bits_uop_ldst_is_rs1 = _RANDOM[10'h3F][22];	// lsu.scala:210:16
        ldq_3_bits_uop_ldst = _RANDOM[10'h3F][28:23];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs1 = {_RANDOM[10'h3F][31:29], _RANDOM[10'h40][2:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_lrs2 = _RANDOM[10'h40][8:3];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs3 = _RANDOM[10'h40][14:9];	// lsu.scala:210:16
        ldq_3_bits_uop_ldst_val = _RANDOM[10'h40][15];	// lsu.scala:210:16
        ldq_3_bits_uop_dst_rtype = _RANDOM[10'h40][17:16];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs1_rtype = _RANDOM[10'h40][19:18];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs2_rtype = _RANDOM[10'h40][21:20];	// lsu.scala:210:16
        ldq_3_bits_uop_frs3_en = _RANDOM[10'h40][22];	// lsu.scala:210:16
        ldq_3_bits_uop_fp_val = _RANDOM[10'h40][23];	// lsu.scala:210:16
        ldq_3_bits_uop_fp_single = _RANDOM[10'h40][24];	// lsu.scala:210:16
        ldq_3_bits_uop_xcpt_pf_if = _RANDOM[10'h40][25];	// lsu.scala:210:16
        ldq_3_bits_uop_xcpt_ae_if = _RANDOM[10'h40][26];	// lsu.scala:210:16
        ldq_3_bits_uop_xcpt_ma_if = _RANDOM[10'h40][27];	// lsu.scala:210:16
        ldq_3_bits_uop_bp_debug_if = _RANDOM[10'h40][28];	// lsu.scala:210:16
        ldq_3_bits_uop_bp_xcpt_if = _RANDOM[10'h40][29];	// lsu.scala:210:16
        ldq_3_bits_uop_debug_fsrc = _RANDOM[10'h40][31:30];	// lsu.scala:210:16
        ldq_3_bits_uop_debug_tsrc = _RANDOM[10'h41][1:0];	// lsu.scala:210:16
        ldq_3_bits_addr_valid = _RANDOM[10'h41][2];	// lsu.scala:210:16
        ldq_3_bits_addr_bits = {_RANDOM[10'h41][31:3], _RANDOM[10'h42][10:0]};	// lsu.scala:210:16
        ldq_3_bits_addr_is_virtual = _RANDOM[10'h42][11];	// lsu.scala:210:16
        ldq_3_bits_addr_is_uncacheable = _RANDOM[10'h42][12];	// lsu.scala:210:16
        ldq_3_bits_executed = _RANDOM[10'h42][13];	// lsu.scala:210:16
        ldq_3_bits_succeeded = _RANDOM[10'h42][14];	// lsu.scala:210:16
        ldq_3_bits_order_fail = _RANDOM[10'h42][15];	// lsu.scala:210:16
        ldq_3_bits_observed = _RANDOM[10'h42][16];	// lsu.scala:210:16
        ldq_3_bits_st_dep_mask = {_RANDOM[10'h42][31:17], _RANDOM[10'h43][8:0]};	// lsu.scala:210:16
        ldq_3_bits_youngest_stq_idx = _RANDOM[10'h43][13:9];	// lsu.scala:210:16
        ldq_3_bits_forward_std_val = _RANDOM[10'h43][14];	// lsu.scala:210:16
        ldq_3_bits_forward_stq_idx = _RANDOM[10'h43][19:15];	// lsu.scala:210:16
        ldq_4_valid = _RANDOM[10'h45][20];	// lsu.scala:210:16
        ldq_4_bits_uop_uopc = _RANDOM[10'h45][27:21];	// lsu.scala:210:16
        ldq_4_bits_uop_inst = {_RANDOM[10'h45][31:28], _RANDOM[10'h46][27:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_debug_inst = {_RANDOM[10'h46][31:28], _RANDOM[10'h47][27:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_is_rvc = _RANDOM[10'h47][28];	// lsu.scala:210:16
        ldq_4_bits_uop_debug_pc =
          {_RANDOM[10'h47][31:29], _RANDOM[10'h48], _RANDOM[10'h49][4:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_iq_type = _RANDOM[10'h49][7:5];	// lsu.scala:210:16
        ldq_4_bits_uop_fu_code = _RANDOM[10'h49][17:8];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_br_type = _RANDOM[10'h49][21:18];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_op1_sel = _RANDOM[10'h49][23:22];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_op2_sel = _RANDOM[10'h49][26:24];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_imm_sel = _RANDOM[10'h49][29:27];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_op_fcn = {_RANDOM[10'h49][31:30], _RANDOM[10'h4A][1:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_fcn_dw = _RANDOM[10'h4A][2];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_csr_cmd = _RANDOM[10'h4A][5:3];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_is_load = _RANDOM[10'h4A][6];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_is_sta = _RANDOM[10'h4A][7];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_is_std = _RANDOM[10'h4A][8];	// lsu.scala:210:16
        ldq_4_bits_uop_iw_state = _RANDOM[10'h4A][10:9];	// lsu.scala:210:16
        ldq_4_bits_uop_iw_p1_poisoned = _RANDOM[10'h4A][11];	// lsu.scala:210:16
        ldq_4_bits_uop_iw_p2_poisoned = _RANDOM[10'h4A][12];	// lsu.scala:210:16
        ldq_4_bits_uop_is_br = _RANDOM[10'h4A][13];	// lsu.scala:210:16
        ldq_4_bits_uop_is_jalr = _RANDOM[10'h4A][14];	// lsu.scala:210:16
        ldq_4_bits_uop_is_jal = _RANDOM[10'h4A][15];	// lsu.scala:210:16
        ldq_4_bits_uop_is_sfb = _RANDOM[10'h4A][16];	// lsu.scala:210:16
        ldq_4_bits_uop_br_mask = {_RANDOM[10'h4A][31:17], _RANDOM[10'h4B][0]};	// lsu.scala:210:16
        ldq_4_bits_uop_br_tag = _RANDOM[10'h4B][4:1];	// lsu.scala:210:16
        ldq_4_bits_uop_ftq_idx = _RANDOM[10'h4B][9:5];	// lsu.scala:210:16
        ldq_4_bits_uop_edge_inst = _RANDOM[10'h4B][10];	// lsu.scala:210:16
        ldq_4_bits_uop_pc_lob = _RANDOM[10'h4B][16:11];	// lsu.scala:210:16
        ldq_4_bits_uop_taken = _RANDOM[10'h4B][17];	// lsu.scala:210:16
        ldq_4_bits_uop_imm_packed = {_RANDOM[10'h4B][31:18], _RANDOM[10'h4C][5:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_csr_addr = _RANDOM[10'h4C][17:6];	// lsu.scala:210:16
        ldq_4_bits_uop_rob_idx = _RANDOM[10'h4C][24:18];	// lsu.scala:210:16
        ldq_4_bits_uop_ldq_idx = _RANDOM[10'h4C][29:25];	// lsu.scala:210:16
        ldq_4_bits_uop_stq_idx = {_RANDOM[10'h4C][31:30], _RANDOM[10'h4D][2:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_rxq_idx = _RANDOM[10'h4D][4:3];	// lsu.scala:210:16
        ldq_4_bits_uop_pdst = _RANDOM[10'h4D][11:5];	// lsu.scala:210:16
        ldq_4_bits_uop_prs1 = _RANDOM[10'h4D][18:12];	// lsu.scala:210:16
        ldq_4_bits_uop_prs2 = _RANDOM[10'h4D][25:19];	// lsu.scala:210:16
        ldq_4_bits_uop_prs3 = {_RANDOM[10'h4D][31:26], _RANDOM[10'h4E][0]};	// lsu.scala:210:16
        ldq_4_bits_uop_ppred = _RANDOM[10'h4E][5:1];	// lsu.scala:210:16
        ldq_4_bits_uop_prs1_busy = _RANDOM[10'h4E][6];	// lsu.scala:210:16
        ldq_4_bits_uop_prs2_busy = _RANDOM[10'h4E][7];	// lsu.scala:210:16
        ldq_4_bits_uop_prs3_busy = _RANDOM[10'h4E][8];	// lsu.scala:210:16
        ldq_4_bits_uop_ppred_busy = _RANDOM[10'h4E][9];	// lsu.scala:210:16
        ldq_4_bits_uop_stale_pdst = _RANDOM[10'h4E][16:10];	// lsu.scala:210:16
        ldq_4_bits_uop_exception = _RANDOM[10'h4E][17];	// lsu.scala:210:16
        ldq_4_bits_uop_exc_cause =
          {_RANDOM[10'h4E][31:18], _RANDOM[10'h4F], _RANDOM[10'h50][17:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_bypassable = _RANDOM[10'h50][18];	// lsu.scala:210:16
        ldq_4_bits_uop_mem_cmd = _RANDOM[10'h50][23:19];	// lsu.scala:210:16
        ldq_4_bits_uop_mem_size = _RANDOM[10'h50][25:24];	// lsu.scala:210:16
        ldq_4_bits_uop_mem_signed = _RANDOM[10'h50][26];	// lsu.scala:210:16
        ldq_4_bits_uop_is_fence = _RANDOM[10'h50][27];	// lsu.scala:210:16
        ldq_4_bits_uop_is_fencei = _RANDOM[10'h50][28];	// lsu.scala:210:16
        ldq_4_bits_uop_is_amo = _RANDOM[10'h50][29];	// lsu.scala:210:16
        ldq_4_bits_uop_uses_ldq = _RANDOM[10'h50][30];	// lsu.scala:210:16
        ldq_4_bits_uop_uses_stq = _RANDOM[10'h50][31];	// lsu.scala:210:16
        ldq_4_bits_uop_is_sys_pc2epc = _RANDOM[10'h51][0];	// lsu.scala:210:16
        ldq_4_bits_uop_is_unique = _RANDOM[10'h51][1];	// lsu.scala:210:16
        ldq_4_bits_uop_flush_on_commit = _RANDOM[10'h51][2];	// lsu.scala:210:16
        ldq_4_bits_uop_ldst_is_rs1 = _RANDOM[10'h51][3];	// lsu.scala:210:16
        ldq_4_bits_uop_ldst = _RANDOM[10'h51][9:4];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs1 = _RANDOM[10'h51][15:10];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs2 = _RANDOM[10'h51][21:16];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs3 = _RANDOM[10'h51][27:22];	// lsu.scala:210:16
        ldq_4_bits_uop_ldst_val = _RANDOM[10'h51][28];	// lsu.scala:210:16
        ldq_4_bits_uop_dst_rtype = _RANDOM[10'h51][30:29];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs1_rtype = {_RANDOM[10'h51][31], _RANDOM[10'h52][0]};	// lsu.scala:210:16
        ldq_4_bits_uop_lrs2_rtype = _RANDOM[10'h52][2:1];	// lsu.scala:210:16
        ldq_4_bits_uop_frs3_en = _RANDOM[10'h52][3];	// lsu.scala:210:16
        ldq_4_bits_uop_fp_val = _RANDOM[10'h52][4];	// lsu.scala:210:16
        ldq_4_bits_uop_fp_single = _RANDOM[10'h52][5];	// lsu.scala:210:16
        ldq_4_bits_uop_xcpt_pf_if = _RANDOM[10'h52][6];	// lsu.scala:210:16
        ldq_4_bits_uop_xcpt_ae_if = _RANDOM[10'h52][7];	// lsu.scala:210:16
        ldq_4_bits_uop_xcpt_ma_if = _RANDOM[10'h52][8];	// lsu.scala:210:16
        ldq_4_bits_uop_bp_debug_if = _RANDOM[10'h52][9];	// lsu.scala:210:16
        ldq_4_bits_uop_bp_xcpt_if = _RANDOM[10'h52][10];	// lsu.scala:210:16
        ldq_4_bits_uop_debug_fsrc = _RANDOM[10'h52][12:11];	// lsu.scala:210:16
        ldq_4_bits_uop_debug_tsrc = _RANDOM[10'h52][14:13];	// lsu.scala:210:16
        ldq_4_bits_addr_valid = _RANDOM[10'h52][15];	// lsu.scala:210:16
        ldq_4_bits_addr_bits = {_RANDOM[10'h52][31:16], _RANDOM[10'h53][23:0]};	// lsu.scala:210:16
        ldq_4_bits_addr_is_virtual = _RANDOM[10'h53][24];	// lsu.scala:210:16
        ldq_4_bits_addr_is_uncacheable = _RANDOM[10'h53][25];	// lsu.scala:210:16
        ldq_4_bits_executed = _RANDOM[10'h53][26];	// lsu.scala:210:16
        ldq_4_bits_succeeded = _RANDOM[10'h53][27];	// lsu.scala:210:16
        ldq_4_bits_order_fail = _RANDOM[10'h53][28];	// lsu.scala:210:16
        ldq_4_bits_observed = _RANDOM[10'h53][29];	// lsu.scala:210:16
        ldq_4_bits_st_dep_mask = {_RANDOM[10'h53][31:30], _RANDOM[10'h54][21:0]};	// lsu.scala:210:16
        ldq_4_bits_youngest_stq_idx = _RANDOM[10'h54][26:22];	// lsu.scala:210:16
        ldq_4_bits_forward_std_val = _RANDOM[10'h54][27];	// lsu.scala:210:16
        ldq_4_bits_forward_stq_idx = {_RANDOM[10'h54][31:28], _RANDOM[10'h55][0]};	// lsu.scala:210:16
        ldq_5_valid = _RANDOM[10'h57][1];	// lsu.scala:210:16
        ldq_5_bits_uop_uopc = _RANDOM[10'h57][8:2];	// lsu.scala:210:16
        ldq_5_bits_uop_inst = {_RANDOM[10'h57][31:9], _RANDOM[10'h58][8:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_debug_inst = {_RANDOM[10'h58][31:9], _RANDOM[10'h59][8:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_is_rvc = _RANDOM[10'h59][9];	// lsu.scala:210:16
        ldq_5_bits_uop_debug_pc = {_RANDOM[10'h59][31:10], _RANDOM[10'h5A][17:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_iq_type = _RANDOM[10'h5A][20:18];	// lsu.scala:210:16
        ldq_5_bits_uop_fu_code = _RANDOM[10'h5A][30:21];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_br_type = {_RANDOM[10'h5A][31], _RANDOM[10'h5B][2:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_op1_sel = _RANDOM[10'h5B][4:3];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_op2_sel = _RANDOM[10'h5B][7:5];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_imm_sel = _RANDOM[10'h5B][10:8];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_op_fcn = _RANDOM[10'h5B][14:11];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_fcn_dw = _RANDOM[10'h5B][15];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_csr_cmd = _RANDOM[10'h5B][18:16];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_is_load = _RANDOM[10'h5B][19];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_is_sta = _RANDOM[10'h5B][20];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_is_std = _RANDOM[10'h5B][21];	// lsu.scala:210:16
        ldq_5_bits_uop_iw_state = _RANDOM[10'h5B][23:22];	// lsu.scala:210:16
        ldq_5_bits_uop_iw_p1_poisoned = _RANDOM[10'h5B][24];	// lsu.scala:210:16
        ldq_5_bits_uop_iw_p2_poisoned = _RANDOM[10'h5B][25];	// lsu.scala:210:16
        ldq_5_bits_uop_is_br = _RANDOM[10'h5B][26];	// lsu.scala:210:16
        ldq_5_bits_uop_is_jalr = _RANDOM[10'h5B][27];	// lsu.scala:210:16
        ldq_5_bits_uop_is_jal = _RANDOM[10'h5B][28];	// lsu.scala:210:16
        ldq_5_bits_uop_is_sfb = _RANDOM[10'h5B][29];	// lsu.scala:210:16
        ldq_5_bits_uop_br_mask = {_RANDOM[10'h5B][31:30], _RANDOM[10'h5C][13:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_br_tag = _RANDOM[10'h5C][17:14];	// lsu.scala:210:16
        ldq_5_bits_uop_ftq_idx = _RANDOM[10'h5C][22:18];	// lsu.scala:210:16
        ldq_5_bits_uop_edge_inst = _RANDOM[10'h5C][23];	// lsu.scala:210:16
        ldq_5_bits_uop_pc_lob = _RANDOM[10'h5C][29:24];	// lsu.scala:210:16
        ldq_5_bits_uop_taken = _RANDOM[10'h5C][30];	// lsu.scala:210:16
        ldq_5_bits_uop_imm_packed = {_RANDOM[10'h5C][31], _RANDOM[10'h5D][18:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_csr_addr = _RANDOM[10'h5D][30:19];	// lsu.scala:210:16
        ldq_5_bits_uop_rob_idx = {_RANDOM[10'h5D][31], _RANDOM[10'h5E][5:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_ldq_idx = _RANDOM[10'h5E][10:6];	// lsu.scala:210:16
        ldq_5_bits_uop_stq_idx = _RANDOM[10'h5E][15:11];	// lsu.scala:210:16
        ldq_5_bits_uop_rxq_idx = _RANDOM[10'h5E][17:16];	// lsu.scala:210:16
        ldq_5_bits_uop_pdst = _RANDOM[10'h5E][24:18];	// lsu.scala:210:16
        ldq_5_bits_uop_prs1 = _RANDOM[10'h5E][31:25];	// lsu.scala:210:16
        ldq_5_bits_uop_prs2 = _RANDOM[10'h5F][6:0];	// lsu.scala:210:16
        ldq_5_bits_uop_prs3 = _RANDOM[10'h5F][13:7];	// lsu.scala:210:16
        ldq_5_bits_uop_ppred = _RANDOM[10'h5F][18:14];	// lsu.scala:210:16
        ldq_5_bits_uop_prs1_busy = _RANDOM[10'h5F][19];	// lsu.scala:210:16
        ldq_5_bits_uop_prs2_busy = _RANDOM[10'h5F][20];	// lsu.scala:210:16
        ldq_5_bits_uop_prs3_busy = _RANDOM[10'h5F][21];	// lsu.scala:210:16
        ldq_5_bits_uop_ppred_busy = _RANDOM[10'h5F][22];	// lsu.scala:210:16
        ldq_5_bits_uop_stale_pdst = _RANDOM[10'h5F][29:23];	// lsu.scala:210:16
        ldq_5_bits_uop_exception = _RANDOM[10'h5F][30];	// lsu.scala:210:16
        ldq_5_bits_uop_exc_cause =
          {_RANDOM[10'h5F][31], _RANDOM[10'h60], _RANDOM[10'h61][30:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_bypassable = _RANDOM[10'h61][31];	// lsu.scala:210:16
        ldq_5_bits_uop_mem_cmd = _RANDOM[10'h62][4:0];	// lsu.scala:210:16
        ldq_5_bits_uop_mem_size = _RANDOM[10'h62][6:5];	// lsu.scala:210:16
        ldq_5_bits_uop_mem_signed = _RANDOM[10'h62][7];	// lsu.scala:210:16
        ldq_5_bits_uop_is_fence = _RANDOM[10'h62][8];	// lsu.scala:210:16
        ldq_5_bits_uop_is_fencei = _RANDOM[10'h62][9];	// lsu.scala:210:16
        ldq_5_bits_uop_is_amo = _RANDOM[10'h62][10];	// lsu.scala:210:16
        ldq_5_bits_uop_uses_ldq = _RANDOM[10'h62][11];	// lsu.scala:210:16
        ldq_5_bits_uop_uses_stq = _RANDOM[10'h62][12];	// lsu.scala:210:16
        ldq_5_bits_uop_is_sys_pc2epc = _RANDOM[10'h62][13];	// lsu.scala:210:16
        ldq_5_bits_uop_is_unique = _RANDOM[10'h62][14];	// lsu.scala:210:16
        ldq_5_bits_uop_flush_on_commit = _RANDOM[10'h62][15];	// lsu.scala:210:16
        ldq_5_bits_uop_ldst_is_rs1 = _RANDOM[10'h62][16];	// lsu.scala:210:16
        ldq_5_bits_uop_ldst = _RANDOM[10'h62][22:17];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs1 = _RANDOM[10'h62][28:23];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs2 = {_RANDOM[10'h62][31:29], _RANDOM[10'h63][2:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_lrs3 = _RANDOM[10'h63][8:3];	// lsu.scala:210:16
        ldq_5_bits_uop_ldst_val = _RANDOM[10'h63][9];	// lsu.scala:210:16
        ldq_5_bits_uop_dst_rtype = _RANDOM[10'h63][11:10];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs1_rtype = _RANDOM[10'h63][13:12];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs2_rtype = _RANDOM[10'h63][15:14];	// lsu.scala:210:16
        ldq_5_bits_uop_frs3_en = _RANDOM[10'h63][16];	// lsu.scala:210:16
        ldq_5_bits_uop_fp_val = _RANDOM[10'h63][17];	// lsu.scala:210:16
        ldq_5_bits_uop_fp_single = _RANDOM[10'h63][18];	// lsu.scala:210:16
        ldq_5_bits_uop_xcpt_pf_if = _RANDOM[10'h63][19];	// lsu.scala:210:16
        ldq_5_bits_uop_xcpt_ae_if = _RANDOM[10'h63][20];	// lsu.scala:210:16
        ldq_5_bits_uop_xcpt_ma_if = _RANDOM[10'h63][21];	// lsu.scala:210:16
        ldq_5_bits_uop_bp_debug_if = _RANDOM[10'h63][22];	// lsu.scala:210:16
        ldq_5_bits_uop_bp_xcpt_if = _RANDOM[10'h63][23];	// lsu.scala:210:16
        ldq_5_bits_uop_debug_fsrc = _RANDOM[10'h63][25:24];	// lsu.scala:210:16
        ldq_5_bits_uop_debug_tsrc = _RANDOM[10'h63][27:26];	// lsu.scala:210:16
        ldq_5_bits_addr_valid = _RANDOM[10'h63][28];	// lsu.scala:210:16
        ldq_5_bits_addr_bits =
          {_RANDOM[10'h63][31:29], _RANDOM[10'h64], _RANDOM[10'h65][4:0]};	// lsu.scala:210:16
        ldq_5_bits_addr_is_virtual = _RANDOM[10'h65][5];	// lsu.scala:210:16
        ldq_5_bits_addr_is_uncacheable = _RANDOM[10'h65][6];	// lsu.scala:210:16
        ldq_5_bits_executed = _RANDOM[10'h65][7];	// lsu.scala:210:16
        ldq_5_bits_succeeded = _RANDOM[10'h65][8];	// lsu.scala:210:16
        ldq_5_bits_order_fail = _RANDOM[10'h65][9];	// lsu.scala:210:16
        ldq_5_bits_observed = _RANDOM[10'h65][10];	// lsu.scala:210:16
        ldq_5_bits_st_dep_mask = {_RANDOM[10'h65][31:11], _RANDOM[10'h66][2:0]};	// lsu.scala:210:16
        ldq_5_bits_youngest_stq_idx = _RANDOM[10'h66][7:3];	// lsu.scala:210:16
        ldq_5_bits_forward_std_val = _RANDOM[10'h66][8];	// lsu.scala:210:16
        ldq_5_bits_forward_stq_idx = _RANDOM[10'h66][13:9];	// lsu.scala:210:16
        ldq_6_valid = _RANDOM[10'h68][14];	// lsu.scala:210:16
        ldq_6_bits_uop_uopc = _RANDOM[10'h68][21:15];	// lsu.scala:210:16
        ldq_6_bits_uop_inst = {_RANDOM[10'h68][31:22], _RANDOM[10'h69][21:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_debug_inst = {_RANDOM[10'h69][31:22], _RANDOM[10'h6A][21:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_is_rvc = _RANDOM[10'h6A][22];	// lsu.scala:210:16
        ldq_6_bits_uop_debug_pc = {_RANDOM[10'h6A][31:23], _RANDOM[10'h6B][30:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_iq_type = {_RANDOM[10'h6B][31], _RANDOM[10'h6C][1:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_fu_code = _RANDOM[10'h6C][11:2];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_br_type = _RANDOM[10'h6C][15:12];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_op1_sel = _RANDOM[10'h6C][17:16];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_op2_sel = _RANDOM[10'h6C][20:18];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_imm_sel = _RANDOM[10'h6C][23:21];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_op_fcn = _RANDOM[10'h6C][27:24];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_fcn_dw = _RANDOM[10'h6C][28];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_csr_cmd = _RANDOM[10'h6C][31:29];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_is_load = _RANDOM[10'h6D][0];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_is_sta = _RANDOM[10'h6D][1];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_is_std = _RANDOM[10'h6D][2];	// lsu.scala:210:16
        ldq_6_bits_uop_iw_state = _RANDOM[10'h6D][4:3];	// lsu.scala:210:16
        ldq_6_bits_uop_iw_p1_poisoned = _RANDOM[10'h6D][5];	// lsu.scala:210:16
        ldq_6_bits_uop_iw_p2_poisoned = _RANDOM[10'h6D][6];	// lsu.scala:210:16
        ldq_6_bits_uop_is_br = _RANDOM[10'h6D][7];	// lsu.scala:210:16
        ldq_6_bits_uop_is_jalr = _RANDOM[10'h6D][8];	// lsu.scala:210:16
        ldq_6_bits_uop_is_jal = _RANDOM[10'h6D][9];	// lsu.scala:210:16
        ldq_6_bits_uop_is_sfb = _RANDOM[10'h6D][10];	// lsu.scala:210:16
        ldq_6_bits_uop_br_mask = _RANDOM[10'h6D][26:11];	// lsu.scala:210:16
        ldq_6_bits_uop_br_tag = _RANDOM[10'h6D][30:27];	// lsu.scala:210:16
        ldq_6_bits_uop_ftq_idx = {_RANDOM[10'h6D][31], _RANDOM[10'h6E][3:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_edge_inst = _RANDOM[10'h6E][4];	// lsu.scala:210:16
        ldq_6_bits_uop_pc_lob = _RANDOM[10'h6E][10:5];	// lsu.scala:210:16
        ldq_6_bits_uop_taken = _RANDOM[10'h6E][11];	// lsu.scala:210:16
        ldq_6_bits_uop_imm_packed = _RANDOM[10'h6E][31:12];	// lsu.scala:210:16
        ldq_6_bits_uop_csr_addr = _RANDOM[10'h6F][11:0];	// lsu.scala:210:16
        ldq_6_bits_uop_rob_idx = _RANDOM[10'h6F][18:12];	// lsu.scala:210:16
        ldq_6_bits_uop_ldq_idx = _RANDOM[10'h6F][23:19];	// lsu.scala:210:16
        ldq_6_bits_uop_stq_idx = _RANDOM[10'h6F][28:24];	// lsu.scala:210:16
        ldq_6_bits_uop_rxq_idx = _RANDOM[10'h6F][30:29];	// lsu.scala:210:16
        ldq_6_bits_uop_pdst = {_RANDOM[10'h6F][31], _RANDOM[10'h70][5:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_prs1 = _RANDOM[10'h70][12:6];	// lsu.scala:210:16
        ldq_6_bits_uop_prs2 = _RANDOM[10'h70][19:13];	// lsu.scala:210:16
        ldq_6_bits_uop_prs3 = _RANDOM[10'h70][26:20];	// lsu.scala:210:16
        ldq_6_bits_uop_ppred = _RANDOM[10'h70][31:27];	// lsu.scala:210:16
        ldq_6_bits_uop_prs1_busy = _RANDOM[10'h71][0];	// lsu.scala:210:16
        ldq_6_bits_uop_prs2_busy = _RANDOM[10'h71][1];	// lsu.scala:210:16
        ldq_6_bits_uop_prs3_busy = _RANDOM[10'h71][2];	// lsu.scala:210:16
        ldq_6_bits_uop_ppred_busy = _RANDOM[10'h71][3];	// lsu.scala:210:16
        ldq_6_bits_uop_stale_pdst = _RANDOM[10'h71][10:4];	// lsu.scala:210:16
        ldq_6_bits_uop_exception = _RANDOM[10'h71][11];	// lsu.scala:210:16
        ldq_6_bits_uop_exc_cause =
          {_RANDOM[10'h71][31:12], _RANDOM[10'h72], _RANDOM[10'h73][11:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_bypassable = _RANDOM[10'h73][12];	// lsu.scala:210:16
        ldq_6_bits_uop_mem_cmd = _RANDOM[10'h73][17:13];	// lsu.scala:210:16
        ldq_6_bits_uop_mem_size = _RANDOM[10'h73][19:18];	// lsu.scala:210:16
        ldq_6_bits_uop_mem_signed = _RANDOM[10'h73][20];	// lsu.scala:210:16
        ldq_6_bits_uop_is_fence = _RANDOM[10'h73][21];	// lsu.scala:210:16
        ldq_6_bits_uop_is_fencei = _RANDOM[10'h73][22];	// lsu.scala:210:16
        ldq_6_bits_uop_is_amo = _RANDOM[10'h73][23];	// lsu.scala:210:16
        ldq_6_bits_uop_uses_ldq = _RANDOM[10'h73][24];	// lsu.scala:210:16
        ldq_6_bits_uop_uses_stq = _RANDOM[10'h73][25];	// lsu.scala:210:16
        ldq_6_bits_uop_is_sys_pc2epc = _RANDOM[10'h73][26];	// lsu.scala:210:16
        ldq_6_bits_uop_is_unique = _RANDOM[10'h73][27];	// lsu.scala:210:16
        ldq_6_bits_uop_flush_on_commit = _RANDOM[10'h73][28];	// lsu.scala:210:16
        ldq_6_bits_uop_ldst_is_rs1 = _RANDOM[10'h73][29];	// lsu.scala:210:16
        ldq_6_bits_uop_ldst = {_RANDOM[10'h73][31:30], _RANDOM[10'h74][3:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_lrs1 = _RANDOM[10'h74][9:4];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs2 = _RANDOM[10'h74][15:10];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs3 = _RANDOM[10'h74][21:16];	// lsu.scala:210:16
        ldq_6_bits_uop_ldst_val = _RANDOM[10'h74][22];	// lsu.scala:210:16
        ldq_6_bits_uop_dst_rtype = _RANDOM[10'h74][24:23];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs1_rtype = _RANDOM[10'h74][26:25];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs2_rtype = _RANDOM[10'h74][28:27];	// lsu.scala:210:16
        ldq_6_bits_uop_frs3_en = _RANDOM[10'h74][29];	// lsu.scala:210:16
        ldq_6_bits_uop_fp_val = _RANDOM[10'h74][30];	// lsu.scala:210:16
        ldq_6_bits_uop_fp_single = _RANDOM[10'h74][31];	// lsu.scala:210:16
        ldq_6_bits_uop_xcpt_pf_if = _RANDOM[10'h75][0];	// lsu.scala:210:16
        ldq_6_bits_uop_xcpt_ae_if = _RANDOM[10'h75][1];	// lsu.scala:210:16
        ldq_6_bits_uop_xcpt_ma_if = _RANDOM[10'h75][2];	// lsu.scala:210:16
        ldq_6_bits_uop_bp_debug_if = _RANDOM[10'h75][3];	// lsu.scala:210:16
        ldq_6_bits_uop_bp_xcpt_if = _RANDOM[10'h75][4];	// lsu.scala:210:16
        ldq_6_bits_uop_debug_fsrc = _RANDOM[10'h75][6:5];	// lsu.scala:210:16
        ldq_6_bits_uop_debug_tsrc = _RANDOM[10'h75][8:7];	// lsu.scala:210:16
        ldq_6_bits_addr_valid = _RANDOM[10'h75][9];	// lsu.scala:210:16
        ldq_6_bits_addr_bits = {_RANDOM[10'h75][31:10], _RANDOM[10'h76][17:0]};	// lsu.scala:210:16
        ldq_6_bits_addr_is_virtual = _RANDOM[10'h76][18];	// lsu.scala:210:16
        ldq_6_bits_addr_is_uncacheable = _RANDOM[10'h76][19];	// lsu.scala:210:16
        ldq_6_bits_executed = _RANDOM[10'h76][20];	// lsu.scala:210:16
        ldq_6_bits_succeeded = _RANDOM[10'h76][21];	// lsu.scala:210:16
        ldq_6_bits_order_fail = _RANDOM[10'h76][22];	// lsu.scala:210:16
        ldq_6_bits_observed = _RANDOM[10'h76][23];	// lsu.scala:210:16
        ldq_6_bits_st_dep_mask = {_RANDOM[10'h76][31:24], _RANDOM[10'h77][15:0]};	// lsu.scala:210:16
        ldq_6_bits_youngest_stq_idx = _RANDOM[10'h77][20:16];	// lsu.scala:210:16
        ldq_6_bits_forward_std_val = _RANDOM[10'h77][21];	// lsu.scala:210:16
        ldq_6_bits_forward_stq_idx = _RANDOM[10'h77][26:22];	// lsu.scala:210:16
        ldq_7_valid = _RANDOM[10'h79][27];	// lsu.scala:210:16
        ldq_7_bits_uop_uopc = {_RANDOM[10'h79][31:28], _RANDOM[10'h7A][2:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_inst = {_RANDOM[10'h7A][31:3], _RANDOM[10'h7B][2:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_debug_inst = {_RANDOM[10'h7B][31:3], _RANDOM[10'h7C][2:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_is_rvc = _RANDOM[10'h7C][3];	// lsu.scala:210:16
        ldq_7_bits_uop_debug_pc = {_RANDOM[10'h7C][31:4], _RANDOM[10'h7D][11:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_iq_type = _RANDOM[10'h7D][14:12];	// lsu.scala:210:16
        ldq_7_bits_uop_fu_code = _RANDOM[10'h7D][24:15];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_br_type = _RANDOM[10'h7D][28:25];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_op1_sel = _RANDOM[10'h7D][30:29];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_op2_sel = {_RANDOM[10'h7D][31], _RANDOM[10'h7E][1:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_imm_sel = _RANDOM[10'h7E][4:2];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_op_fcn = _RANDOM[10'h7E][8:5];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_fcn_dw = _RANDOM[10'h7E][9];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_csr_cmd = _RANDOM[10'h7E][12:10];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_is_load = _RANDOM[10'h7E][13];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_is_sta = _RANDOM[10'h7E][14];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_is_std = _RANDOM[10'h7E][15];	// lsu.scala:210:16
        ldq_7_bits_uop_iw_state = _RANDOM[10'h7E][17:16];	// lsu.scala:210:16
        ldq_7_bits_uop_iw_p1_poisoned = _RANDOM[10'h7E][18];	// lsu.scala:210:16
        ldq_7_bits_uop_iw_p2_poisoned = _RANDOM[10'h7E][19];	// lsu.scala:210:16
        ldq_7_bits_uop_is_br = _RANDOM[10'h7E][20];	// lsu.scala:210:16
        ldq_7_bits_uop_is_jalr = _RANDOM[10'h7E][21];	// lsu.scala:210:16
        ldq_7_bits_uop_is_jal = _RANDOM[10'h7E][22];	// lsu.scala:210:16
        ldq_7_bits_uop_is_sfb = _RANDOM[10'h7E][23];	// lsu.scala:210:16
        ldq_7_bits_uop_br_mask = {_RANDOM[10'h7E][31:24], _RANDOM[10'h7F][7:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_br_tag = _RANDOM[10'h7F][11:8];	// lsu.scala:210:16
        ldq_7_bits_uop_ftq_idx = _RANDOM[10'h7F][16:12];	// lsu.scala:210:16
        ldq_7_bits_uop_edge_inst = _RANDOM[10'h7F][17];	// lsu.scala:210:16
        ldq_7_bits_uop_pc_lob = _RANDOM[10'h7F][23:18];	// lsu.scala:210:16
        ldq_7_bits_uop_taken = _RANDOM[10'h7F][24];	// lsu.scala:210:16
        ldq_7_bits_uop_imm_packed = {_RANDOM[10'h7F][31:25], _RANDOM[10'h80][12:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_csr_addr = _RANDOM[10'h80][24:13];	// lsu.scala:210:16
        ldq_7_bits_uop_rob_idx = _RANDOM[10'h80][31:25];	// lsu.scala:210:16
        ldq_7_bits_uop_ldq_idx = _RANDOM[10'h81][4:0];	// lsu.scala:210:16
        ldq_7_bits_uop_stq_idx = _RANDOM[10'h81][9:5];	// lsu.scala:210:16
        ldq_7_bits_uop_rxq_idx = _RANDOM[10'h81][11:10];	// lsu.scala:210:16
        ldq_7_bits_uop_pdst = _RANDOM[10'h81][18:12];	// lsu.scala:210:16
        ldq_7_bits_uop_prs1 = _RANDOM[10'h81][25:19];	// lsu.scala:210:16
        ldq_7_bits_uop_prs2 = {_RANDOM[10'h81][31:26], _RANDOM[10'h82][0]};	// lsu.scala:210:16
        ldq_7_bits_uop_prs3 = _RANDOM[10'h82][7:1];	// lsu.scala:210:16
        ldq_7_bits_uop_ppred = _RANDOM[10'h82][12:8];	// lsu.scala:210:16
        ldq_7_bits_uop_prs1_busy = _RANDOM[10'h82][13];	// lsu.scala:210:16
        ldq_7_bits_uop_prs2_busy = _RANDOM[10'h82][14];	// lsu.scala:210:16
        ldq_7_bits_uop_prs3_busy = _RANDOM[10'h82][15];	// lsu.scala:210:16
        ldq_7_bits_uop_ppred_busy = _RANDOM[10'h82][16];	// lsu.scala:210:16
        ldq_7_bits_uop_stale_pdst = _RANDOM[10'h82][23:17];	// lsu.scala:210:16
        ldq_7_bits_uop_exception = _RANDOM[10'h82][24];	// lsu.scala:210:16
        ldq_7_bits_uop_exc_cause =
          {_RANDOM[10'h82][31:25], _RANDOM[10'h83], _RANDOM[10'h84][24:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_bypassable = _RANDOM[10'h84][25];	// lsu.scala:210:16
        ldq_7_bits_uop_mem_cmd = _RANDOM[10'h84][30:26];	// lsu.scala:210:16
        ldq_7_bits_uop_mem_size = {_RANDOM[10'h84][31], _RANDOM[10'h85][0]};	// lsu.scala:210:16
        ldq_7_bits_uop_mem_signed = _RANDOM[10'h85][1];	// lsu.scala:210:16
        ldq_7_bits_uop_is_fence = _RANDOM[10'h85][2];	// lsu.scala:210:16
        ldq_7_bits_uop_is_fencei = _RANDOM[10'h85][3];	// lsu.scala:210:16
        ldq_7_bits_uop_is_amo = _RANDOM[10'h85][4];	// lsu.scala:210:16
        ldq_7_bits_uop_uses_ldq = _RANDOM[10'h85][5];	// lsu.scala:210:16
        ldq_7_bits_uop_uses_stq = _RANDOM[10'h85][6];	// lsu.scala:210:16
        ldq_7_bits_uop_is_sys_pc2epc = _RANDOM[10'h85][7];	// lsu.scala:210:16
        ldq_7_bits_uop_is_unique = _RANDOM[10'h85][8];	// lsu.scala:210:16
        ldq_7_bits_uop_flush_on_commit = _RANDOM[10'h85][9];	// lsu.scala:210:16
        ldq_7_bits_uop_ldst_is_rs1 = _RANDOM[10'h85][10];	// lsu.scala:210:16
        ldq_7_bits_uop_ldst = _RANDOM[10'h85][16:11];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs1 = _RANDOM[10'h85][22:17];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs2 = _RANDOM[10'h85][28:23];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs3 = {_RANDOM[10'h85][31:29], _RANDOM[10'h86][2:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_ldst_val = _RANDOM[10'h86][3];	// lsu.scala:210:16
        ldq_7_bits_uop_dst_rtype = _RANDOM[10'h86][5:4];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs1_rtype = _RANDOM[10'h86][7:6];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs2_rtype = _RANDOM[10'h86][9:8];	// lsu.scala:210:16
        ldq_7_bits_uop_frs3_en = _RANDOM[10'h86][10];	// lsu.scala:210:16
        ldq_7_bits_uop_fp_val = _RANDOM[10'h86][11];	// lsu.scala:210:16
        ldq_7_bits_uop_fp_single = _RANDOM[10'h86][12];	// lsu.scala:210:16
        ldq_7_bits_uop_xcpt_pf_if = _RANDOM[10'h86][13];	// lsu.scala:210:16
        ldq_7_bits_uop_xcpt_ae_if = _RANDOM[10'h86][14];	// lsu.scala:210:16
        ldq_7_bits_uop_xcpt_ma_if = _RANDOM[10'h86][15];	// lsu.scala:210:16
        ldq_7_bits_uop_bp_debug_if = _RANDOM[10'h86][16];	// lsu.scala:210:16
        ldq_7_bits_uop_bp_xcpt_if = _RANDOM[10'h86][17];	// lsu.scala:210:16
        ldq_7_bits_uop_debug_fsrc = _RANDOM[10'h86][19:18];	// lsu.scala:210:16
        ldq_7_bits_uop_debug_tsrc = _RANDOM[10'h86][21:20];	// lsu.scala:210:16
        ldq_7_bits_addr_valid = _RANDOM[10'h86][22];	// lsu.scala:210:16
        ldq_7_bits_addr_bits = {_RANDOM[10'h86][31:23], _RANDOM[10'h87][30:0]};	// lsu.scala:210:16
        ldq_7_bits_addr_is_virtual = _RANDOM[10'h87][31];	// lsu.scala:210:16
        ldq_7_bits_addr_is_uncacheable = _RANDOM[10'h88][0];	// lsu.scala:210:16
        ldq_7_bits_executed = _RANDOM[10'h88][1];	// lsu.scala:210:16
        ldq_7_bits_succeeded = _RANDOM[10'h88][2];	// lsu.scala:210:16
        ldq_7_bits_order_fail = _RANDOM[10'h88][3];	// lsu.scala:210:16
        ldq_7_bits_observed = _RANDOM[10'h88][4];	// lsu.scala:210:16
        ldq_7_bits_st_dep_mask = _RANDOM[10'h88][28:5];	// lsu.scala:210:16
        ldq_7_bits_youngest_stq_idx = {_RANDOM[10'h88][31:29], _RANDOM[10'h89][1:0]};	// lsu.scala:210:16
        ldq_7_bits_forward_std_val = _RANDOM[10'h89][2];	// lsu.scala:210:16
        ldq_7_bits_forward_stq_idx = _RANDOM[10'h89][7:3];	// lsu.scala:210:16
        ldq_8_valid = _RANDOM[10'h8B][8];	// lsu.scala:210:16
        ldq_8_bits_uop_uopc = _RANDOM[10'h8B][15:9];	// lsu.scala:210:16
        ldq_8_bits_uop_inst = {_RANDOM[10'h8B][31:16], _RANDOM[10'h8C][15:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_debug_inst = {_RANDOM[10'h8C][31:16], _RANDOM[10'h8D][15:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_is_rvc = _RANDOM[10'h8D][16];	// lsu.scala:210:16
        ldq_8_bits_uop_debug_pc = {_RANDOM[10'h8D][31:17], _RANDOM[10'h8E][24:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_iq_type = _RANDOM[10'h8E][27:25];	// lsu.scala:210:16
        ldq_8_bits_uop_fu_code = {_RANDOM[10'h8E][31:28], _RANDOM[10'h8F][5:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_br_type = _RANDOM[10'h8F][9:6];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_op1_sel = _RANDOM[10'h8F][11:10];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_op2_sel = _RANDOM[10'h8F][14:12];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_imm_sel = _RANDOM[10'h8F][17:15];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_op_fcn = _RANDOM[10'h8F][21:18];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_fcn_dw = _RANDOM[10'h8F][22];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_csr_cmd = _RANDOM[10'h8F][25:23];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_is_load = _RANDOM[10'h8F][26];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_is_sta = _RANDOM[10'h8F][27];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_is_std = _RANDOM[10'h8F][28];	// lsu.scala:210:16
        ldq_8_bits_uop_iw_state = _RANDOM[10'h8F][30:29];	// lsu.scala:210:16
        ldq_8_bits_uop_iw_p1_poisoned = _RANDOM[10'h8F][31];	// lsu.scala:210:16
        ldq_8_bits_uop_iw_p2_poisoned = _RANDOM[10'h90][0];	// lsu.scala:210:16
        ldq_8_bits_uop_is_br = _RANDOM[10'h90][1];	// lsu.scala:210:16
        ldq_8_bits_uop_is_jalr = _RANDOM[10'h90][2];	// lsu.scala:210:16
        ldq_8_bits_uop_is_jal = _RANDOM[10'h90][3];	// lsu.scala:210:16
        ldq_8_bits_uop_is_sfb = _RANDOM[10'h90][4];	// lsu.scala:210:16
        ldq_8_bits_uop_br_mask = _RANDOM[10'h90][20:5];	// lsu.scala:210:16
        ldq_8_bits_uop_br_tag = _RANDOM[10'h90][24:21];	// lsu.scala:210:16
        ldq_8_bits_uop_ftq_idx = _RANDOM[10'h90][29:25];	// lsu.scala:210:16
        ldq_8_bits_uop_edge_inst = _RANDOM[10'h90][30];	// lsu.scala:210:16
        ldq_8_bits_uop_pc_lob = {_RANDOM[10'h90][31], _RANDOM[10'h91][4:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_taken = _RANDOM[10'h91][5];	// lsu.scala:210:16
        ldq_8_bits_uop_imm_packed = _RANDOM[10'h91][25:6];	// lsu.scala:210:16
        ldq_8_bits_uop_csr_addr = {_RANDOM[10'h91][31:26], _RANDOM[10'h92][5:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_rob_idx = _RANDOM[10'h92][12:6];	// lsu.scala:210:16
        ldq_8_bits_uop_ldq_idx = _RANDOM[10'h92][17:13];	// lsu.scala:210:16
        ldq_8_bits_uop_stq_idx = _RANDOM[10'h92][22:18];	// lsu.scala:210:16
        ldq_8_bits_uop_rxq_idx = _RANDOM[10'h92][24:23];	// lsu.scala:210:16
        ldq_8_bits_uop_pdst = _RANDOM[10'h92][31:25];	// lsu.scala:210:16
        ldq_8_bits_uop_prs1 = _RANDOM[10'h93][6:0];	// lsu.scala:210:16
        ldq_8_bits_uop_prs2 = _RANDOM[10'h93][13:7];	// lsu.scala:210:16
        ldq_8_bits_uop_prs3 = _RANDOM[10'h93][20:14];	// lsu.scala:210:16
        ldq_8_bits_uop_ppred = _RANDOM[10'h93][25:21];	// lsu.scala:210:16
        ldq_8_bits_uop_prs1_busy = _RANDOM[10'h93][26];	// lsu.scala:210:16
        ldq_8_bits_uop_prs2_busy = _RANDOM[10'h93][27];	// lsu.scala:210:16
        ldq_8_bits_uop_prs3_busy = _RANDOM[10'h93][28];	// lsu.scala:210:16
        ldq_8_bits_uop_ppred_busy = _RANDOM[10'h93][29];	// lsu.scala:210:16
        ldq_8_bits_uop_stale_pdst = {_RANDOM[10'h93][31:30], _RANDOM[10'h94][4:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_exception = _RANDOM[10'h94][5];	// lsu.scala:210:16
        ldq_8_bits_uop_exc_cause =
          {_RANDOM[10'h94][31:6], _RANDOM[10'h95], _RANDOM[10'h96][5:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_bypassable = _RANDOM[10'h96][6];	// lsu.scala:210:16
        ldq_8_bits_uop_mem_cmd = _RANDOM[10'h96][11:7];	// lsu.scala:210:16
        ldq_8_bits_uop_mem_size = _RANDOM[10'h96][13:12];	// lsu.scala:210:16
        ldq_8_bits_uop_mem_signed = _RANDOM[10'h96][14];	// lsu.scala:210:16
        ldq_8_bits_uop_is_fence = _RANDOM[10'h96][15];	// lsu.scala:210:16
        ldq_8_bits_uop_is_fencei = _RANDOM[10'h96][16];	// lsu.scala:210:16
        ldq_8_bits_uop_is_amo = _RANDOM[10'h96][17];	// lsu.scala:210:16
        ldq_8_bits_uop_uses_ldq = _RANDOM[10'h96][18];	// lsu.scala:210:16
        ldq_8_bits_uop_uses_stq = _RANDOM[10'h96][19];	// lsu.scala:210:16
        ldq_8_bits_uop_is_sys_pc2epc = _RANDOM[10'h96][20];	// lsu.scala:210:16
        ldq_8_bits_uop_is_unique = _RANDOM[10'h96][21];	// lsu.scala:210:16
        ldq_8_bits_uop_flush_on_commit = _RANDOM[10'h96][22];	// lsu.scala:210:16
        ldq_8_bits_uop_ldst_is_rs1 = _RANDOM[10'h96][23];	// lsu.scala:210:16
        ldq_8_bits_uop_ldst = _RANDOM[10'h96][29:24];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs1 = {_RANDOM[10'h96][31:30], _RANDOM[10'h97][3:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_lrs2 = _RANDOM[10'h97][9:4];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs3 = _RANDOM[10'h97][15:10];	// lsu.scala:210:16
        ldq_8_bits_uop_ldst_val = _RANDOM[10'h97][16];	// lsu.scala:210:16
        ldq_8_bits_uop_dst_rtype = _RANDOM[10'h97][18:17];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs1_rtype = _RANDOM[10'h97][20:19];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs2_rtype = _RANDOM[10'h97][22:21];	// lsu.scala:210:16
        ldq_8_bits_uop_frs3_en = _RANDOM[10'h97][23];	// lsu.scala:210:16
        ldq_8_bits_uop_fp_val = _RANDOM[10'h97][24];	// lsu.scala:210:16
        ldq_8_bits_uop_fp_single = _RANDOM[10'h97][25];	// lsu.scala:210:16
        ldq_8_bits_uop_xcpt_pf_if = _RANDOM[10'h97][26];	// lsu.scala:210:16
        ldq_8_bits_uop_xcpt_ae_if = _RANDOM[10'h97][27];	// lsu.scala:210:16
        ldq_8_bits_uop_xcpt_ma_if = _RANDOM[10'h97][28];	// lsu.scala:210:16
        ldq_8_bits_uop_bp_debug_if = _RANDOM[10'h97][29];	// lsu.scala:210:16
        ldq_8_bits_uop_bp_xcpt_if = _RANDOM[10'h97][30];	// lsu.scala:210:16
        ldq_8_bits_uop_debug_fsrc = {_RANDOM[10'h97][31], _RANDOM[10'h98][0]};	// lsu.scala:210:16
        ldq_8_bits_uop_debug_tsrc = _RANDOM[10'h98][2:1];	// lsu.scala:210:16
        ldq_8_bits_addr_valid = _RANDOM[10'h98][3];	// lsu.scala:210:16
        ldq_8_bits_addr_bits = {_RANDOM[10'h98][31:4], _RANDOM[10'h99][11:0]};	// lsu.scala:210:16
        ldq_8_bits_addr_is_virtual = _RANDOM[10'h99][12];	// lsu.scala:210:16
        ldq_8_bits_addr_is_uncacheable = _RANDOM[10'h99][13];	// lsu.scala:210:16
        ldq_8_bits_executed = _RANDOM[10'h99][14];	// lsu.scala:210:16
        ldq_8_bits_succeeded = _RANDOM[10'h99][15];	// lsu.scala:210:16
        ldq_8_bits_order_fail = _RANDOM[10'h99][16];	// lsu.scala:210:16
        ldq_8_bits_observed = _RANDOM[10'h99][17];	// lsu.scala:210:16
        ldq_8_bits_st_dep_mask = {_RANDOM[10'h99][31:18], _RANDOM[10'h9A][9:0]};	// lsu.scala:210:16
        ldq_8_bits_youngest_stq_idx = _RANDOM[10'h9A][14:10];	// lsu.scala:210:16
        ldq_8_bits_forward_std_val = _RANDOM[10'h9A][15];	// lsu.scala:210:16
        ldq_8_bits_forward_stq_idx = _RANDOM[10'h9A][20:16];	// lsu.scala:210:16
        ldq_9_valid = _RANDOM[10'h9C][21];	// lsu.scala:210:16
        ldq_9_bits_uop_uopc = _RANDOM[10'h9C][28:22];	// lsu.scala:210:16
        ldq_9_bits_uop_inst = {_RANDOM[10'h9C][31:29], _RANDOM[10'h9D][28:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_debug_inst = {_RANDOM[10'h9D][31:29], _RANDOM[10'h9E][28:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_is_rvc = _RANDOM[10'h9E][29];	// lsu.scala:210:16
        ldq_9_bits_uop_debug_pc =
          {_RANDOM[10'h9E][31:30], _RANDOM[10'h9F], _RANDOM[10'hA0][5:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_iq_type = _RANDOM[10'hA0][8:6];	// lsu.scala:210:16
        ldq_9_bits_uop_fu_code = _RANDOM[10'hA0][18:9];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_br_type = _RANDOM[10'hA0][22:19];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_op1_sel = _RANDOM[10'hA0][24:23];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_op2_sel = _RANDOM[10'hA0][27:25];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_imm_sel = _RANDOM[10'hA0][30:28];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_op_fcn = {_RANDOM[10'hA0][31], _RANDOM[10'hA1][2:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_fcn_dw = _RANDOM[10'hA1][3];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_csr_cmd = _RANDOM[10'hA1][6:4];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_is_load = _RANDOM[10'hA1][7];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_is_sta = _RANDOM[10'hA1][8];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_is_std = _RANDOM[10'hA1][9];	// lsu.scala:210:16
        ldq_9_bits_uop_iw_state = _RANDOM[10'hA1][11:10];	// lsu.scala:210:16
        ldq_9_bits_uop_iw_p1_poisoned = _RANDOM[10'hA1][12];	// lsu.scala:210:16
        ldq_9_bits_uop_iw_p2_poisoned = _RANDOM[10'hA1][13];	// lsu.scala:210:16
        ldq_9_bits_uop_is_br = _RANDOM[10'hA1][14];	// lsu.scala:210:16
        ldq_9_bits_uop_is_jalr = _RANDOM[10'hA1][15];	// lsu.scala:210:16
        ldq_9_bits_uop_is_jal = _RANDOM[10'hA1][16];	// lsu.scala:210:16
        ldq_9_bits_uop_is_sfb = _RANDOM[10'hA1][17];	// lsu.scala:210:16
        ldq_9_bits_uop_br_mask = {_RANDOM[10'hA1][31:18], _RANDOM[10'hA2][1:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_br_tag = _RANDOM[10'hA2][5:2];	// lsu.scala:210:16
        ldq_9_bits_uop_ftq_idx = _RANDOM[10'hA2][10:6];	// lsu.scala:210:16
        ldq_9_bits_uop_edge_inst = _RANDOM[10'hA2][11];	// lsu.scala:210:16
        ldq_9_bits_uop_pc_lob = _RANDOM[10'hA2][17:12];	// lsu.scala:210:16
        ldq_9_bits_uop_taken = _RANDOM[10'hA2][18];	// lsu.scala:210:16
        ldq_9_bits_uop_imm_packed = {_RANDOM[10'hA2][31:19], _RANDOM[10'hA3][6:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_csr_addr = _RANDOM[10'hA3][18:7];	// lsu.scala:210:16
        ldq_9_bits_uop_rob_idx = _RANDOM[10'hA3][25:19];	// lsu.scala:210:16
        ldq_9_bits_uop_ldq_idx = _RANDOM[10'hA3][30:26];	// lsu.scala:210:16
        ldq_9_bits_uop_stq_idx = {_RANDOM[10'hA3][31], _RANDOM[10'hA4][3:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_rxq_idx = _RANDOM[10'hA4][5:4];	// lsu.scala:210:16
        ldq_9_bits_uop_pdst = _RANDOM[10'hA4][12:6];	// lsu.scala:210:16
        ldq_9_bits_uop_prs1 = _RANDOM[10'hA4][19:13];	// lsu.scala:210:16
        ldq_9_bits_uop_prs2 = _RANDOM[10'hA4][26:20];	// lsu.scala:210:16
        ldq_9_bits_uop_prs3 = {_RANDOM[10'hA4][31:27], _RANDOM[10'hA5][1:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_ppred = _RANDOM[10'hA5][6:2];	// lsu.scala:210:16
        ldq_9_bits_uop_prs1_busy = _RANDOM[10'hA5][7];	// lsu.scala:210:16
        ldq_9_bits_uop_prs2_busy = _RANDOM[10'hA5][8];	// lsu.scala:210:16
        ldq_9_bits_uop_prs3_busy = _RANDOM[10'hA5][9];	// lsu.scala:210:16
        ldq_9_bits_uop_ppred_busy = _RANDOM[10'hA5][10];	// lsu.scala:210:16
        ldq_9_bits_uop_stale_pdst = _RANDOM[10'hA5][17:11];	// lsu.scala:210:16
        ldq_9_bits_uop_exception = _RANDOM[10'hA5][18];	// lsu.scala:210:16
        ldq_9_bits_uop_exc_cause =
          {_RANDOM[10'hA5][31:19], _RANDOM[10'hA6], _RANDOM[10'hA7][18:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_bypassable = _RANDOM[10'hA7][19];	// lsu.scala:210:16
        ldq_9_bits_uop_mem_cmd = _RANDOM[10'hA7][24:20];	// lsu.scala:210:16
        ldq_9_bits_uop_mem_size = _RANDOM[10'hA7][26:25];	// lsu.scala:210:16
        ldq_9_bits_uop_mem_signed = _RANDOM[10'hA7][27];	// lsu.scala:210:16
        ldq_9_bits_uop_is_fence = _RANDOM[10'hA7][28];	// lsu.scala:210:16
        ldq_9_bits_uop_is_fencei = _RANDOM[10'hA7][29];	// lsu.scala:210:16
        ldq_9_bits_uop_is_amo = _RANDOM[10'hA7][30];	// lsu.scala:210:16
        ldq_9_bits_uop_uses_ldq = _RANDOM[10'hA7][31];	// lsu.scala:210:16
        ldq_9_bits_uop_uses_stq = _RANDOM[10'hA8][0];	// lsu.scala:210:16
        ldq_9_bits_uop_is_sys_pc2epc = _RANDOM[10'hA8][1];	// lsu.scala:210:16
        ldq_9_bits_uop_is_unique = _RANDOM[10'hA8][2];	// lsu.scala:210:16
        ldq_9_bits_uop_flush_on_commit = _RANDOM[10'hA8][3];	// lsu.scala:210:16
        ldq_9_bits_uop_ldst_is_rs1 = _RANDOM[10'hA8][4];	// lsu.scala:210:16
        ldq_9_bits_uop_ldst = _RANDOM[10'hA8][10:5];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs1 = _RANDOM[10'hA8][16:11];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs2 = _RANDOM[10'hA8][22:17];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs3 = _RANDOM[10'hA8][28:23];	// lsu.scala:210:16
        ldq_9_bits_uop_ldst_val = _RANDOM[10'hA8][29];	// lsu.scala:210:16
        ldq_9_bits_uop_dst_rtype = _RANDOM[10'hA8][31:30];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs1_rtype = _RANDOM[10'hA9][1:0];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs2_rtype = _RANDOM[10'hA9][3:2];	// lsu.scala:210:16
        ldq_9_bits_uop_frs3_en = _RANDOM[10'hA9][4];	// lsu.scala:210:16
        ldq_9_bits_uop_fp_val = _RANDOM[10'hA9][5];	// lsu.scala:210:16
        ldq_9_bits_uop_fp_single = _RANDOM[10'hA9][6];	// lsu.scala:210:16
        ldq_9_bits_uop_xcpt_pf_if = _RANDOM[10'hA9][7];	// lsu.scala:210:16
        ldq_9_bits_uop_xcpt_ae_if = _RANDOM[10'hA9][8];	// lsu.scala:210:16
        ldq_9_bits_uop_xcpt_ma_if = _RANDOM[10'hA9][9];	// lsu.scala:210:16
        ldq_9_bits_uop_bp_debug_if = _RANDOM[10'hA9][10];	// lsu.scala:210:16
        ldq_9_bits_uop_bp_xcpt_if = _RANDOM[10'hA9][11];	// lsu.scala:210:16
        ldq_9_bits_uop_debug_fsrc = _RANDOM[10'hA9][13:12];	// lsu.scala:210:16
        ldq_9_bits_uop_debug_tsrc = _RANDOM[10'hA9][15:14];	// lsu.scala:210:16
        ldq_9_bits_addr_valid = _RANDOM[10'hA9][16];	// lsu.scala:210:16
        ldq_9_bits_addr_bits = {_RANDOM[10'hA9][31:17], _RANDOM[10'hAA][24:0]};	// lsu.scala:210:16
        ldq_9_bits_addr_is_virtual = _RANDOM[10'hAA][25];	// lsu.scala:210:16
        ldq_9_bits_addr_is_uncacheable = _RANDOM[10'hAA][26];	// lsu.scala:210:16
        ldq_9_bits_executed = _RANDOM[10'hAA][27];	// lsu.scala:210:16
        ldq_9_bits_succeeded = _RANDOM[10'hAA][28];	// lsu.scala:210:16
        ldq_9_bits_order_fail = _RANDOM[10'hAA][29];	// lsu.scala:210:16
        ldq_9_bits_observed = _RANDOM[10'hAA][30];	// lsu.scala:210:16
        ldq_9_bits_st_dep_mask = {_RANDOM[10'hAA][31], _RANDOM[10'hAB][22:0]};	// lsu.scala:210:16
        ldq_9_bits_youngest_stq_idx = _RANDOM[10'hAB][27:23];	// lsu.scala:210:16
        ldq_9_bits_forward_std_val = _RANDOM[10'hAB][28];	// lsu.scala:210:16
        ldq_9_bits_forward_stq_idx = {_RANDOM[10'hAB][31:29], _RANDOM[10'hAC][1:0]};	// lsu.scala:210:16
        ldq_10_valid = _RANDOM[10'hAE][2];	// lsu.scala:210:16
        ldq_10_bits_uop_uopc = _RANDOM[10'hAE][9:3];	// lsu.scala:210:16
        ldq_10_bits_uop_inst = {_RANDOM[10'hAE][31:10], _RANDOM[10'hAF][9:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_debug_inst = {_RANDOM[10'hAF][31:10], _RANDOM[10'hB0][9:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_is_rvc = _RANDOM[10'hB0][10];	// lsu.scala:210:16
        ldq_10_bits_uop_debug_pc = {_RANDOM[10'hB0][31:11], _RANDOM[10'hB1][18:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_iq_type = _RANDOM[10'hB1][21:19];	// lsu.scala:210:16
        ldq_10_bits_uop_fu_code = _RANDOM[10'hB1][31:22];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_br_type = _RANDOM[10'hB2][3:0];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_op1_sel = _RANDOM[10'hB2][5:4];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_op2_sel = _RANDOM[10'hB2][8:6];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_imm_sel = _RANDOM[10'hB2][11:9];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_op_fcn = _RANDOM[10'hB2][15:12];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_fcn_dw = _RANDOM[10'hB2][16];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_csr_cmd = _RANDOM[10'hB2][19:17];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_is_load = _RANDOM[10'hB2][20];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_is_sta = _RANDOM[10'hB2][21];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_is_std = _RANDOM[10'hB2][22];	// lsu.scala:210:16
        ldq_10_bits_uop_iw_state = _RANDOM[10'hB2][24:23];	// lsu.scala:210:16
        ldq_10_bits_uop_iw_p1_poisoned = _RANDOM[10'hB2][25];	// lsu.scala:210:16
        ldq_10_bits_uop_iw_p2_poisoned = _RANDOM[10'hB2][26];	// lsu.scala:210:16
        ldq_10_bits_uop_is_br = _RANDOM[10'hB2][27];	// lsu.scala:210:16
        ldq_10_bits_uop_is_jalr = _RANDOM[10'hB2][28];	// lsu.scala:210:16
        ldq_10_bits_uop_is_jal = _RANDOM[10'hB2][29];	// lsu.scala:210:16
        ldq_10_bits_uop_is_sfb = _RANDOM[10'hB2][30];	// lsu.scala:210:16
        ldq_10_bits_uop_br_mask = {_RANDOM[10'hB2][31], _RANDOM[10'hB3][14:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_br_tag = _RANDOM[10'hB3][18:15];	// lsu.scala:210:16
        ldq_10_bits_uop_ftq_idx = _RANDOM[10'hB3][23:19];	// lsu.scala:210:16
        ldq_10_bits_uop_edge_inst = _RANDOM[10'hB3][24];	// lsu.scala:210:16
        ldq_10_bits_uop_pc_lob = _RANDOM[10'hB3][30:25];	// lsu.scala:210:16
        ldq_10_bits_uop_taken = _RANDOM[10'hB3][31];	// lsu.scala:210:16
        ldq_10_bits_uop_imm_packed = _RANDOM[10'hB4][19:0];	// lsu.scala:210:16
        ldq_10_bits_uop_csr_addr = _RANDOM[10'hB4][31:20];	// lsu.scala:210:16
        ldq_10_bits_uop_rob_idx = _RANDOM[10'hB5][6:0];	// lsu.scala:210:16
        ldq_10_bits_uop_ldq_idx = _RANDOM[10'hB5][11:7];	// lsu.scala:210:16
        ldq_10_bits_uop_stq_idx = _RANDOM[10'hB5][16:12];	// lsu.scala:210:16
        ldq_10_bits_uop_rxq_idx = _RANDOM[10'hB5][18:17];	// lsu.scala:210:16
        ldq_10_bits_uop_pdst = _RANDOM[10'hB5][25:19];	// lsu.scala:210:16
        ldq_10_bits_uop_prs1 = {_RANDOM[10'hB5][31:26], _RANDOM[10'hB6][0]};	// lsu.scala:210:16
        ldq_10_bits_uop_prs2 = _RANDOM[10'hB6][7:1];	// lsu.scala:210:16
        ldq_10_bits_uop_prs3 = _RANDOM[10'hB6][14:8];	// lsu.scala:210:16
        ldq_10_bits_uop_ppred = _RANDOM[10'hB6][19:15];	// lsu.scala:210:16
        ldq_10_bits_uop_prs1_busy = _RANDOM[10'hB6][20];	// lsu.scala:210:16
        ldq_10_bits_uop_prs2_busy = _RANDOM[10'hB6][21];	// lsu.scala:210:16
        ldq_10_bits_uop_prs3_busy = _RANDOM[10'hB6][22];	// lsu.scala:210:16
        ldq_10_bits_uop_ppred_busy = _RANDOM[10'hB6][23];	// lsu.scala:210:16
        ldq_10_bits_uop_stale_pdst = _RANDOM[10'hB6][30:24];	// lsu.scala:210:16
        ldq_10_bits_uop_exception = _RANDOM[10'hB6][31];	// lsu.scala:210:16
        ldq_10_bits_uop_exc_cause = {_RANDOM[10'hB7], _RANDOM[10'hB8]};	// lsu.scala:210:16
        ldq_10_bits_uop_bypassable = _RANDOM[10'hB9][0];	// lsu.scala:210:16
        ldq_10_bits_uop_mem_cmd = _RANDOM[10'hB9][5:1];	// lsu.scala:210:16
        ldq_10_bits_uop_mem_size = _RANDOM[10'hB9][7:6];	// lsu.scala:210:16
        ldq_10_bits_uop_mem_signed = _RANDOM[10'hB9][8];	// lsu.scala:210:16
        ldq_10_bits_uop_is_fence = _RANDOM[10'hB9][9];	// lsu.scala:210:16
        ldq_10_bits_uop_is_fencei = _RANDOM[10'hB9][10];	// lsu.scala:210:16
        ldq_10_bits_uop_is_amo = _RANDOM[10'hB9][11];	// lsu.scala:210:16
        ldq_10_bits_uop_uses_ldq = _RANDOM[10'hB9][12];	// lsu.scala:210:16
        ldq_10_bits_uop_uses_stq = _RANDOM[10'hB9][13];	// lsu.scala:210:16
        ldq_10_bits_uop_is_sys_pc2epc = _RANDOM[10'hB9][14];	// lsu.scala:210:16
        ldq_10_bits_uop_is_unique = _RANDOM[10'hB9][15];	// lsu.scala:210:16
        ldq_10_bits_uop_flush_on_commit = _RANDOM[10'hB9][16];	// lsu.scala:210:16
        ldq_10_bits_uop_ldst_is_rs1 = _RANDOM[10'hB9][17];	// lsu.scala:210:16
        ldq_10_bits_uop_ldst = _RANDOM[10'hB9][23:18];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs1 = _RANDOM[10'hB9][29:24];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs2 = {_RANDOM[10'hB9][31:30], _RANDOM[10'hBA][3:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_lrs3 = _RANDOM[10'hBA][9:4];	// lsu.scala:210:16
        ldq_10_bits_uop_ldst_val = _RANDOM[10'hBA][10];	// lsu.scala:210:16
        ldq_10_bits_uop_dst_rtype = _RANDOM[10'hBA][12:11];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs1_rtype = _RANDOM[10'hBA][14:13];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs2_rtype = _RANDOM[10'hBA][16:15];	// lsu.scala:210:16
        ldq_10_bits_uop_frs3_en = _RANDOM[10'hBA][17];	// lsu.scala:210:16
        ldq_10_bits_uop_fp_val = _RANDOM[10'hBA][18];	// lsu.scala:210:16
        ldq_10_bits_uop_fp_single = _RANDOM[10'hBA][19];	// lsu.scala:210:16
        ldq_10_bits_uop_xcpt_pf_if = _RANDOM[10'hBA][20];	// lsu.scala:210:16
        ldq_10_bits_uop_xcpt_ae_if = _RANDOM[10'hBA][21];	// lsu.scala:210:16
        ldq_10_bits_uop_xcpt_ma_if = _RANDOM[10'hBA][22];	// lsu.scala:210:16
        ldq_10_bits_uop_bp_debug_if = _RANDOM[10'hBA][23];	// lsu.scala:210:16
        ldq_10_bits_uop_bp_xcpt_if = _RANDOM[10'hBA][24];	// lsu.scala:210:16
        ldq_10_bits_uop_debug_fsrc = _RANDOM[10'hBA][26:25];	// lsu.scala:210:16
        ldq_10_bits_uop_debug_tsrc = _RANDOM[10'hBA][28:27];	// lsu.scala:210:16
        ldq_10_bits_addr_valid = _RANDOM[10'hBA][29];	// lsu.scala:210:16
        ldq_10_bits_addr_bits =
          {_RANDOM[10'hBA][31:30], _RANDOM[10'hBB], _RANDOM[10'hBC][5:0]};	// lsu.scala:210:16
        ldq_10_bits_addr_is_virtual = _RANDOM[10'hBC][6];	// lsu.scala:210:16
        ldq_10_bits_addr_is_uncacheable = _RANDOM[10'hBC][7];	// lsu.scala:210:16
        ldq_10_bits_executed = _RANDOM[10'hBC][8];	// lsu.scala:210:16
        ldq_10_bits_succeeded = _RANDOM[10'hBC][9];	// lsu.scala:210:16
        ldq_10_bits_order_fail = _RANDOM[10'hBC][10];	// lsu.scala:210:16
        ldq_10_bits_observed = _RANDOM[10'hBC][11];	// lsu.scala:210:16
        ldq_10_bits_st_dep_mask = {_RANDOM[10'hBC][31:12], _RANDOM[10'hBD][3:0]};	// lsu.scala:210:16
        ldq_10_bits_youngest_stq_idx = _RANDOM[10'hBD][8:4];	// lsu.scala:210:16
        ldq_10_bits_forward_std_val = _RANDOM[10'hBD][9];	// lsu.scala:210:16
        ldq_10_bits_forward_stq_idx = _RANDOM[10'hBD][14:10];	// lsu.scala:210:16
        ldq_11_valid = _RANDOM[10'hBF][15];	// lsu.scala:210:16
        ldq_11_bits_uop_uopc = _RANDOM[10'hBF][22:16];	// lsu.scala:210:16
        ldq_11_bits_uop_inst = {_RANDOM[10'hBF][31:23], _RANDOM[10'hC0][22:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_debug_inst = {_RANDOM[10'hC0][31:23], _RANDOM[10'hC1][22:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_is_rvc = _RANDOM[10'hC1][23];	// lsu.scala:210:16
        ldq_11_bits_uop_debug_pc = {_RANDOM[10'hC1][31:24], _RANDOM[10'hC2]};	// lsu.scala:210:16
        ldq_11_bits_uop_iq_type = _RANDOM[10'hC3][2:0];	// lsu.scala:210:16
        ldq_11_bits_uop_fu_code = _RANDOM[10'hC3][12:3];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_br_type = _RANDOM[10'hC3][16:13];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_op1_sel = _RANDOM[10'hC3][18:17];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_op2_sel = _RANDOM[10'hC3][21:19];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_imm_sel = _RANDOM[10'hC3][24:22];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_op_fcn = _RANDOM[10'hC3][28:25];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_fcn_dw = _RANDOM[10'hC3][29];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_csr_cmd = {_RANDOM[10'hC3][31:30], _RANDOM[10'hC4][0]};	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_is_load = _RANDOM[10'hC4][1];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_is_sta = _RANDOM[10'hC4][2];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_is_std = _RANDOM[10'hC4][3];	// lsu.scala:210:16
        ldq_11_bits_uop_iw_state = _RANDOM[10'hC4][5:4];	// lsu.scala:210:16
        ldq_11_bits_uop_iw_p1_poisoned = _RANDOM[10'hC4][6];	// lsu.scala:210:16
        ldq_11_bits_uop_iw_p2_poisoned = _RANDOM[10'hC4][7];	// lsu.scala:210:16
        ldq_11_bits_uop_is_br = _RANDOM[10'hC4][8];	// lsu.scala:210:16
        ldq_11_bits_uop_is_jalr = _RANDOM[10'hC4][9];	// lsu.scala:210:16
        ldq_11_bits_uop_is_jal = _RANDOM[10'hC4][10];	// lsu.scala:210:16
        ldq_11_bits_uop_is_sfb = _RANDOM[10'hC4][11];	// lsu.scala:210:16
        ldq_11_bits_uop_br_mask = _RANDOM[10'hC4][27:12];	// lsu.scala:210:16
        ldq_11_bits_uop_br_tag = _RANDOM[10'hC4][31:28];	// lsu.scala:210:16
        ldq_11_bits_uop_ftq_idx = _RANDOM[10'hC5][4:0];	// lsu.scala:210:16
        ldq_11_bits_uop_edge_inst = _RANDOM[10'hC5][5];	// lsu.scala:210:16
        ldq_11_bits_uop_pc_lob = _RANDOM[10'hC5][11:6];	// lsu.scala:210:16
        ldq_11_bits_uop_taken = _RANDOM[10'hC5][12];	// lsu.scala:210:16
        ldq_11_bits_uop_imm_packed = {_RANDOM[10'hC5][31:13], _RANDOM[10'hC6][0]};	// lsu.scala:210:16
        ldq_11_bits_uop_csr_addr = _RANDOM[10'hC6][12:1];	// lsu.scala:210:16
        ldq_11_bits_uop_rob_idx = _RANDOM[10'hC6][19:13];	// lsu.scala:210:16
        ldq_11_bits_uop_ldq_idx = _RANDOM[10'hC6][24:20];	// lsu.scala:210:16
        ldq_11_bits_uop_stq_idx = _RANDOM[10'hC6][29:25];	// lsu.scala:210:16
        ldq_11_bits_uop_rxq_idx = _RANDOM[10'hC6][31:30];	// lsu.scala:210:16
        ldq_11_bits_uop_pdst = _RANDOM[10'hC7][6:0];	// lsu.scala:210:16
        ldq_11_bits_uop_prs1 = _RANDOM[10'hC7][13:7];	// lsu.scala:210:16
        ldq_11_bits_uop_prs2 = _RANDOM[10'hC7][20:14];	// lsu.scala:210:16
        ldq_11_bits_uop_prs3 = _RANDOM[10'hC7][27:21];	// lsu.scala:210:16
        ldq_11_bits_uop_ppred = {_RANDOM[10'hC7][31:28], _RANDOM[10'hC8][0]};	// lsu.scala:210:16
        ldq_11_bits_uop_prs1_busy = _RANDOM[10'hC8][1];	// lsu.scala:210:16
        ldq_11_bits_uop_prs2_busy = _RANDOM[10'hC8][2];	// lsu.scala:210:16
        ldq_11_bits_uop_prs3_busy = _RANDOM[10'hC8][3];	// lsu.scala:210:16
        ldq_11_bits_uop_ppred_busy = _RANDOM[10'hC8][4];	// lsu.scala:210:16
        ldq_11_bits_uop_stale_pdst = _RANDOM[10'hC8][11:5];	// lsu.scala:210:16
        ldq_11_bits_uop_exception = _RANDOM[10'hC8][12];	// lsu.scala:210:16
        ldq_11_bits_uop_exc_cause =
          {_RANDOM[10'hC8][31:13], _RANDOM[10'hC9], _RANDOM[10'hCA][12:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_bypassable = _RANDOM[10'hCA][13];	// lsu.scala:210:16
        ldq_11_bits_uop_mem_cmd = _RANDOM[10'hCA][18:14];	// lsu.scala:210:16
        ldq_11_bits_uop_mem_size = _RANDOM[10'hCA][20:19];	// lsu.scala:210:16
        ldq_11_bits_uop_mem_signed = _RANDOM[10'hCA][21];	// lsu.scala:210:16
        ldq_11_bits_uop_is_fence = _RANDOM[10'hCA][22];	// lsu.scala:210:16
        ldq_11_bits_uop_is_fencei = _RANDOM[10'hCA][23];	// lsu.scala:210:16
        ldq_11_bits_uop_is_amo = _RANDOM[10'hCA][24];	// lsu.scala:210:16
        ldq_11_bits_uop_uses_ldq = _RANDOM[10'hCA][25];	// lsu.scala:210:16
        ldq_11_bits_uop_uses_stq = _RANDOM[10'hCA][26];	// lsu.scala:210:16
        ldq_11_bits_uop_is_sys_pc2epc = _RANDOM[10'hCA][27];	// lsu.scala:210:16
        ldq_11_bits_uop_is_unique = _RANDOM[10'hCA][28];	// lsu.scala:210:16
        ldq_11_bits_uop_flush_on_commit = _RANDOM[10'hCA][29];	// lsu.scala:210:16
        ldq_11_bits_uop_ldst_is_rs1 = _RANDOM[10'hCA][30];	// lsu.scala:210:16
        ldq_11_bits_uop_ldst = {_RANDOM[10'hCA][31], _RANDOM[10'hCB][4:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_lrs1 = _RANDOM[10'hCB][10:5];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs2 = _RANDOM[10'hCB][16:11];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs3 = _RANDOM[10'hCB][22:17];	// lsu.scala:210:16
        ldq_11_bits_uop_ldst_val = _RANDOM[10'hCB][23];	// lsu.scala:210:16
        ldq_11_bits_uop_dst_rtype = _RANDOM[10'hCB][25:24];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs1_rtype = _RANDOM[10'hCB][27:26];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs2_rtype = _RANDOM[10'hCB][29:28];	// lsu.scala:210:16
        ldq_11_bits_uop_frs3_en = _RANDOM[10'hCB][30];	// lsu.scala:210:16
        ldq_11_bits_uop_fp_val = _RANDOM[10'hCB][31];	// lsu.scala:210:16
        ldq_11_bits_uop_fp_single = _RANDOM[10'hCC][0];	// lsu.scala:210:16
        ldq_11_bits_uop_xcpt_pf_if = _RANDOM[10'hCC][1];	// lsu.scala:210:16
        ldq_11_bits_uop_xcpt_ae_if = _RANDOM[10'hCC][2];	// lsu.scala:210:16
        ldq_11_bits_uop_xcpt_ma_if = _RANDOM[10'hCC][3];	// lsu.scala:210:16
        ldq_11_bits_uop_bp_debug_if = _RANDOM[10'hCC][4];	// lsu.scala:210:16
        ldq_11_bits_uop_bp_xcpt_if = _RANDOM[10'hCC][5];	// lsu.scala:210:16
        ldq_11_bits_uop_debug_fsrc = _RANDOM[10'hCC][7:6];	// lsu.scala:210:16
        ldq_11_bits_uop_debug_tsrc = _RANDOM[10'hCC][9:8];	// lsu.scala:210:16
        ldq_11_bits_addr_valid = _RANDOM[10'hCC][10];	// lsu.scala:210:16
        ldq_11_bits_addr_bits = {_RANDOM[10'hCC][31:11], _RANDOM[10'hCD][18:0]};	// lsu.scala:210:16
        ldq_11_bits_addr_is_virtual = _RANDOM[10'hCD][19];	// lsu.scala:210:16
        ldq_11_bits_addr_is_uncacheable = _RANDOM[10'hCD][20];	// lsu.scala:210:16
        ldq_11_bits_executed = _RANDOM[10'hCD][21];	// lsu.scala:210:16
        ldq_11_bits_succeeded = _RANDOM[10'hCD][22];	// lsu.scala:210:16
        ldq_11_bits_order_fail = _RANDOM[10'hCD][23];	// lsu.scala:210:16
        ldq_11_bits_observed = _RANDOM[10'hCD][24];	// lsu.scala:210:16
        ldq_11_bits_st_dep_mask = {_RANDOM[10'hCD][31:25], _RANDOM[10'hCE][16:0]};	// lsu.scala:210:16
        ldq_11_bits_youngest_stq_idx = _RANDOM[10'hCE][21:17];	// lsu.scala:210:16
        ldq_11_bits_forward_std_val = _RANDOM[10'hCE][22];	// lsu.scala:210:16
        ldq_11_bits_forward_stq_idx = _RANDOM[10'hCE][27:23];	// lsu.scala:210:16
        ldq_12_valid = _RANDOM[10'hD0][28];	// lsu.scala:210:16
        ldq_12_bits_uop_uopc = {_RANDOM[10'hD0][31:29], _RANDOM[10'hD1][3:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_inst = {_RANDOM[10'hD1][31:4], _RANDOM[10'hD2][3:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_debug_inst = {_RANDOM[10'hD2][31:4], _RANDOM[10'hD3][3:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_is_rvc = _RANDOM[10'hD3][4];	// lsu.scala:210:16
        ldq_12_bits_uop_debug_pc = {_RANDOM[10'hD3][31:5], _RANDOM[10'hD4][12:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_iq_type = _RANDOM[10'hD4][15:13];	// lsu.scala:210:16
        ldq_12_bits_uop_fu_code = _RANDOM[10'hD4][25:16];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_br_type = _RANDOM[10'hD4][29:26];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_op1_sel = _RANDOM[10'hD4][31:30];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_op2_sel = _RANDOM[10'hD5][2:0];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_imm_sel = _RANDOM[10'hD5][5:3];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_op_fcn = _RANDOM[10'hD5][9:6];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_fcn_dw = _RANDOM[10'hD5][10];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_csr_cmd = _RANDOM[10'hD5][13:11];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_is_load = _RANDOM[10'hD5][14];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_is_sta = _RANDOM[10'hD5][15];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_is_std = _RANDOM[10'hD5][16];	// lsu.scala:210:16
        ldq_12_bits_uop_iw_state = _RANDOM[10'hD5][18:17];	// lsu.scala:210:16
        ldq_12_bits_uop_iw_p1_poisoned = _RANDOM[10'hD5][19];	// lsu.scala:210:16
        ldq_12_bits_uop_iw_p2_poisoned = _RANDOM[10'hD5][20];	// lsu.scala:210:16
        ldq_12_bits_uop_is_br = _RANDOM[10'hD5][21];	// lsu.scala:210:16
        ldq_12_bits_uop_is_jalr = _RANDOM[10'hD5][22];	// lsu.scala:210:16
        ldq_12_bits_uop_is_jal = _RANDOM[10'hD5][23];	// lsu.scala:210:16
        ldq_12_bits_uop_is_sfb = _RANDOM[10'hD5][24];	// lsu.scala:210:16
        ldq_12_bits_uop_br_mask = {_RANDOM[10'hD5][31:25], _RANDOM[10'hD6][8:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_br_tag = _RANDOM[10'hD6][12:9];	// lsu.scala:210:16
        ldq_12_bits_uop_ftq_idx = _RANDOM[10'hD6][17:13];	// lsu.scala:210:16
        ldq_12_bits_uop_edge_inst = _RANDOM[10'hD6][18];	// lsu.scala:210:16
        ldq_12_bits_uop_pc_lob = _RANDOM[10'hD6][24:19];	// lsu.scala:210:16
        ldq_12_bits_uop_taken = _RANDOM[10'hD6][25];	// lsu.scala:210:16
        ldq_12_bits_uop_imm_packed = {_RANDOM[10'hD6][31:26], _RANDOM[10'hD7][13:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_csr_addr = _RANDOM[10'hD7][25:14];	// lsu.scala:210:16
        ldq_12_bits_uop_rob_idx = {_RANDOM[10'hD7][31:26], _RANDOM[10'hD8][0]};	// lsu.scala:210:16
        ldq_12_bits_uop_ldq_idx = _RANDOM[10'hD8][5:1];	// lsu.scala:210:16
        ldq_12_bits_uop_stq_idx = _RANDOM[10'hD8][10:6];	// lsu.scala:210:16
        ldq_12_bits_uop_rxq_idx = _RANDOM[10'hD8][12:11];	// lsu.scala:210:16
        ldq_12_bits_uop_pdst = _RANDOM[10'hD8][19:13];	// lsu.scala:210:16
        ldq_12_bits_uop_prs1 = _RANDOM[10'hD8][26:20];	// lsu.scala:210:16
        ldq_12_bits_uop_prs2 = {_RANDOM[10'hD8][31:27], _RANDOM[10'hD9][1:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_prs3 = _RANDOM[10'hD9][8:2];	// lsu.scala:210:16
        ldq_12_bits_uop_ppred = _RANDOM[10'hD9][13:9];	// lsu.scala:210:16
        ldq_12_bits_uop_prs1_busy = _RANDOM[10'hD9][14];	// lsu.scala:210:16
        ldq_12_bits_uop_prs2_busy = _RANDOM[10'hD9][15];	// lsu.scala:210:16
        ldq_12_bits_uop_prs3_busy = _RANDOM[10'hD9][16];	// lsu.scala:210:16
        ldq_12_bits_uop_ppred_busy = _RANDOM[10'hD9][17];	// lsu.scala:210:16
        ldq_12_bits_uop_stale_pdst = _RANDOM[10'hD9][24:18];	// lsu.scala:210:16
        ldq_12_bits_uop_exception = _RANDOM[10'hD9][25];	// lsu.scala:210:16
        ldq_12_bits_uop_exc_cause =
          {_RANDOM[10'hD9][31:26], _RANDOM[10'hDA], _RANDOM[10'hDB][25:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_bypassable = _RANDOM[10'hDB][26];	// lsu.scala:210:16
        ldq_12_bits_uop_mem_cmd = _RANDOM[10'hDB][31:27];	// lsu.scala:210:16
        ldq_12_bits_uop_mem_size = _RANDOM[10'hDC][1:0];	// lsu.scala:210:16
        ldq_12_bits_uop_mem_signed = _RANDOM[10'hDC][2];	// lsu.scala:210:16
        ldq_12_bits_uop_is_fence = _RANDOM[10'hDC][3];	// lsu.scala:210:16
        ldq_12_bits_uop_is_fencei = _RANDOM[10'hDC][4];	// lsu.scala:210:16
        ldq_12_bits_uop_is_amo = _RANDOM[10'hDC][5];	// lsu.scala:210:16
        ldq_12_bits_uop_uses_ldq = _RANDOM[10'hDC][6];	// lsu.scala:210:16
        ldq_12_bits_uop_uses_stq = _RANDOM[10'hDC][7];	// lsu.scala:210:16
        ldq_12_bits_uop_is_sys_pc2epc = _RANDOM[10'hDC][8];	// lsu.scala:210:16
        ldq_12_bits_uop_is_unique = _RANDOM[10'hDC][9];	// lsu.scala:210:16
        ldq_12_bits_uop_flush_on_commit = _RANDOM[10'hDC][10];	// lsu.scala:210:16
        ldq_12_bits_uop_ldst_is_rs1 = _RANDOM[10'hDC][11];	// lsu.scala:210:16
        ldq_12_bits_uop_ldst = _RANDOM[10'hDC][17:12];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs1 = _RANDOM[10'hDC][23:18];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs2 = _RANDOM[10'hDC][29:24];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs3 = {_RANDOM[10'hDC][31:30], _RANDOM[10'hDD][3:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_ldst_val = _RANDOM[10'hDD][4];	// lsu.scala:210:16
        ldq_12_bits_uop_dst_rtype = _RANDOM[10'hDD][6:5];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs1_rtype = _RANDOM[10'hDD][8:7];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs2_rtype = _RANDOM[10'hDD][10:9];	// lsu.scala:210:16
        ldq_12_bits_uop_frs3_en = _RANDOM[10'hDD][11];	// lsu.scala:210:16
        ldq_12_bits_uop_fp_val = _RANDOM[10'hDD][12];	// lsu.scala:210:16
        ldq_12_bits_uop_fp_single = _RANDOM[10'hDD][13];	// lsu.scala:210:16
        ldq_12_bits_uop_xcpt_pf_if = _RANDOM[10'hDD][14];	// lsu.scala:210:16
        ldq_12_bits_uop_xcpt_ae_if = _RANDOM[10'hDD][15];	// lsu.scala:210:16
        ldq_12_bits_uop_xcpt_ma_if = _RANDOM[10'hDD][16];	// lsu.scala:210:16
        ldq_12_bits_uop_bp_debug_if = _RANDOM[10'hDD][17];	// lsu.scala:210:16
        ldq_12_bits_uop_bp_xcpt_if = _RANDOM[10'hDD][18];	// lsu.scala:210:16
        ldq_12_bits_uop_debug_fsrc = _RANDOM[10'hDD][20:19];	// lsu.scala:210:16
        ldq_12_bits_uop_debug_tsrc = _RANDOM[10'hDD][22:21];	// lsu.scala:210:16
        ldq_12_bits_addr_valid = _RANDOM[10'hDD][23];	// lsu.scala:210:16
        ldq_12_bits_addr_bits = {_RANDOM[10'hDD][31:24], _RANDOM[10'hDE]};	// lsu.scala:210:16
        ldq_12_bits_addr_is_virtual = _RANDOM[10'hDF][0];	// lsu.scala:210:16
        ldq_12_bits_addr_is_uncacheable = _RANDOM[10'hDF][1];	// lsu.scala:210:16
        ldq_12_bits_executed = _RANDOM[10'hDF][2];	// lsu.scala:210:16
        ldq_12_bits_succeeded = _RANDOM[10'hDF][3];	// lsu.scala:210:16
        ldq_12_bits_order_fail = _RANDOM[10'hDF][4];	// lsu.scala:210:16
        ldq_12_bits_observed = _RANDOM[10'hDF][5];	// lsu.scala:210:16
        ldq_12_bits_st_dep_mask = _RANDOM[10'hDF][29:6];	// lsu.scala:210:16
        ldq_12_bits_youngest_stq_idx = {_RANDOM[10'hDF][31:30], _RANDOM[10'hE0][2:0]};	// lsu.scala:210:16
        ldq_12_bits_forward_std_val = _RANDOM[10'hE0][3];	// lsu.scala:210:16
        ldq_12_bits_forward_stq_idx = _RANDOM[10'hE0][8:4];	// lsu.scala:210:16
        ldq_13_valid = _RANDOM[10'hE2][9];	// lsu.scala:210:16
        ldq_13_bits_uop_uopc = _RANDOM[10'hE2][16:10];	// lsu.scala:210:16
        ldq_13_bits_uop_inst = {_RANDOM[10'hE2][31:17], _RANDOM[10'hE3][16:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_debug_inst = {_RANDOM[10'hE3][31:17], _RANDOM[10'hE4][16:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_is_rvc = _RANDOM[10'hE4][17];	// lsu.scala:210:16
        ldq_13_bits_uop_debug_pc = {_RANDOM[10'hE4][31:18], _RANDOM[10'hE5][25:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_iq_type = _RANDOM[10'hE5][28:26];	// lsu.scala:210:16
        ldq_13_bits_uop_fu_code = {_RANDOM[10'hE5][31:29], _RANDOM[10'hE6][6:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_br_type = _RANDOM[10'hE6][10:7];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_op1_sel = _RANDOM[10'hE6][12:11];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_op2_sel = _RANDOM[10'hE6][15:13];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_imm_sel = _RANDOM[10'hE6][18:16];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_op_fcn = _RANDOM[10'hE6][22:19];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_fcn_dw = _RANDOM[10'hE6][23];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_csr_cmd = _RANDOM[10'hE6][26:24];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_is_load = _RANDOM[10'hE6][27];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_is_sta = _RANDOM[10'hE6][28];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_is_std = _RANDOM[10'hE6][29];	// lsu.scala:210:16
        ldq_13_bits_uop_iw_state = _RANDOM[10'hE6][31:30];	// lsu.scala:210:16
        ldq_13_bits_uop_iw_p1_poisoned = _RANDOM[10'hE7][0];	// lsu.scala:210:16
        ldq_13_bits_uop_iw_p2_poisoned = _RANDOM[10'hE7][1];	// lsu.scala:210:16
        ldq_13_bits_uop_is_br = _RANDOM[10'hE7][2];	// lsu.scala:210:16
        ldq_13_bits_uop_is_jalr = _RANDOM[10'hE7][3];	// lsu.scala:210:16
        ldq_13_bits_uop_is_jal = _RANDOM[10'hE7][4];	// lsu.scala:210:16
        ldq_13_bits_uop_is_sfb = _RANDOM[10'hE7][5];	// lsu.scala:210:16
        ldq_13_bits_uop_br_mask = _RANDOM[10'hE7][21:6];	// lsu.scala:210:16
        ldq_13_bits_uop_br_tag = _RANDOM[10'hE7][25:22];	// lsu.scala:210:16
        ldq_13_bits_uop_ftq_idx = _RANDOM[10'hE7][30:26];	// lsu.scala:210:16
        ldq_13_bits_uop_edge_inst = _RANDOM[10'hE7][31];	// lsu.scala:210:16
        ldq_13_bits_uop_pc_lob = _RANDOM[10'hE8][5:0];	// lsu.scala:210:16
        ldq_13_bits_uop_taken = _RANDOM[10'hE8][6];	// lsu.scala:210:16
        ldq_13_bits_uop_imm_packed = _RANDOM[10'hE8][26:7];	// lsu.scala:210:16
        ldq_13_bits_uop_csr_addr = {_RANDOM[10'hE8][31:27], _RANDOM[10'hE9][6:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_rob_idx = _RANDOM[10'hE9][13:7];	// lsu.scala:210:16
        ldq_13_bits_uop_ldq_idx = _RANDOM[10'hE9][18:14];	// lsu.scala:210:16
        ldq_13_bits_uop_stq_idx = _RANDOM[10'hE9][23:19];	// lsu.scala:210:16
        ldq_13_bits_uop_rxq_idx = _RANDOM[10'hE9][25:24];	// lsu.scala:210:16
        ldq_13_bits_uop_pdst = {_RANDOM[10'hE9][31:26], _RANDOM[10'hEA][0]};	// lsu.scala:210:16
        ldq_13_bits_uop_prs1 = _RANDOM[10'hEA][7:1];	// lsu.scala:210:16
        ldq_13_bits_uop_prs2 = _RANDOM[10'hEA][14:8];	// lsu.scala:210:16
        ldq_13_bits_uop_prs3 = _RANDOM[10'hEA][21:15];	// lsu.scala:210:16
        ldq_13_bits_uop_ppred = _RANDOM[10'hEA][26:22];	// lsu.scala:210:16
        ldq_13_bits_uop_prs1_busy = _RANDOM[10'hEA][27];	// lsu.scala:210:16
        ldq_13_bits_uop_prs2_busy = _RANDOM[10'hEA][28];	// lsu.scala:210:16
        ldq_13_bits_uop_prs3_busy = _RANDOM[10'hEA][29];	// lsu.scala:210:16
        ldq_13_bits_uop_ppred_busy = _RANDOM[10'hEA][30];	// lsu.scala:210:16
        ldq_13_bits_uop_stale_pdst = {_RANDOM[10'hEA][31], _RANDOM[10'hEB][5:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_exception = _RANDOM[10'hEB][6];	// lsu.scala:210:16
        ldq_13_bits_uop_exc_cause =
          {_RANDOM[10'hEB][31:7], _RANDOM[10'hEC], _RANDOM[10'hED][6:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_bypassable = _RANDOM[10'hED][7];	// lsu.scala:210:16
        ldq_13_bits_uop_mem_cmd = _RANDOM[10'hED][12:8];	// lsu.scala:210:16
        ldq_13_bits_uop_mem_size = _RANDOM[10'hED][14:13];	// lsu.scala:210:16
        ldq_13_bits_uop_mem_signed = _RANDOM[10'hED][15];	// lsu.scala:210:16
        ldq_13_bits_uop_is_fence = _RANDOM[10'hED][16];	// lsu.scala:210:16
        ldq_13_bits_uop_is_fencei = _RANDOM[10'hED][17];	// lsu.scala:210:16
        ldq_13_bits_uop_is_amo = _RANDOM[10'hED][18];	// lsu.scala:210:16
        ldq_13_bits_uop_uses_ldq = _RANDOM[10'hED][19];	// lsu.scala:210:16
        ldq_13_bits_uop_uses_stq = _RANDOM[10'hED][20];	// lsu.scala:210:16
        ldq_13_bits_uop_is_sys_pc2epc = _RANDOM[10'hED][21];	// lsu.scala:210:16
        ldq_13_bits_uop_is_unique = _RANDOM[10'hED][22];	// lsu.scala:210:16
        ldq_13_bits_uop_flush_on_commit = _RANDOM[10'hED][23];	// lsu.scala:210:16
        ldq_13_bits_uop_ldst_is_rs1 = _RANDOM[10'hED][24];	// lsu.scala:210:16
        ldq_13_bits_uop_ldst = _RANDOM[10'hED][30:25];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs1 = {_RANDOM[10'hED][31], _RANDOM[10'hEE][4:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_lrs2 = _RANDOM[10'hEE][10:5];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs3 = _RANDOM[10'hEE][16:11];	// lsu.scala:210:16
        ldq_13_bits_uop_ldst_val = _RANDOM[10'hEE][17];	// lsu.scala:210:16
        ldq_13_bits_uop_dst_rtype = _RANDOM[10'hEE][19:18];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs1_rtype = _RANDOM[10'hEE][21:20];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs2_rtype = _RANDOM[10'hEE][23:22];	// lsu.scala:210:16
        ldq_13_bits_uop_frs3_en = _RANDOM[10'hEE][24];	// lsu.scala:210:16
        ldq_13_bits_uop_fp_val = _RANDOM[10'hEE][25];	// lsu.scala:210:16
        ldq_13_bits_uop_fp_single = _RANDOM[10'hEE][26];	// lsu.scala:210:16
        ldq_13_bits_uop_xcpt_pf_if = _RANDOM[10'hEE][27];	// lsu.scala:210:16
        ldq_13_bits_uop_xcpt_ae_if = _RANDOM[10'hEE][28];	// lsu.scala:210:16
        ldq_13_bits_uop_xcpt_ma_if = _RANDOM[10'hEE][29];	// lsu.scala:210:16
        ldq_13_bits_uop_bp_debug_if = _RANDOM[10'hEE][30];	// lsu.scala:210:16
        ldq_13_bits_uop_bp_xcpt_if = _RANDOM[10'hEE][31];	// lsu.scala:210:16
        ldq_13_bits_uop_debug_fsrc = _RANDOM[10'hEF][1:0];	// lsu.scala:210:16
        ldq_13_bits_uop_debug_tsrc = _RANDOM[10'hEF][3:2];	// lsu.scala:210:16
        ldq_13_bits_addr_valid = _RANDOM[10'hEF][4];	// lsu.scala:210:16
        ldq_13_bits_addr_bits = {_RANDOM[10'hEF][31:5], _RANDOM[10'hF0][12:0]};	// lsu.scala:210:16
        ldq_13_bits_addr_is_virtual = _RANDOM[10'hF0][13];	// lsu.scala:210:16
        ldq_13_bits_addr_is_uncacheable = _RANDOM[10'hF0][14];	// lsu.scala:210:16
        ldq_13_bits_executed = _RANDOM[10'hF0][15];	// lsu.scala:210:16
        ldq_13_bits_succeeded = _RANDOM[10'hF0][16];	// lsu.scala:210:16
        ldq_13_bits_order_fail = _RANDOM[10'hF0][17];	// lsu.scala:210:16
        ldq_13_bits_observed = _RANDOM[10'hF0][18];	// lsu.scala:210:16
        ldq_13_bits_st_dep_mask = {_RANDOM[10'hF0][31:19], _RANDOM[10'hF1][10:0]};	// lsu.scala:210:16
        ldq_13_bits_youngest_stq_idx = _RANDOM[10'hF1][15:11];	// lsu.scala:210:16
        ldq_13_bits_forward_std_val = _RANDOM[10'hF1][16];	// lsu.scala:210:16
        ldq_13_bits_forward_stq_idx = _RANDOM[10'hF1][21:17];	// lsu.scala:210:16
        ldq_14_valid = _RANDOM[10'hF3][22];	// lsu.scala:210:16
        ldq_14_bits_uop_uopc = _RANDOM[10'hF3][29:23];	// lsu.scala:210:16
        ldq_14_bits_uop_inst = {_RANDOM[10'hF3][31:30], _RANDOM[10'hF4][29:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_debug_inst = {_RANDOM[10'hF4][31:30], _RANDOM[10'hF5][29:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_is_rvc = _RANDOM[10'hF5][30];	// lsu.scala:210:16
        ldq_14_bits_uop_debug_pc =
          {_RANDOM[10'hF5][31], _RANDOM[10'hF6], _RANDOM[10'hF7][6:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_iq_type = _RANDOM[10'hF7][9:7];	// lsu.scala:210:16
        ldq_14_bits_uop_fu_code = _RANDOM[10'hF7][19:10];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_br_type = _RANDOM[10'hF7][23:20];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_op1_sel = _RANDOM[10'hF7][25:24];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_op2_sel = _RANDOM[10'hF7][28:26];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_imm_sel = _RANDOM[10'hF7][31:29];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_op_fcn = _RANDOM[10'hF8][3:0];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_fcn_dw = _RANDOM[10'hF8][4];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_csr_cmd = _RANDOM[10'hF8][7:5];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_is_load = _RANDOM[10'hF8][8];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_is_sta = _RANDOM[10'hF8][9];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_is_std = _RANDOM[10'hF8][10];	// lsu.scala:210:16
        ldq_14_bits_uop_iw_state = _RANDOM[10'hF8][12:11];	// lsu.scala:210:16
        ldq_14_bits_uop_iw_p1_poisoned = _RANDOM[10'hF8][13];	// lsu.scala:210:16
        ldq_14_bits_uop_iw_p2_poisoned = _RANDOM[10'hF8][14];	// lsu.scala:210:16
        ldq_14_bits_uop_is_br = _RANDOM[10'hF8][15];	// lsu.scala:210:16
        ldq_14_bits_uop_is_jalr = _RANDOM[10'hF8][16];	// lsu.scala:210:16
        ldq_14_bits_uop_is_jal = _RANDOM[10'hF8][17];	// lsu.scala:210:16
        ldq_14_bits_uop_is_sfb = _RANDOM[10'hF8][18];	// lsu.scala:210:16
        ldq_14_bits_uop_br_mask = {_RANDOM[10'hF8][31:19], _RANDOM[10'hF9][2:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_br_tag = _RANDOM[10'hF9][6:3];	// lsu.scala:210:16
        ldq_14_bits_uop_ftq_idx = _RANDOM[10'hF9][11:7];	// lsu.scala:210:16
        ldq_14_bits_uop_edge_inst = _RANDOM[10'hF9][12];	// lsu.scala:210:16
        ldq_14_bits_uop_pc_lob = _RANDOM[10'hF9][18:13];	// lsu.scala:210:16
        ldq_14_bits_uop_taken = _RANDOM[10'hF9][19];	// lsu.scala:210:16
        ldq_14_bits_uop_imm_packed = {_RANDOM[10'hF9][31:20], _RANDOM[10'hFA][7:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_csr_addr = _RANDOM[10'hFA][19:8];	// lsu.scala:210:16
        ldq_14_bits_uop_rob_idx = _RANDOM[10'hFA][26:20];	// lsu.scala:210:16
        ldq_14_bits_uop_ldq_idx = _RANDOM[10'hFA][31:27];	// lsu.scala:210:16
        ldq_14_bits_uop_stq_idx = _RANDOM[10'hFB][4:0];	// lsu.scala:210:16
        ldq_14_bits_uop_rxq_idx = _RANDOM[10'hFB][6:5];	// lsu.scala:210:16
        ldq_14_bits_uop_pdst = _RANDOM[10'hFB][13:7];	// lsu.scala:210:16
        ldq_14_bits_uop_prs1 = _RANDOM[10'hFB][20:14];	// lsu.scala:210:16
        ldq_14_bits_uop_prs2 = _RANDOM[10'hFB][27:21];	// lsu.scala:210:16
        ldq_14_bits_uop_prs3 = {_RANDOM[10'hFB][31:28], _RANDOM[10'hFC][2:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_ppred = _RANDOM[10'hFC][7:3];	// lsu.scala:210:16
        ldq_14_bits_uop_prs1_busy = _RANDOM[10'hFC][8];	// lsu.scala:210:16
        ldq_14_bits_uop_prs2_busy = _RANDOM[10'hFC][9];	// lsu.scala:210:16
        ldq_14_bits_uop_prs3_busy = _RANDOM[10'hFC][10];	// lsu.scala:210:16
        ldq_14_bits_uop_ppred_busy = _RANDOM[10'hFC][11];	// lsu.scala:210:16
        ldq_14_bits_uop_stale_pdst = _RANDOM[10'hFC][18:12];	// lsu.scala:210:16
        ldq_14_bits_uop_exception = _RANDOM[10'hFC][19];	// lsu.scala:210:16
        ldq_14_bits_uop_exc_cause =
          {_RANDOM[10'hFC][31:20], _RANDOM[10'hFD], _RANDOM[10'hFE][19:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_bypassable = _RANDOM[10'hFE][20];	// lsu.scala:210:16
        ldq_14_bits_uop_mem_cmd = _RANDOM[10'hFE][25:21];	// lsu.scala:210:16
        ldq_14_bits_uop_mem_size = _RANDOM[10'hFE][27:26];	// lsu.scala:210:16
        ldq_14_bits_uop_mem_signed = _RANDOM[10'hFE][28];	// lsu.scala:210:16
        ldq_14_bits_uop_is_fence = _RANDOM[10'hFE][29];	// lsu.scala:210:16
        ldq_14_bits_uop_is_fencei = _RANDOM[10'hFE][30];	// lsu.scala:210:16
        ldq_14_bits_uop_is_amo = _RANDOM[10'hFE][31];	// lsu.scala:210:16
        ldq_14_bits_uop_uses_ldq = _RANDOM[10'hFF][0];	// lsu.scala:210:16
        ldq_14_bits_uop_uses_stq = _RANDOM[10'hFF][1];	// lsu.scala:210:16
        ldq_14_bits_uop_is_sys_pc2epc = _RANDOM[10'hFF][2];	// lsu.scala:210:16
        ldq_14_bits_uop_is_unique = _RANDOM[10'hFF][3];	// lsu.scala:210:16
        ldq_14_bits_uop_flush_on_commit = _RANDOM[10'hFF][4];	// lsu.scala:210:16
        ldq_14_bits_uop_ldst_is_rs1 = _RANDOM[10'hFF][5];	// lsu.scala:210:16
        ldq_14_bits_uop_ldst = _RANDOM[10'hFF][11:6];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs1 = _RANDOM[10'hFF][17:12];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs2 = _RANDOM[10'hFF][23:18];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs3 = _RANDOM[10'hFF][29:24];	// lsu.scala:210:16
        ldq_14_bits_uop_ldst_val = _RANDOM[10'hFF][30];	// lsu.scala:210:16
        ldq_14_bits_uop_dst_rtype = {_RANDOM[10'hFF][31], _RANDOM[10'h100][0]};	// lsu.scala:210:16
        ldq_14_bits_uop_lrs1_rtype = _RANDOM[10'h100][2:1];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs2_rtype = _RANDOM[10'h100][4:3];	// lsu.scala:210:16
        ldq_14_bits_uop_frs3_en = _RANDOM[10'h100][5];	// lsu.scala:210:16
        ldq_14_bits_uop_fp_val = _RANDOM[10'h100][6];	// lsu.scala:210:16
        ldq_14_bits_uop_fp_single = _RANDOM[10'h100][7];	// lsu.scala:210:16
        ldq_14_bits_uop_xcpt_pf_if = _RANDOM[10'h100][8];	// lsu.scala:210:16
        ldq_14_bits_uop_xcpt_ae_if = _RANDOM[10'h100][9];	// lsu.scala:210:16
        ldq_14_bits_uop_xcpt_ma_if = _RANDOM[10'h100][10];	// lsu.scala:210:16
        ldq_14_bits_uop_bp_debug_if = _RANDOM[10'h100][11];	// lsu.scala:210:16
        ldq_14_bits_uop_bp_xcpt_if = _RANDOM[10'h100][12];	// lsu.scala:210:16
        ldq_14_bits_uop_debug_fsrc = _RANDOM[10'h100][14:13];	// lsu.scala:210:16
        ldq_14_bits_uop_debug_tsrc = _RANDOM[10'h100][16:15];	// lsu.scala:210:16
        ldq_14_bits_addr_valid = _RANDOM[10'h100][17];	// lsu.scala:210:16
        ldq_14_bits_addr_bits = {_RANDOM[10'h100][31:18], _RANDOM[10'h101][25:0]};	// lsu.scala:210:16
        ldq_14_bits_addr_is_virtual = _RANDOM[10'h101][26];	// lsu.scala:210:16
        ldq_14_bits_addr_is_uncacheable = _RANDOM[10'h101][27];	// lsu.scala:210:16
        ldq_14_bits_executed = _RANDOM[10'h101][28];	// lsu.scala:210:16
        ldq_14_bits_succeeded = _RANDOM[10'h101][29];	// lsu.scala:210:16
        ldq_14_bits_order_fail = _RANDOM[10'h101][30];	// lsu.scala:210:16
        ldq_14_bits_observed = _RANDOM[10'h101][31];	// lsu.scala:210:16
        ldq_14_bits_st_dep_mask = _RANDOM[10'h102][23:0];	// lsu.scala:210:16
        ldq_14_bits_youngest_stq_idx = _RANDOM[10'h102][28:24];	// lsu.scala:210:16
        ldq_14_bits_forward_std_val = _RANDOM[10'h102][29];	// lsu.scala:210:16
        ldq_14_bits_forward_stq_idx = {_RANDOM[10'h102][31:30], _RANDOM[10'h103][2:0]};	// lsu.scala:210:16
        ldq_15_valid = _RANDOM[10'h105][3];	// lsu.scala:210:16
        ldq_15_bits_uop_uopc = _RANDOM[10'h105][10:4];	// lsu.scala:210:16
        ldq_15_bits_uop_inst = {_RANDOM[10'h105][31:11], _RANDOM[10'h106][10:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_debug_inst = {_RANDOM[10'h106][31:11], _RANDOM[10'h107][10:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_is_rvc = _RANDOM[10'h107][11];	// lsu.scala:210:16
        ldq_15_bits_uop_debug_pc = {_RANDOM[10'h107][31:12], _RANDOM[10'h108][19:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_iq_type = _RANDOM[10'h108][22:20];	// lsu.scala:210:16
        ldq_15_bits_uop_fu_code = {_RANDOM[10'h108][31:23], _RANDOM[10'h109][0]};	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_br_type = _RANDOM[10'h109][4:1];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_op1_sel = _RANDOM[10'h109][6:5];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_op2_sel = _RANDOM[10'h109][9:7];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_imm_sel = _RANDOM[10'h109][12:10];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_op_fcn = _RANDOM[10'h109][16:13];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_fcn_dw = _RANDOM[10'h109][17];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_csr_cmd = _RANDOM[10'h109][20:18];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_is_load = _RANDOM[10'h109][21];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_is_sta = _RANDOM[10'h109][22];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_is_std = _RANDOM[10'h109][23];	// lsu.scala:210:16
        ldq_15_bits_uop_iw_state = _RANDOM[10'h109][25:24];	// lsu.scala:210:16
        ldq_15_bits_uop_iw_p1_poisoned = _RANDOM[10'h109][26];	// lsu.scala:210:16
        ldq_15_bits_uop_iw_p2_poisoned = _RANDOM[10'h109][27];	// lsu.scala:210:16
        ldq_15_bits_uop_is_br = _RANDOM[10'h109][28];	// lsu.scala:210:16
        ldq_15_bits_uop_is_jalr = _RANDOM[10'h109][29];	// lsu.scala:210:16
        ldq_15_bits_uop_is_jal = _RANDOM[10'h109][30];	// lsu.scala:210:16
        ldq_15_bits_uop_is_sfb = _RANDOM[10'h109][31];	// lsu.scala:210:16
        ldq_15_bits_uop_br_mask = _RANDOM[10'h10A][15:0];	// lsu.scala:210:16
        ldq_15_bits_uop_br_tag = _RANDOM[10'h10A][19:16];	// lsu.scala:210:16
        ldq_15_bits_uop_ftq_idx = _RANDOM[10'h10A][24:20];	// lsu.scala:210:16
        ldq_15_bits_uop_edge_inst = _RANDOM[10'h10A][25];	// lsu.scala:210:16
        ldq_15_bits_uop_pc_lob = _RANDOM[10'h10A][31:26];	// lsu.scala:210:16
        ldq_15_bits_uop_taken = _RANDOM[10'h10B][0];	// lsu.scala:210:16
        ldq_15_bits_uop_imm_packed = _RANDOM[10'h10B][20:1];	// lsu.scala:210:16
        ldq_15_bits_uop_csr_addr = {_RANDOM[10'h10B][31:21], _RANDOM[10'h10C][0]};	// lsu.scala:210:16
        ldq_15_bits_uop_rob_idx = _RANDOM[10'h10C][7:1];	// lsu.scala:210:16
        ldq_15_bits_uop_ldq_idx = _RANDOM[10'h10C][12:8];	// lsu.scala:210:16
        ldq_15_bits_uop_stq_idx = _RANDOM[10'h10C][17:13];	// lsu.scala:210:16
        ldq_15_bits_uop_rxq_idx = _RANDOM[10'h10C][19:18];	// lsu.scala:210:16
        ldq_15_bits_uop_pdst = _RANDOM[10'h10C][26:20];	// lsu.scala:210:16
        ldq_15_bits_uop_prs1 = {_RANDOM[10'h10C][31:27], _RANDOM[10'h10D][1:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_prs2 = _RANDOM[10'h10D][8:2];	// lsu.scala:210:16
        ldq_15_bits_uop_prs3 = _RANDOM[10'h10D][15:9];	// lsu.scala:210:16
        ldq_15_bits_uop_ppred = _RANDOM[10'h10D][20:16];	// lsu.scala:210:16
        ldq_15_bits_uop_prs1_busy = _RANDOM[10'h10D][21];	// lsu.scala:210:16
        ldq_15_bits_uop_prs2_busy = _RANDOM[10'h10D][22];	// lsu.scala:210:16
        ldq_15_bits_uop_prs3_busy = _RANDOM[10'h10D][23];	// lsu.scala:210:16
        ldq_15_bits_uop_ppred_busy = _RANDOM[10'h10D][24];	// lsu.scala:210:16
        ldq_15_bits_uop_stale_pdst = _RANDOM[10'h10D][31:25];	// lsu.scala:210:16
        ldq_15_bits_uop_exception = _RANDOM[10'h10E][0];	// lsu.scala:210:16
        ldq_15_bits_uop_exc_cause =
          {_RANDOM[10'h10E][31:1], _RANDOM[10'h10F], _RANDOM[10'h110][0]};	// lsu.scala:210:16
        ldq_15_bits_uop_bypassable = _RANDOM[10'h110][1];	// lsu.scala:210:16
        ldq_15_bits_uop_mem_cmd = _RANDOM[10'h110][6:2];	// lsu.scala:210:16
        ldq_15_bits_uop_mem_size = _RANDOM[10'h110][8:7];	// lsu.scala:210:16
        ldq_15_bits_uop_mem_signed = _RANDOM[10'h110][9];	// lsu.scala:210:16
        ldq_15_bits_uop_is_fence = _RANDOM[10'h110][10];	// lsu.scala:210:16
        ldq_15_bits_uop_is_fencei = _RANDOM[10'h110][11];	// lsu.scala:210:16
        ldq_15_bits_uop_is_amo = _RANDOM[10'h110][12];	// lsu.scala:210:16
        ldq_15_bits_uop_uses_ldq = _RANDOM[10'h110][13];	// lsu.scala:210:16
        ldq_15_bits_uop_uses_stq = _RANDOM[10'h110][14];	// lsu.scala:210:16
        ldq_15_bits_uop_is_sys_pc2epc = _RANDOM[10'h110][15];	// lsu.scala:210:16
        ldq_15_bits_uop_is_unique = _RANDOM[10'h110][16];	// lsu.scala:210:16
        ldq_15_bits_uop_flush_on_commit = _RANDOM[10'h110][17];	// lsu.scala:210:16
        ldq_15_bits_uop_ldst_is_rs1 = _RANDOM[10'h110][18];	// lsu.scala:210:16
        ldq_15_bits_uop_ldst = _RANDOM[10'h110][24:19];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs1 = _RANDOM[10'h110][30:25];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs2 = {_RANDOM[10'h110][31], _RANDOM[10'h111][4:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_lrs3 = _RANDOM[10'h111][10:5];	// lsu.scala:210:16
        ldq_15_bits_uop_ldst_val = _RANDOM[10'h111][11];	// lsu.scala:210:16
        ldq_15_bits_uop_dst_rtype = _RANDOM[10'h111][13:12];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs1_rtype = _RANDOM[10'h111][15:14];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs2_rtype = _RANDOM[10'h111][17:16];	// lsu.scala:210:16
        ldq_15_bits_uop_frs3_en = _RANDOM[10'h111][18];	// lsu.scala:210:16
        ldq_15_bits_uop_fp_val = _RANDOM[10'h111][19];	// lsu.scala:210:16
        ldq_15_bits_uop_fp_single = _RANDOM[10'h111][20];	// lsu.scala:210:16
        ldq_15_bits_uop_xcpt_pf_if = _RANDOM[10'h111][21];	// lsu.scala:210:16
        ldq_15_bits_uop_xcpt_ae_if = _RANDOM[10'h111][22];	// lsu.scala:210:16
        ldq_15_bits_uop_xcpt_ma_if = _RANDOM[10'h111][23];	// lsu.scala:210:16
        ldq_15_bits_uop_bp_debug_if = _RANDOM[10'h111][24];	// lsu.scala:210:16
        ldq_15_bits_uop_bp_xcpt_if = _RANDOM[10'h111][25];	// lsu.scala:210:16
        ldq_15_bits_uop_debug_fsrc = _RANDOM[10'h111][27:26];	// lsu.scala:210:16
        ldq_15_bits_uop_debug_tsrc = _RANDOM[10'h111][29:28];	// lsu.scala:210:16
        ldq_15_bits_addr_valid = _RANDOM[10'h111][30];	// lsu.scala:210:16
        ldq_15_bits_addr_bits =
          {_RANDOM[10'h111][31], _RANDOM[10'h112], _RANDOM[10'h113][6:0]};	// lsu.scala:210:16
        ldq_15_bits_addr_is_virtual = _RANDOM[10'h113][7];	// lsu.scala:210:16
        ldq_15_bits_addr_is_uncacheable = _RANDOM[10'h113][8];	// lsu.scala:210:16
        ldq_15_bits_executed = _RANDOM[10'h113][9];	// lsu.scala:210:16
        ldq_15_bits_succeeded = _RANDOM[10'h113][10];	// lsu.scala:210:16
        ldq_15_bits_order_fail = _RANDOM[10'h113][11];	// lsu.scala:210:16
        ldq_15_bits_observed = _RANDOM[10'h113][12];	// lsu.scala:210:16
        ldq_15_bits_st_dep_mask = {_RANDOM[10'h113][31:13], _RANDOM[10'h114][4:0]};	// lsu.scala:210:16
        ldq_15_bits_youngest_stq_idx = _RANDOM[10'h114][9:5];	// lsu.scala:210:16
        ldq_15_bits_forward_std_val = _RANDOM[10'h114][10];	// lsu.scala:210:16
        ldq_15_bits_forward_stq_idx = _RANDOM[10'h114][15:11];	// lsu.scala:210:16
        ldq_16_valid = _RANDOM[10'h116][16];	// lsu.scala:210:16
        ldq_16_bits_uop_uopc = _RANDOM[10'h116][23:17];	// lsu.scala:210:16
        ldq_16_bits_uop_inst = {_RANDOM[10'h116][31:24], _RANDOM[10'h117][23:0]};	// lsu.scala:210:16
        ldq_16_bits_uop_debug_inst = {_RANDOM[10'h117][31:24], _RANDOM[10'h118][23:0]};	// lsu.scala:210:16
        ldq_16_bits_uop_is_rvc = _RANDOM[10'h118][24];	// lsu.scala:210:16
        ldq_16_bits_uop_debug_pc =
          {_RANDOM[10'h118][31:25], _RANDOM[10'h119], _RANDOM[10'h11A][0]};	// lsu.scala:210:16
        ldq_16_bits_uop_iq_type = _RANDOM[10'h11A][3:1];	// lsu.scala:210:16
        ldq_16_bits_uop_fu_code = _RANDOM[10'h11A][13:4];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_br_type = _RANDOM[10'h11A][17:14];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_op1_sel = _RANDOM[10'h11A][19:18];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_op2_sel = _RANDOM[10'h11A][22:20];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_imm_sel = _RANDOM[10'h11A][25:23];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_op_fcn = _RANDOM[10'h11A][29:26];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_fcn_dw = _RANDOM[10'h11A][30];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h11A][31], _RANDOM[10'h11B][1:0]};	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_is_load = _RANDOM[10'h11B][2];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_is_sta = _RANDOM[10'h11B][3];	// lsu.scala:210:16
        ldq_16_bits_uop_ctrl_is_std = _RANDOM[10'h11B][4];	// lsu.scala:210:16
        ldq_16_bits_uop_iw_state = _RANDOM[10'h11B][6:5];	// lsu.scala:210:16
        ldq_16_bits_uop_iw_p1_poisoned = _RANDOM[10'h11B][7];	// lsu.scala:210:16
        ldq_16_bits_uop_iw_p2_poisoned = _RANDOM[10'h11B][8];	// lsu.scala:210:16
        ldq_16_bits_uop_is_br = _RANDOM[10'h11B][9];	// lsu.scala:210:16
        ldq_16_bits_uop_is_jalr = _RANDOM[10'h11B][10];	// lsu.scala:210:16
        ldq_16_bits_uop_is_jal = _RANDOM[10'h11B][11];	// lsu.scala:210:16
        ldq_16_bits_uop_is_sfb = _RANDOM[10'h11B][12];	// lsu.scala:210:16
        ldq_16_bits_uop_br_mask = _RANDOM[10'h11B][28:13];	// lsu.scala:210:16
        ldq_16_bits_uop_br_tag = {_RANDOM[10'h11B][31:29], _RANDOM[10'h11C][0]};	// lsu.scala:210:16
        ldq_16_bits_uop_ftq_idx = _RANDOM[10'h11C][5:1];	// lsu.scala:210:16
        ldq_16_bits_uop_edge_inst = _RANDOM[10'h11C][6];	// lsu.scala:210:16
        ldq_16_bits_uop_pc_lob = _RANDOM[10'h11C][12:7];	// lsu.scala:210:16
        ldq_16_bits_uop_taken = _RANDOM[10'h11C][13];	// lsu.scala:210:16
        ldq_16_bits_uop_imm_packed = {_RANDOM[10'h11C][31:14], _RANDOM[10'h11D][1:0]};	// lsu.scala:210:16
        ldq_16_bits_uop_csr_addr = _RANDOM[10'h11D][13:2];	// lsu.scala:210:16
        ldq_16_bits_uop_rob_idx = _RANDOM[10'h11D][20:14];	// lsu.scala:210:16
        ldq_16_bits_uop_ldq_idx = _RANDOM[10'h11D][25:21];	// lsu.scala:210:16
        ldq_16_bits_uop_stq_idx = _RANDOM[10'h11D][30:26];	// lsu.scala:210:16
        ldq_16_bits_uop_rxq_idx = {_RANDOM[10'h11D][31], _RANDOM[10'h11E][0]};	// lsu.scala:210:16
        ldq_16_bits_uop_pdst = _RANDOM[10'h11E][7:1];	// lsu.scala:210:16
        ldq_16_bits_uop_prs1 = _RANDOM[10'h11E][14:8];	// lsu.scala:210:16
        ldq_16_bits_uop_prs2 = _RANDOM[10'h11E][21:15];	// lsu.scala:210:16
        ldq_16_bits_uop_prs3 = _RANDOM[10'h11E][28:22];	// lsu.scala:210:16
        ldq_16_bits_uop_ppred = {_RANDOM[10'h11E][31:29], _RANDOM[10'h11F][1:0]};	// lsu.scala:210:16
        ldq_16_bits_uop_prs1_busy = _RANDOM[10'h11F][2];	// lsu.scala:210:16
        ldq_16_bits_uop_prs2_busy = _RANDOM[10'h11F][3];	// lsu.scala:210:16
        ldq_16_bits_uop_prs3_busy = _RANDOM[10'h11F][4];	// lsu.scala:210:16
        ldq_16_bits_uop_ppred_busy = _RANDOM[10'h11F][5];	// lsu.scala:210:16
        ldq_16_bits_uop_stale_pdst = _RANDOM[10'h11F][12:6];	// lsu.scala:210:16
        ldq_16_bits_uop_exception = _RANDOM[10'h11F][13];	// lsu.scala:210:16
        ldq_16_bits_uop_exc_cause =
          {_RANDOM[10'h11F][31:14], _RANDOM[10'h120], _RANDOM[10'h121][13:0]};	// lsu.scala:210:16
        ldq_16_bits_uop_bypassable = _RANDOM[10'h121][14];	// lsu.scala:210:16
        ldq_16_bits_uop_mem_cmd = _RANDOM[10'h121][19:15];	// lsu.scala:210:16
        ldq_16_bits_uop_mem_size = _RANDOM[10'h121][21:20];	// lsu.scala:210:16
        ldq_16_bits_uop_mem_signed = _RANDOM[10'h121][22];	// lsu.scala:210:16
        ldq_16_bits_uop_is_fence = _RANDOM[10'h121][23];	// lsu.scala:210:16
        ldq_16_bits_uop_is_fencei = _RANDOM[10'h121][24];	// lsu.scala:210:16
        ldq_16_bits_uop_is_amo = _RANDOM[10'h121][25];	// lsu.scala:210:16
        ldq_16_bits_uop_uses_ldq = _RANDOM[10'h121][26];	// lsu.scala:210:16
        ldq_16_bits_uop_uses_stq = _RANDOM[10'h121][27];	// lsu.scala:210:16
        ldq_16_bits_uop_is_sys_pc2epc = _RANDOM[10'h121][28];	// lsu.scala:210:16
        ldq_16_bits_uop_is_unique = _RANDOM[10'h121][29];	// lsu.scala:210:16
        ldq_16_bits_uop_flush_on_commit = _RANDOM[10'h121][30];	// lsu.scala:210:16
        ldq_16_bits_uop_ldst_is_rs1 = _RANDOM[10'h121][31];	// lsu.scala:210:16
        ldq_16_bits_uop_ldst = _RANDOM[10'h122][5:0];	// lsu.scala:210:16
        ldq_16_bits_uop_lrs1 = _RANDOM[10'h122][11:6];	// lsu.scala:210:16
        ldq_16_bits_uop_lrs2 = _RANDOM[10'h122][17:12];	// lsu.scala:210:16
        ldq_16_bits_uop_lrs3 = _RANDOM[10'h122][23:18];	// lsu.scala:210:16
        ldq_16_bits_uop_ldst_val = _RANDOM[10'h122][24];	// lsu.scala:210:16
        ldq_16_bits_uop_dst_rtype = _RANDOM[10'h122][26:25];	// lsu.scala:210:16
        ldq_16_bits_uop_lrs1_rtype = _RANDOM[10'h122][28:27];	// lsu.scala:210:16
        ldq_16_bits_uop_lrs2_rtype = _RANDOM[10'h122][30:29];	// lsu.scala:210:16
        ldq_16_bits_uop_frs3_en = _RANDOM[10'h122][31];	// lsu.scala:210:16
        ldq_16_bits_uop_fp_val = _RANDOM[10'h123][0];	// lsu.scala:210:16
        ldq_16_bits_uop_fp_single = _RANDOM[10'h123][1];	// lsu.scala:210:16
        ldq_16_bits_uop_xcpt_pf_if = _RANDOM[10'h123][2];	// lsu.scala:210:16
        ldq_16_bits_uop_xcpt_ae_if = _RANDOM[10'h123][3];	// lsu.scala:210:16
        ldq_16_bits_uop_xcpt_ma_if = _RANDOM[10'h123][4];	// lsu.scala:210:16
        ldq_16_bits_uop_bp_debug_if = _RANDOM[10'h123][5];	// lsu.scala:210:16
        ldq_16_bits_uop_bp_xcpt_if = _RANDOM[10'h123][6];	// lsu.scala:210:16
        ldq_16_bits_uop_debug_fsrc = _RANDOM[10'h123][8:7];	// lsu.scala:210:16
        ldq_16_bits_uop_debug_tsrc = _RANDOM[10'h123][10:9];	// lsu.scala:210:16
        ldq_16_bits_addr_valid = _RANDOM[10'h123][11];	// lsu.scala:210:16
        ldq_16_bits_addr_bits = {_RANDOM[10'h123][31:12], _RANDOM[10'h124][19:0]};	// lsu.scala:210:16
        ldq_16_bits_addr_is_virtual = _RANDOM[10'h124][20];	// lsu.scala:210:16
        ldq_16_bits_addr_is_uncacheable = _RANDOM[10'h124][21];	// lsu.scala:210:16
        ldq_16_bits_executed = _RANDOM[10'h124][22];	// lsu.scala:210:16
        ldq_16_bits_succeeded = _RANDOM[10'h124][23];	// lsu.scala:210:16
        ldq_16_bits_order_fail = _RANDOM[10'h124][24];	// lsu.scala:210:16
        ldq_16_bits_observed = _RANDOM[10'h124][25];	// lsu.scala:210:16
        ldq_16_bits_st_dep_mask = {_RANDOM[10'h124][31:26], _RANDOM[10'h125][17:0]};	// lsu.scala:210:16
        ldq_16_bits_youngest_stq_idx = _RANDOM[10'h125][22:18];	// lsu.scala:210:16
        ldq_16_bits_forward_std_val = _RANDOM[10'h125][23];	// lsu.scala:210:16
        ldq_16_bits_forward_stq_idx = _RANDOM[10'h125][28:24];	// lsu.scala:210:16
        ldq_17_valid = _RANDOM[10'h127][29];	// lsu.scala:210:16
        ldq_17_bits_uop_uopc = {_RANDOM[10'h127][31:30], _RANDOM[10'h128][4:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_inst = {_RANDOM[10'h128][31:5], _RANDOM[10'h129][4:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_debug_inst = {_RANDOM[10'h129][31:5], _RANDOM[10'h12A][4:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_is_rvc = _RANDOM[10'h12A][5];	// lsu.scala:210:16
        ldq_17_bits_uop_debug_pc = {_RANDOM[10'h12A][31:6], _RANDOM[10'h12B][13:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_iq_type = _RANDOM[10'h12B][16:14];	// lsu.scala:210:16
        ldq_17_bits_uop_fu_code = _RANDOM[10'h12B][26:17];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_br_type = _RANDOM[10'h12B][30:27];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_op1_sel = {_RANDOM[10'h12B][31], _RANDOM[10'h12C][0]};	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_op2_sel = _RANDOM[10'h12C][3:1];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_imm_sel = _RANDOM[10'h12C][6:4];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_op_fcn = _RANDOM[10'h12C][10:7];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_fcn_dw = _RANDOM[10'h12C][11];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_csr_cmd = _RANDOM[10'h12C][14:12];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_is_load = _RANDOM[10'h12C][15];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_is_sta = _RANDOM[10'h12C][16];	// lsu.scala:210:16
        ldq_17_bits_uop_ctrl_is_std = _RANDOM[10'h12C][17];	// lsu.scala:210:16
        ldq_17_bits_uop_iw_state = _RANDOM[10'h12C][19:18];	// lsu.scala:210:16
        ldq_17_bits_uop_iw_p1_poisoned = _RANDOM[10'h12C][20];	// lsu.scala:210:16
        ldq_17_bits_uop_iw_p2_poisoned = _RANDOM[10'h12C][21];	// lsu.scala:210:16
        ldq_17_bits_uop_is_br = _RANDOM[10'h12C][22];	// lsu.scala:210:16
        ldq_17_bits_uop_is_jalr = _RANDOM[10'h12C][23];	// lsu.scala:210:16
        ldq_17_bits_uop_is_jal = _RANDOM[10'h12C][24];	// lsu.scala:210:16
        ldq_17_bits_uop_is_sfb = _RANDOM[10'h12C][25];	// lsu.scala:210:16
        ldq_17_bits_uop_br_mask = {_RANDOM[10'h12C][31:26], _RANDOM[10'h12D][9:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_br_tag = _RANDOM[10'h12D][13:10];	// lsu.scala:210:16
        ldq_17_bits_uop_ftq_idx = _RANDOM[10'h12D][18:14];	// lsu.scala:210:16
        ldq_17_bits_uop_edge_inst = _RANDOM[10'h12D][19];	// lsu.scala:210:16
        ldq_17_bits_uop_pc_lob = _RANDOM[10'h12D][25:20];	// lsu.scala:210:16
        ldq_17_bits_uop_taken = _RANDOM[10'h12D][26];	// lsu.scala:210:16
        ldq_17_bits_uop_imm_packed = {_RANDOM[10'h12D][31:27], _RANDOM[10'h12E][14:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_csr_addr = _RANDOM[10'h12E][26:15];	// lsu.scala:210:16
        ldq_17_bits_uop_rob_idx = {_RANDOM[10'h12E][31:27], _RANDOM[10'h12F][1:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_ldq_idx = _RANDOM[10'h12F][6:2];	// lsu.scala:210:16
        ldq_17_bits_uop_stq_idx = _RANDOM[10'h12F][11:7];	// lsu.scala:210:16
        ldq_17_bits_uop_rxq_idx = _RANDOM[10'h12F][13:12];	// lsu.scala:210:16
        ldq_17_bits_uop_pdst = _RANDOM[10'h12F][20:14];	// lsu.scala:210:16
        ldq_17_bits_uop_prs1 = _RANDOM[10'h12F][27:21];	// lsu.scala:210:16
        ldq_17_bits_uop_prs2 = {_RANDOM[10'h12F][31:28], _RANDOM[10'h130][2:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_prs3 = _RANDOM[10'h130][9:3];	// lsu.scala:210:16
        ldq_17_bits_uop_ppred = _RANDOM[10'h130][14:10];	// lsu.scala:210:16
        ldq_17_bits_uop_prs1_busy = _RANDOM[10'h130][15];	// lsu.scala:210:16
        ldq_17_bits_uop_prs2_busy = _RANDOM[10'h130][16];	// lsu.scala:210:16
        ldq_17_bits_uop_prs3_busy = _RANDOM[10'h130][17];	// lsu.scala:210:16
        ldq_17_bits_uop_ppred_busy = _RANDOM[10'h130][18];	// lsu.scala:210:16
        ldq_17_bits_uop_stale_pdst = _RANDOM[10'h130][25:19];	// lsu.scala:210:16
        ldq_17_bits_uop_exception = _RANDOM[10'h130][26];	// lsu.scala:210:16
        ldq_17_bits_uop_exc_cause =
          {_RANDOM[10'h130][31:27], _RANDOM[10'h131], _RANDOM[10'h132][26:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_bypassable = _RANDOM[10'h132][27];	// lsu.scala:210:16
        ldq_17_bits_uop_mem_cmd = {_RANDOM[10'h132][31:28], _RANDOM[10'h133][0]};	// lsu.scala:210:16
        ldq_17_bits_uop_mem_size = _RANDOM[10'h133][2:1];	// lsu.scala:210:16
        ldq_17_bits_uop_mem_signed = _RANDOM[10'h133][3];	// lsu.scala:210:16
        ldq_17_bits_uop_is_fence = _RANDOM[10'h133][4];	// lsu.scala:210:16
        ldq_17_bits_uop_is_fencei = _RANDOM[10'h133][5];	// lsu.scala:210:16
        ldq_17_bits_uop_is_amo = _RANDOM[10'h133][6];	// lsu.scala:210:16
        ldq_17_bits_uop_uses_ldq = _RANDOM[10'h133][7];	// lsu.scala:210:16
        ldq_17_bits_uop_uses_stq = _RANDOM[10'h133][8];	// lsu.scala:210:16
        ldq_17_bits_uop_is_sys_pc2epc = _RANDOM[10'h133][9];	// lsu.scala:210:16
        ldq_17_bits_uop_is_unique = _RANDOM[10'h133][10];	// lsu.scala:210:16
        ldq_17_bits_uop_flush_on_commit = _RANDOM[10'h133][11];	// lsu.scala:210:16
        ldq_17_bits_uop_ldst_is_rs1 = _RANDOM[10'h133][12];	// lsu.scala:210:16
        ldq_17_bits_uop_ldst = _RANDOM[10'h133][18:13];	// lsu.scala:210:16
        ldq_17_bits_uop_lrs1 = _RANDOM[10'h133][24:19];	// lsu.scala:210:16
        ldq_17_bits_uop_lrs2 = _RANDOM[10'h133][30:25];	// lsu.scala:210:16
        ldq_17_bits_uop_lrs3 = {_RANDOM[10'h133][31], _RANDOM[10'h134][4:0]};	// lsu.scala:210:16
        ldq_17_bits_uop_ldst_val = _RANDOM[10'h134][5];	// lsu.scala:210:16
        ldq_17_bits_uop_dst_rtype = _RANDOM[10'h134][7:6];	// lsu.scala:210:16
        ldq_17_bits_uop_lrs1_rtype = _RANDOM[10'h134][9:8];	// lsu.scala:210:16
        ldq_17_bits_uop_lrs2_rtype = _RANDOM[10'h134][11:10];	// lsu.scala:210:16
        ldq_17_bits_uop_frs3_en = _RANDOM[10'h134][12];	// lsu.scala:210:16
        ldq_17_bits_uop_fp_val = _RANDOM[10'h134][13];	// lsu.scala:210:16
        ldq_17_bits_uop_fp_single = _RANDOM[10'h134][14];	// lsu.scala:210:16
        ldq_17_bits_uop_xcpt_pf_if = _RANDOM[10'h134][15];	// lsu.scala:210:16
        ldq_17_bits_uop_xcpt_ae_if = _RANDOM[10'h134][16];	// lsu.scala:210:16
        ldq_17_bits_uop_xcpt_ma_if = _RANDOM[10'h134][17];	// lsu.scala:210:16
        ldq_17_bits_uop_bp_debug_if = _RANDOM[10'h134][18];	// lsu.scala:210:16
        ldq_17_bits_uop_bp_xcpt_if = _RANDOM[10'h134][19];	// lsu.scala:210:16
        ldq_17_bits_uop_debug_fsrc = _RANDOM[10'h134][21:20];	// lsu.scala:210:16
        ldq_17_bits_uop_debug_tsrc = _RANDOM[10'h134][23:22];	// lsu.scala:210:16
        ldq_17_bits_addr_valid = _RANDOM[10'h134][24];	// lsu.scala:210:16
        ldq_17_bits_addr_bits =
          {_RANDOM[10'h134][31:25], _RANDOM[10'h135], _RANDOM[10'h136][0]};	// lsu.scala:210:16
        ldq_17_bits_addr_is_virtual = _RANDOM[10'h136][1];	// lsu.scala:210:16
        ldq_17_bits_addr_is_uncacheable = _RANDOM[10'h136][2];	// lsu.scala:210:16
        ldq_17_bits_executed = _RANDOM[10'h136][3];	// lsu.scala:210:16
        ldq_17_bits_succeeded = _RANDOM[10'h136][4];	// lsu.scala:210:16
        ldq_17_bits_order_fail = _RANDOM[10'h136][5];	// lsu.scala:210:16
        ldq_17_bits_observed = _RANDOM[10'h136][6];	// lsu.scala:210:16
        ldq_17_bits_st_dep_mask = _RANDOM[10'h136][30:7];	// lsu.scala:210:16
        ldq_17_bits_youngest_stq_idx = {_RANDOM[10'h136][31], _RANDOM[10'h137][3:0]};	// lsu.scala:210:16
        ldq_17_bits_forward_std_val = _RANDOM[10'h137][4];	// lsu.scala:210:16
        ldq_17_bits_forward_stq_idx = _RANDOM[10'h137][9:5];	// lsu.scala:210:16
        ldq_18_valid = _RANDOM[10'h139][10];	// lsu.scala:210:16
        ldq_18_bits_uop_uopc = _RANDOM[10'h139][17:11];	// lsu.scala:210:16
        ldq_18_bits_uop_inst = {_RANDOM[10'h139][31:18], _RANDOM[10'h13A][17:0]};	// lsu.scala:210:16
        ldq_18_bits_uop_debug_inst = {_RANDOM[10'h13A][31:18], _RANDOM[10'h13B][17:0]};	// lsu.scala:210:16
        ldq_18_bits_uop_is_rvc = _RANDOM[10'h13B][18];	// lsu.scala:210:16
        ldq_18_bits_uop_debug_pc = {_RANDOM[10'h13B][31:19], _RANDOM[10'h13C][26:0]};	// lsu.scala:210:16
        ldq_18_bits_uop_iq_type = _RANDOM[10'h13C][29:27];	// lsu.scala:210:16
        ldq_18_bits_uop_fu_code = {_RANDOM[10'h13C][31:30], _RANDOM[10'h13D][7:0]};	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_br_type = _RANDOM[10'h13D][11:8];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_op1_sel = _RANDOM[10'h13D][13:12];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_op2_sel = _RANDOM[10'h13D][16:14];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_imm_sel = _RANDOM[10'h13D][19:17];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_op_fcn = _RANDOM[10'h13D][23:20];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_fcn_dw = _RANDOM[10'h13D][24];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_csr_cmd = _RANDOM[10'h13D][27:25];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_is_load = _RANDOM[10'h13D][28];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_is_sta = _RANDOM[10'h13D][29];	// lsu.scala:210:16
        ldq_18_bits_uop_ctrl_is_std = _RANDOM[10'h13D][30];	// lsu.scala:210:16
        ldq_18_bits_uop_iw_state = {_RANDOM[10'h13D][31], _RANDOM[10'h13E][0]};	// lsu.scala:210:16
        ldq_18_bits_uop_iw_p1_poisoned = _RANDOM[10'h13E][1];	// lsu.scala:210:16
        ldq_18_bits_uop_iw_p2_poisoned = _RANDOM[10'h13E][2];	// lsu.scala:210:16
        ldq_18_bits_uop_is_br = _RANDOM[10'h13E][3];	// lsu.scala:210:16
        ldq_18_bits_uop_is_jalr = _RANDOM[10'h13E][4];	// lsu.scala:210:16
        ldq_18_bits_uop_is_jal = _RANDOM[10'h13E][5];	// lsu.scala:210:16
        ldq_18_bits_uop_is_sfb = _RANDOM[10'h13E][6];	// lsu.scala:210:16
        ldq_18_bits_uop_br_mask = _RANDOM[10'h13E][22:7];	// lsu.scala:210:16
        ldq_18_bits_uop_br_tag = _RANDOM[10'h13E][26:23];	// lsu.scala:210:16
        ldq_18_bits_uop_ftq_idx = _RANDOM[10'h13E][31:27];	// lsu.scala:210:16
        ldq_18_bits_uop_edge_inst = _RANDOM[10'h13F][0];	// lsu.scala:210:16
        ldq_18_bits_uop_pc_lob = _RANDOM[10'h13F][6:1];	// lsu.scala:210:16
        ldq_18_bits_uop_taken = _RANDOM[10'h13F][7];	// lsu.scala:210:16
        ldq_18_bits_uop_imm_packed = _RANDOM[10'h13F][27:8];	// lsu.scala:210:16
        ldq_18_bits_uop_csr_addr = {_RANDOM[10'h13F][31:28], _RANDOM[10'h140][7:0]};	// lsu.scala:210:16
        ldq_18_bits_uop_rob_idx = _RANDOM[10'h140][14:8];	// lsu.scala:210:16
        ldq_18_bits_uop_ldq_idx = _RANDOM[10'h140][19:15];	// lsu.scala:210:16
        ldq_18_bits_uop_stq_idx = _RANDOM[10'h140][24:20];	// lsu.scala:210:16
        ldq_18_bits_uop_rxq_idx = _RANDOM[10'h140][26:25];	// lsu.scala:210:16
        ldq_18_bits_uop_pdst = {_RANDOM[10'h140][31:27], _RANDOM[10'h141][1:0]};	// lsu.scala:210:16
        ldq_18_bits_uop_prs1 = _RANDOM[10'h141][8:2];	// lsu.scala:210:16
        ldq_18_bits_uop_prs2 = _RANDOM[10'h141][15:9];	// lsu.scala:210:16
        ldq_18_bits_uop_prs3 = _RANDOM[10'h141][22:16];	// lsu.scala:210:16
        ldq_18_bits_uop_ppred = _RANDOM[10'h141][27:23];	// lsu.scala:210:16
        ldq_18_bits_uop_prs1_busy = _RANDOM[10'h141][28];	// lsu.scala:210:16
        ldq_18_bits_uop_prs2_busy = _RANDOM[10'h141][29];	// lsu.scala:210:16
        ldq_18_bits_uop_prs3_busy = _RANDOM[10'h141][30];	// lsu.scala:210:16
        ldq_18_bits_uop_ppred_busy = _RANDOM[10'h141][31];	// lsu.scala:210:16
        ldq_18_bits_uop_stale_pdst = _RANDOM[10'h142][6:0];	// lsu.scala:210:16
        ldq_18_bits_uop_exception = _RANDOM[10'h142][7];	// lsu.scala:210:16
        ldq_18_bits_uop_exc_cause =
          {_RANDOM[10'h142][31:8], _RANDOM[10'h143], _RANDOM[10'h144][7:0]};	// lsu.scala:210:16
        ldq_18_bits_uop_bypassable = _RANDOM[10'h144][8];	// lsu.scala:210:16
        ldq_18_bits_uop_mem_cmd = _RANDOM[10'h144][13:9];	// lsu.scala:210:16
        ldq_18_bits_uop_mem_size = _RANDOM[10'h144][15:14];	// lsu.scala:210:16
        ldq_18_bits_uop_mem_signed = _RANDOM[10'h144][16];	// lsu.scala:210:16
        ldq_18_bits_uop_is_fence = _RANDOM[10'h144][17];	// lsu.scala:210:16
        ldq_18_bits_uop_is_fencei = _RANDOM[10'h144][18];	// lsu.scala:210:16
        ldq_18_bits_uop_is_amo = _RANDOM[10'h144][19];	// lsu.scala:210:16
        ldq_18_bits_uop_uses_ldq = _RANDOM[10'h144][20];	// lsu.scala:210:16
        ldq_18_bits_uop_uses_stq = _RANDOM[10'h144][21];	// lsu.scala:210:16
        ldq_18_bits_uop_is_sys_pc2epc = _RANDOM[10'h144][22];	// lsu.scala:210:16
        ldq_18_bits_uop_is_unique = _RANDOM[10'h144][23];	// lsu.scala:210:16
        ldq_18_bits_uop_flush_on_commit = _RANDOM[10'h144][24];	// lsu.scala:210:16
        ldq_18_bits_uop_ldst_is_rs1 = _RANDOM[10'h144][25];	// lsu.scala:210:16
        ldq_18_bits_uop_ldst = _RANDOM[10'h144][31:26];	// lsu.scala:210:16
        ldq_18_bits_uop_lrs1 = _RANDOM[10'h145][5:0];	// lsu.scala:210:16
        ldq_18_bits_uop_lrs2 = _RANDOM[10'h145][11:6];	// lsu.scala:210:16
        ldq_18_bits_uop_lrs3 = _RANDOM[10'h145][17:12];	// lsu.scala:210:16
        ldq_18_bits_uop_ldst_val = _RANDOM[10'h145][18];	// lsu.scala:210:16
        ldq_18_bits_uop_dst_rtype = _RANDOM[10'h145][20:19];	// lsu.scala:210:16
        ldq_18_bits_uop_lrs1_rtype = _RANDOM[10'h145][22:21];	// lsu.scala:210:16
        ldq_18_bits_uop_lrs2_rtype = _RANDOM[10'h145][24:23];	// lsu.scala:210:16
        ldq_18_bits_uop_frs3_en = _RANDOM[10'h145][25];	// lsu.scala:210:16
        ldq_18_bits_uop_fp_val = _RANDOM[10'h145][26];	// lsu.scala:210:16
        ldq_18_bits_uop_fp_single = _RANDOM[10'h145][27];	// lsu.scala:210:16
        ldq_18_bits_uop_xcpt_pf_if = _RANDOM[10'h145][28];	// lsu.scala:210:16
        ldq_18_bits_uop_xcpt_ae_if = _RANDOM[10'h145][29];	// lsu.scala:210:16
        ldq_18_bits_uop_xcpt_ma_if = _RANDOM[10'h145][30];	// lsu.scala:210:16
        ldq_18_bits_uop_bp_debug_if = _RANDOM[10'h145][31];	// lsu.scala:210:16
        ldq_18_bits_uop_bp_xcpt_if = _RANDOM[10'h146][0];	// lsu.scala:210:16
        ldq_18_bits_uop_debug_fsrc = _RANDOM[10'h146][2:1];	// lsu.scala:210:16
        ldq_18_bits_uop_debug_tsrc = _RANDOM[10'h146][4:3];	// lsu.scala:210:16
        ldq_18_bits_addr_valid = _RANDOM[10'h146][5];	// lsu.scala:210:16
        ldq_18_bits_addr_bits = {_RANDOM[10'h146][31:6], _RANDOM[10'h147][13:0]};	// lsu.scala:210:16
        ldq_18_bits_addr_is_virtual = _RANDOM[10'h147][14];	// lsu.scala:210:16
        ldq_18_bits_addr_is_uncacheable = _RANDOM[10'h147][15];	// lsu.scala:210:16
        ldq_18_bits_executed = _RANDOM[10'h147][16];	// lsu.scala:210:16
        ldq_18_bits_succeeded = _RANDOM[10'h147][17];	// lsu.scala:210:16
        ldq_18_bits_order_fail = _RANDOM[10'h147][18];	// lsu.scala:210:16
        ldq_18_bits_observed = _RANDOM[10'h147][19];	// lsu.scala:210:16
        ldq_18_bits_st_dep_mask = {_RANDOM[10'h147][31:20], _RANDOM[10'h148][11:0]};	// lsu.scala:210:16
        ldq_18_bits_youngest_stq_idx = _RANDOM[10'h148][16:12];	// lsu.scala:210:16
        ldq_18_bits_forward_std_val = _RANDOM[10'h148][17];	// lsu.scala:210:16
        ldq_18_bits_forward_stq_idx = _RANDOM[10'h148][22:18];	// lsu.scala:210:16
        ldq_19_valid = _RANDOM[10'h14A][23];	// lsu.scala:210:16
        ldq_19_bits_uop_uopc = _RANDOM[10'h14A][30:24];	// lsu.scala:210:16
        ldq_19_bits_uop_inst = {_RANDOM[10'h14A][31], _RANDOM[10'h14B][30:0]};	// lsu.scala:210:16
        ldq_19_bits_uop_debug_inst = {_RANDOM[10'h14B][31], _RANDOM[10'h14C][30:0]};	// lsu.scala:210:16
        ldq_19_bits_uop_is_rvc = _RANDOM[10'h14C][31];	// lsu.scala:210:16
        ldq_19_bits_uop_debug_pc = {_RANDOM[10'h14D], _RANDOM[10'h14E][7:0]};	// lsu.scala:210:16
        ldq_19_bits_uop_iq_type = _RANDOM[10'h14E][10:8];	// lsu.scala:210:16
        ldq_19_bits_uop_fu_code = _RANDOM[10'h14E][20:11];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_br_type = _RANDOM[10'h14E][24:21];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_op1_sel = _RANDOM[10'h14E][26:25];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_op2_sel = _RANDOM[10'h14E][29:27];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_imm_sel = {_RANDOM[10'h14E][31:30], _RANDOM[10'h14F][0]};	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_op_fcn = _RANDOM[10'h14F][4:1];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_fcn_dw = _RANDOM[10'h14F][5];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_csr_cmd = _RANDOM[10'h14F][8:6];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_is_load = _RANDOM[10'h14F][9];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_is_sta = _RANDOM[10'h14F][10];	// lsu.scala:210:16
        ldq_19_bits_uop_ctrl_is_std = _RANDOM[10'h14F][11];	// lsu.scala:210:16
        ldq_19_bits_uop_iw_state = _RANDOM[10'h14F][13:12];	// lsu.scala:210:16
        ldq_19_bits_uop_iw_p1_poisoned = _RANDOM[10'h14F][14];	// lsu.scala:210:16
        ldq_19_bits_uop_iw_p2_poisoned = _RANDOM[10'h14F][15];	// lsu.scala:210:16
        ldq_19_bits_uop_is_br = _RANDOM[10'h14F][16];	// lsu.scala:210:16
        ldq_19_bits_uop_is_jalr = _RANDOM[10'h14F][17];	// lsu.scala:210:16
        ldq_19_bits_uop_is_jal = _RANDOM[10'h14F][18];	// lsu.scala:210:16
        ldq_19_bits_uop_is_sfb = _RANDOM[10'h14F][19];	// lsu.scala:210:16
        ldq_19_bits_uop_br_mask = {_RANDOM[10'h14F][31:20], _RANDOM[10'h150][3:0]};	// lsu.scala:210:16
        ldq_19_bits_uop_br_tag = _RANDOM[10'h150][7:4];	// lsu.scala:210:16
        ldq_19_bits_uop_ftq_idx = _RANDOM[10'h150][12:8];	// lsu.scala:210:16
        ldq_19_bits_uop_edge_inst = _RANDOM[10'h150][13];	// lsu.scala:210:16
        ldq_19_bits_uop_pc_lob = _RANDOM[10'h150][19:14];	// lsu.scala:210:16
        ldq_19_bits_uop_taken = _RANDOM[10'h150][20];	// lsu.scala:210:16
        ldq_19_bits_uop_imm_packed = {_RANDOM[10'h150][31:21], _RANDOM[10'h151][8:0]};	// lsu.scala:210:16
        ldq_19_bits_uop_csr_addr = _RANDOM[10'h151][20:9];	// lsu.scala:210:16
        ldq_19_bits_uop_rob_idx = _RANDOM[10'h151][27:21];	// lsu.scala:210:16
        ldq_19_bits_uop_ldq_idx = {_RANDOM[10'h151][31:28], _RANDOM[10'h152][0]};	// lsu.scala:210:16
        ldq_19_bits_uop_stq_idx = _RANDOM[10'h152][5:1];	// lsu.scala:210:16
        ldq_19_bits_uop_rxq_idx = _RANDOM[10'h152][7:6];	// lsu.scala:210:16
        ldq_19_bits_uop_pdst = _RANDOM[10'h152][14:8];	// lsu.scala:210:16
        ldq_19_bits_uop_prs1 = _RANDOM[10'h152][21:15];	// lsu.scala:210:16
        ldq_19_bits_uop_prs2 = _RANDOM[10'h152][28:22];	// lsu.scala:210:16
        ldq_19_bits_uop_prs3 = {_RANDOM[10'h152][31:29], _RANDOM[10'h153][3:0]};	// lsu.scala:210:16
        ldq_19_bits_uop_ppred = _RANDOM[10'h153][8:4];	// lsu.scala:210:16
        ldq_19_bits_uop_prs1_busy = _RANDOM[10'h153][9];	// lsu.scala:210:16
        ldq_19_bits_uop_prs2_busy = _RANDOM[10'h153][10];	// lsu.scala:210:16
        ldq_19_bits_uop_prs3_busy = _RANDOM[10'h153][11];	// lsu.scala:210:16
        ldq_19_bits_uop_ppred_busy = _RANDOM[10'h153][12];	// lsu.scala:210:16
        ldq_19_bits_uop_stale_pdst = _RANDOM[10'h153][19:13];	// lsu.scala:210:16
        ldq_19_bits_uop_exception = _RANDOM[10'h153][20];	// lsu.scala:210:16
        ldq_19_bits_uop_exc_cause =
          {_RANDOM[10'h153][31:21], _RANDOM[10'h154], _RANDOM[10'h155][20:0]};	// lsu.scala:210:16
        ldq_19_bits_uop_bypassable = _RANDOM[10'h155][21];	// lsu.scala:210:16
        ldq_19_bits_uop_mem_cmd = _RANDOM[10'h155][26:22];	// lsu.scala:210:16
        ldq_19_bits_uop_mem_size = _RANDOM[10'h155][28:27];	// lsu.scala:210:16
        ldq_19_bits_uop_mem_signed = _RANDOM[10'h155][29];	// lsu.scala:210:16
        ldq_19_bits_uop_is_fence = _RANDOM[10'h155][30];	// lsu.scala:210:16
        ldq_19_bits_uop_is_fencei = _RANDOM[10'h155][31];	// lsu.scala:210:16
        ldq_19_bits_uop_is_amo = _RANDOM[10'h156][0];	// lsu.scala:210:16
        ldq_19_bits_uop_uses_ldq = _RANDOM[10'h156][1];	// lsu.scala:210:16
        ldq_19_bits_uop_uses_stq = _RANDOM[10'h156][2];	// lsu.scala:210:16
        ldq_19_bits_uop_is_sys_pc2epc = _RANDOM[10'h156][3];	// lsu.scala:210:16
        ldq_19_bits_uop_is_unique = _RANDOM[10'h156][4];	// lsu.scala:210:16
        ldq_19_bits_uop_flush_on_commit = _RANDOM[10'h156][5];	// lsu.scala:210:16
        ldq_19_bits_uop_ldst_is_rs1 = _RANDOM[10'h156][6];	// lsu.scala:210:16
        ldq_19_bits_uop_ldst = _RANDOM[10'h156][12:7];	// lsu.scala:210:16
        ldq_19_bits_uop_lrs1 = _RANDOM[10'h156][18:13];	// lsu.scala:210:16
        ldq_19_bits_uop_lrs2 = _RANDOM[10'h156][24:19];	// lsu.scala:210:16
        ldq_19_bits_uop_lrs3 = _RANDOM[10'h156][30:25];	// lsu.scala:210:16
        ldq_19_bits_uop_ldst_val = _RANDOM[10'h156][31];	// lsu.scala:210:16
        ldq_19_bits_uop_dst_rtype = _RANDOM[10'h157][1:0];	// lsu.scala:210:16
        ldq_19_bits_uop_lrs1_rtype = _RANDOM[10'h157][3:2];	// lsu.scala:210:16
        ldq_19_bits_uop_lrs2_rtype = _RANDOM[10'h157][5:4];	// lsu.scala:210:16
        ldq_19_bits_uop_frs3_en = _RANDOM[10'h157][6];	// lsu.scala:210:16
        ldq_19_bits_uop_fp_val = _RANDOM[10'h157][7];	// lsu.scala:210:16
        ldq_19_bits_uop_fp_single = _RANDOM[10'h157][8];	// lsu.scala:210:16
        ldq_19_bits_uop_xcpt_pf_if = _RANDOM[10'h157][9];	// lsu.scala:210:16
        ldq_19_bits_uop_xcpt_ae_if = _RANDOM[10'h157][10];	// lsu.scala:210:16
        ldq_19_bits_uop_xcpt_ma_if = _RANDOM[10'h157][11];	// lsu.scala:210:16
        ldq_19_bits_uop_bp_debug_if = _RANDOM[10'h157][12];	// lsu.scala:210:16
        ldq_19_bits_uop_bp_xcpt_if = _RANDOM[10'h157][13];	// lsu.scala:210:16
        ldq_19_bits_uop_debug_fsrc = _RANDOM[10'h157][15:14];	// lsu.scala:210:16
        ldq_19_bits_uop_debug_tsrc = _RANDOM[10'h157][17:16];	// lsu.scala:210:16
        ldq_19_bits_addr_valid = _RANDOM[10'h157][18];	// lsu.scala:210:16
        ldq_19_bits_addr_bits = {_RANDOM[10'h157][31:19], _RANDOM[10'h158][26:0]};	// lsu.scala:210:16
        ldq_19_bits_addr_is_virtual = _RANDOM[10'h158][27];	// lsu.scala:210:16
        ldq_19_bits_addr_is_uncacheable = _RANDOM[10'h158][28];	// lsu.scala:210:16
        ldq_19_bits_executed = _RANDOM[10'h158][29];	// lsu.scala:210:16
        ldq_19_bits_succeeded = _RANDOM[10'h158][30];	// lsu.scala:210:16
        ldq_19_bits_order_fail = _RANDOM[10'h158][31];	// lsu.scala:210:16
        ldq_19_bits_observed = _RANDOM[10'h159][0];	// lsu.scala:210:16
        ldq_19_bits_st_dep_mask = _RANDOM[10'h159][24:1];	// lsu.scala:210:16
        ldq_19_bits_youngest_stq_idx = _RANDOM[10'h159][29:25];	// lsu.scala:210:16
        ldq_19_bits_forward_std_val = _RANDOM[10'h159][30];	// lsu.scala:210:16
        ldq_19_bits_forward_stq_idx = {_RANDOM[10'h159][31], _RANDOM[10'h15A][3:0]};	// lsu.scala:210:16
        ldq_20_valid = _RANDOM[10'h15C][4];	// lsu.scala:210:16
        ldq_20_bits_uop_uopc = _RANDOM[10'h15C][11:5];	// lsu.scala:210:16
        ldq_20_bits_uop_inst = {_RANDOM[10'h15C][31:12], _RANDOM[10'h15D][11:0]};	// lsu.scala:210:16
        ldq_20_bits_uop_debug_inst = {_RANDOM[10'h15D][31:12], _RANDOM[10'h15E][11:0]};	// lsu.scala:210:16
        ldq_20_bits_uop_is_rvc = _RANDOM[10'h15E][12];	// lsu.scala:210:16
        ldq_20_bits_uop_debug_pc = {_RANDOM[10'h15E][31:13], _RANDOM[10'h15F][20:0]};	// lsu.scala:210:16
        ldq_20_bits_uop_iq_type = _RANDOM[10'h15F][23:21];	// lsu.scala:210:16
        ldq_20_bits_uop_fu_code = {_RANDOM[10'h15F][31:24], _RANDOM[10'h160][1:0]};	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_br_type = _RANDOM[10'h160][5:2];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_op1_sel = _RANDOM[10'h160][7:6];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_op2_sel = _RANDOM[10'h160][10:8];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_imm_sel = _RANDOM[10'h160][13:11];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_op_fcn = _RANDOM[10'h160][17:14];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_fcn_dw = _RANDOM[10'h160][18];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_csr_cmd = _RANDOM[10'h160][21:19];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_is_load = _RANDOM[10'h160][22];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_is_sta = _RANDOM[10'h160][23];	// lsu.scala:210:16
        ldq_20_bits_uop_ctrl_is_std = _RANDOM[10'h160][24];	// lsu.scala:210:16
        ldq_20_bits_uop_iw_state = _RANDOM[10'h160][26:25];	// lsu.scala:210:16
        ldq_20_bits_uop_iw_p1_poisoned = _RANDOM[10'h160][27];	// lsu.scala:210:16
        ldq_20_bits_uop_iw_p2_poisoned = _RANDOM[10'h160][28];	// lsu.scala:210:16
        ldq_20_bits_uop_is_br = _RANDOM[10'h160][29];	// lsu.scala:210:16
        ldq_20_bits_uop_is_jalr = _RANDOM[10'h160][30];	// lsu.scala:210:16
        ldq_20_bits_uop_is_jal = _RANDOM[10'h160][31];	// lsu.scala:210:16
        ldq_20_bits_uop_is_sfb = _RANDOM[10'h161][0];	// lsu.scala:210:16
        ldq_20_bits_uop_br_mask = _RANDOM[10'h161][16:1];	// lsu.scala:210:16
        ldq_20_bits_uop_br_tag = _RANDOM[10'h161][20:17];	// lsu.scala:210:16
        ldq_20_bits_uop_ftq_idx = _RANDOM[10'h161][25:21];	// lsu.scala:210:16
        ldq_20_bits_uop_edge_inst = _RANDOM[10'h161][26];	// lsu.scala:210:16
        ldq_20_bits_uop_pc_lob = {_RANDOM[10'h161][31:27], _RANDOM[10'h162][0]};	// lsu.scala:210:16
        ldq_20_bits_uop_taken = _RANDOM[10'h162][1];	// lsu.scala:210:16
        ldq_20_bits_uop_imm_packed = _RANDOM[10'h162][21:2];	// lsu.scala:210:16
        ldq_20_bits_uop_csr_addr = {_RANDOM[10'h162][31:22], _RANDOM[10'h163][1:0]};	// lsu.scala:210:16
        ldq_20_bits_uop_rob_idx = _RANDOM[10'h163][8:2];	// lsu.scala:210:16
        ldq_20_bits_uop_ldq_idx = _RANDOM[10'h163][13:9];	// lsu.scala:210:16
        ldq_20_bits_uop_stq_idx = _RANDOM[10'h163][18:14];	// lsu.scala:210:16
        ldq_20_bits_uop_rxq_idx = _RANDOM[10'h163][20:19];	// lsu.scala:210:16
        ldq_20_bits_uop_pdst = _RANDOM[10'h163][27:21];	// lsu.scala:210:16
        ldq_20_bits_uop_prs1 = {_RANDOM[10'h163][31:28], _RANDOM[10'h164][2:0]};	// lsu.scala:210:16
        ldq_20_bits_uop_prs2 = _RANDOM[10'h164][9:3];	// lsu.scala:210:16
        ldq_20_bits_uop_prs3 = _RANDOM[10'h164][16:10];	// lsu.scala:210:16
        ldq_20_bits_uop_ppred = _RANDOM[10'h164][21:17];	// lsu.scala:210:16
        ldq_20_bits_uop_prs1_busy = _RANDOM[10'h164][22];	// lsu.scala:210:16
        ldq_20_bits_uop_prs2_busy = _RANDOM[10'h164][23];	// lsu.scala:210:16
        ldq_20_bits_uop_prs3_busy = _RANDOM[10'h164][24];	// lsu.scala:210:16
        ldq_20_bits_uop_ppred_busy = _RANDOM[10'h164][25];	// lsu.scala:210:16
        ldq_20_bits_uop_stale_pdst = {_RANDOM[10'h164][31:26], _RANDOM[10'h165][0]};	// lsu.scala:210:16
        ldq_20_bits_uop_exception = _RANDOM[10'h165][1];	// lsu.scala:210:16
        ldq_20_bits_uop_exc_cause =
          {_RANDOM[10'h165][31:2], _RANDOM[10'h166], _RANDOM[10'h167][1:0]};	// lsu.scala:210:16
        ldq_20_bits_uop_bypassable = _RANDOM[10'h167][2];	// lsu.scala:210:16
        ldq_20_bits_uop_mem_cmd = _RANDOM[10'h167][7:3];	// lsu.scala:210:16
        ldq_20_bits_uop_mem_size = _RANDOM[10'h167][9:8];	// lsu.scala:210:16
        ldq_20_bits_uop_mem_signed = _RANDOM[10'h167][10];	// lsu.scala:210:16
        ldq_20_bits_uop_is_fence = _RANDOM[10'h167][11];	// lsu.scala:210:16
        ldq_20_bits_uop_is_fencei = _RANDOM[10'h167][12];	// lsu.scala:210:16
        ldq_20_bits_uop_is_amo = _RANDOM[10'h167][13];	// lsu.scala:210:16
        ldq_20_bits_uop_uses_ldq = _RANDOM[10'h167][14];	// lsu.scala:210:16
        ldq_20_bits_uop_uses_stq = _RANDOM[10'h167][15];	// lsu.scala:210:16
        ldq_20_bits_uop_is_sys_pc2epc = _RANDOM[10'h167][16];	// lsu.scala:210:16
        ldq_20_bits_uop_is_unique = _RANDOM[10'h167][17];	// lsu.scala:210:16
        ldq_20_bits_uop_flush_on_commit = _RANDOM[10'h167][18];	// lsu.scala:210:16
        ldq_20_bits_uop_ldst_is_rs1 = _RANDOM[10'h167][19];	// lsu.scala:210:16
        ldq_20_bits_uop_ldst = _RANDOM[10'h167][25:20];	// lsu.scala:210:16
        ldq_20_bits_uop_lrs1 = _RANDOM[10'h167][31:26];	// lsu.scala:210:16
        ldq_20_bits_uop_lrs2 = _RANDOM[10'h168][5:0];	// lsu.scala:210:16
        ldq_20_bits_uop_lrs3 = _RANDOM[10'h168][11:6];	// lsu.scala:210:16
        ldq_20_bits_uop_ldst_val = _RANDOM[10'h168][12];	// lsu.scala:210:16
        ldq_20_bits_uop_dst_rtype = _RANDOM[10'h168][14:13];	// lsu.scala:210:16
        ldq_20_bits_uop_lrs1_rtype = _RANDOM[10'h168][16:15];	// lsu.scala:210:16
        ldq_20_bits_uop_lrs2_rtype = _RANDOM[10'h168][18:17];	// lsu.scala:210:16
        ldq_20_bits_uop_frs3_en = _RANDOM[10'h168][19];	// lsu.scala:210:16
        ldq_20_bits_uop_fp_val = _RANDOM[10'h168][20];	// lsu.scala:210:16
        ldq_20_bits_uop_fp_single = _RANDOM[10'h168][21];	// lsu.scala:210:16
        ldq_20_bits_uop_xcpt_pf_if = _RANDOM[10'h168][22];	// lsu.scala:210:16
        ldq_20_bits_uop_xcpt_ae_if = _RANDOM[10'h168][23];	// lsu.scala:210:16
        ldq_20_bits_uop_xcpt_ma_if = _RANDOM[10'h168][24];	// lsu.scala:210:16
        ldq_20_bits_uop_bp_debug_if = _RANDOM[10'h168][25];	// lsu.scala:210:16
        ldq_20_bits_uop_bp_xcpt_if = _RANDOM[10'h168][26];	// lsu.scala:210:16
        ldq_20_bits_uop_debug_fsrc = _RANDOM[10'h168][28:27];	// lsu.scala:210:16
        ldq_20_bits_uop_debug_tsrc = _RANDOM[10'h168][30:29];	// lsu.scala:210:16
        ldq_20_bits_addr_valid = _RANDOM[10'h168][31];	// lsu.scala:210:16
        ldq_20_bits_addr_bits = {_RANDOM[10'h169], _RANDOM[10'h16A][7:0]};	// lsu.scala:210:16
        ldq_20_bits_addr_is_virtual = _RANDOM[10'h16A][8];	// lsu.scala:210:16
        ldq_20_bits_addr_is_uncacheable = _RANDOM[10'h16A][9];	// lsu.scala:210:16
        ldq_20_bits_executed = _RANDOM[10'h16A][10];	// lsu.scala:210:16
        ldq_20_bits_succeeded = _RANDOM[10'h16A][11];	// lsu.scala:210:16
        ldq_20_bits_order_fail = _RANDOM[10'h16A][12];	// lsu.scala:210:16
        ldq_20_bits_observed = _RANDOM[10'h16A][13];	// lsu.scala:210:16
        ldq_20_bits_st_dep_mask = {_RANDOM[10'h16A][31:14], _RANDOM[10'h16B][5:0]};	// lsu.scala:210:16
        ldq_20_bits_youngest_stq_idx = _RANDOM[10'h16B][10:6];	// lsu.scala:210:16
        ldq_20_bits_forward_std_val = _RANDOM[10'h16B][11];	// lsu.scala:210:16
        ldq_20_bits_forward_stq_idx = _RANDOM[10'h16B][16:12];	// lsu.scala:210:16
        ldq_21_valid = _RANDOM[10'h16D][17];	// lsu.scala:210:16
        ldq_21_bits_uop_uopc = _RANDOM[10'h16D][24:18];	// lsu.scala:210:16
        ldq_21_bits_uop_inst = {_RANDOM[10'h16D][31:25], _RANDOM[10'h16E][24:0]};	// lsu.scala:210:16
        ldq_21_bits_uop_debug_inst = {_RANDOM[10'h16E][31:25], _RANDOM[10'h16F][24:0]};	// lsu.scala:210:16
        ldq_21_bits_uop_is_rvc = _RANDOM[10'h16F][25];	// lsu.scala:210:16
        ldq_21_bits_uop_debug_pc =
          {_RANDOM[10'h16F][31:26], _RANDOM[10'h170], _RANDOM[10'h171][1:0]};	// lsu.scala:210:16
        ldq_21_bits_uop_iq_type = _RANDOM[10'h171][4:2];	// lsu.scala:210:16
        ldq_21_bits_uop_fu_code = _RANDOM[10'h171][14:5];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_br_type = _RANDOM[10'h171][18:15];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_op1_sel = _RANDOM[10'h171][20:19];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_op2_sel = _RANDOM[10'h171][23:21];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_imm_sel = _RANDOM[10'h171][26:24];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_op_fcn = _RANDOM[10'h171][30:27];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_fcn_dw = _RANDOM[10'h171][31];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_csr_cmd = _RANDOM[10'h172][2:0];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_is_load = _RANDOM[10'h172][3];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_is_sta = _RANDOM[10'h172][4];	// lsu.scala:210:16
        ldq_21_bits_uop_ctrl_is_std = _RANDOM[10'h172][5];	// lsu.scala:210:16
        ldq_21_bits_uop_iw_state = _RANDOM[10'h172][7:6];	// lsu.scala:210:16
        ldq_21_bits_uop_iw_p1_poisoned = _RANDOM[10'h172][8];	// lsu.scala:210:16
        ldq_21_bits_uop_iw_p2_poisoned = _RANDOM[10'h172][9];	// lsu.scala:210:16
        ldq_21_bits_uop_is_br = _RANDOM[10'h172][10];	// lsu.scala:210:16
        ldq_21_bits_uop_is_jalr = _RANDOM[10'h172][11];	// lsu.scala:210:16
        ldq_21_bits_uop_is_jal = _RANDOM[10'h172][12];	// lsu.scala:210:16
        ldq_21_bits_uop_is_sfb = _RANDOM[10'h172][13];	// lsu.scala:210:16
        ldq_21_bits_uop_br_mask = _RANDOM[10'h172][29:14];	// lsu.scala:210:16
        ldq_21_bits_uop_br_tag = {_RANDOM[10'h172][31:30], _RANDOM[10'h173][1:0]};	// lsu.scala:210:16
        ldq_21_bits_uop_ftq_idx = _RANDOM[10'h173][6:2];	// lsu.scala:210:16
        ldq_21_bits_uop_edge_inst = _RANDOM[10'h173][7];	// lsu.scala:210:16
        ldq_21_bits_uop_pc_lob = _RANDOM[10'h173][13:8];	// lsu.scala:210:16
        ldq_21_bits_uop_taken = _RANDOM[10'h173][14];	// lsu.scala:210:16
        ldq_21_bits_uop_imm_packed = {_RANDOM[10'h173][31:15], _RANDOM[10'h174][2:0]};	// lsu.scala:210:16
        ldq_21_bits_uop_csr_addr = _RANDOM[10'h174][14:3];	// lsu.scala:210:16
        ldq_21_bits_uop_rob_idx = _RANDOM[10'h174][21:15];	// lsu.scala:210:16
        ldq_21_bits_uop_ldq_idx = _RANDOM[10'h174][26:22];	// lsu.scala:210:16
        ldq_21_bits_uop_stq_idx = _RANDOM[10'h174][31:27];	// lsu.scala:210:16
        ldq_21_bits_uop_rxq_idx = _RANDOM[10'h175][1:0];	// lsu.scala:210:16
        ldq_21_bits_uop_pdst = _RANDOM[10'h175][8:2];	// lsu.scala:210:16
        ldq_21_bits_uop_prs1 = _RANDOM[10'h175][15:9];	// lsu.scala:210:16
        ldq_21_bits_uop_prs2 = _RANDOM[10'h175][22:16];	// lsu.scala:210:16
        ldq_21_bits_uop_prs3 = _RANDOM[10'h175][29:23];	// lsu.scala:210:16
        ldq_21_bits_uop_ppred = {_RANDOM[10'h175][31:30], _RANDOM[10'h176][2:0]};	// lsu.scala:210:16
        ldq_21_bits_uop_prs1_busy = _RANDOM[10'h176][3];	// lsu.scala:210:16
        ldq_21_bits_uop_prs2_busy = _RANDOM[10'h176][4];	// lsu.scala:210:16
        ldq_21_bits_uop_prs3_busy = _RANDOM[10'h176][5];	// lsu.scala:210:16
        ldq_21_bits_uop_ppred_busy = _RANDOM[10'h176][6];	// lsu.scala:210:16
        ldq_21_bits_uop_stale_pdst = _RANDOM[10'h176][13:7];	// lsu.scala:210:16
        ldq_21_bits_uop_exception = _RANDOM[10'h176][14];	// lsu.scala:210:16
        ldq_21_bits_uop_exc_cause =
          {_RANDOM[10'h176][31:15], _RANDOM[10'h177], _RANDOM[10'h178][14:0]};	// lsu.scala:210:16
        ldq_21_bits_uop_bypassable = _RANDOM[10'h178][15];	// lsu.scala:210:16
        ldq_21_bits_uop_mem_cmd = _RANDOM[10'h178][20:16];	// lsu.scala:210:16
        ldq_21_bits_uop_mem_size = _RANDOM[10'h178][22:21];	// lsu.scala:210:16
        ldq_21_bits_uop_mem_signed = _RANDOM[10'h178][23];	// lsu.scala:210:16
        ldq_21_bits_uop_is_fence = _RANDOM[10'h178][24];	// lsu.scala:210:16
        ldq_21_bits_uop_is_fencei = _RANDOM[10'h178][25];	// lsu.scala:210:16
        ldq_21_bits_uop_is_amo = _RANDOM[10'h178][26];	// lsu.scala:210:16
        ldq_21_bits_uop_uses_ldq = _RANDOM[10'h178][27];	// lsu.scala:210:16
        ldq_21_bits_uop_uses_stq = _RANDOM[10'h178][28];	// lsu.scala:210:16
        ldq_21_bits_uop_is_sys_pc2epc = _RANDOM[10'h178][29];	// lsu.scala:210:16
        ldq_21_bits_uop_is_unique = _RANDOM[10'h178][30];	// lsu.scala:210:16
        ldq_21_bits_uop_flush_on_commit = _RANDOM[10'h178][31];	// lsu.scala:210:16
        ldq_21_bits_uop_ldst_is_rs1 = _RANDOM[10'h179][0];	// lsu.scala:210:16
        ldq_21_bits_uop_ldst = _RANDOM[10'h179][6:1];	// lsu.scala:210:16
        ldq_21_bits_uop_lrs1 = _RANDOM[10'h179][12:7];	// lsu.scala:210:16
        ldq_21_bits_uop_lrs2 = _RANDOM[10'h179][18:13];	// lsu.scala:210:16
        ldq_21_bits_uop_lrs3 = _RANDOM[10'h179][24:19];	// lsu.scala:210:16
        ldq_21_bits_uop_ldst_val = _RANDOM[10'h179][25];	// lsu.scala:210:16
        ldq_21_bits_uop_dst_rtype = _RANDOM[10'h179][27:26];	// lsu.scala:210:16
        ldq_21_bits_uop_lrs1_rtype = _RANDOM[10'h179][29:28];	// lsu.scala:210:16
        ldq_21_bits_uop_lrs2_rtype = _RANDOM[10'h179][31:30];	// lsu.scala:210:16
        ldq_21_bits_uop_frs3_en = _RANDOM[10'h17A][0];	// lsu.scala:210:16
        ldq_21_bits_uop_fp_val = _RANDOM[10'h17A][1];	// lsu.scala:210:16
        ldq_21_bits_uop_fp_single = _RANDOM[10'h17A][2];	// lsu.scala:210:16
        ldq_21_bits_uop_xcpt_pf_if = _RANDOM[10'h17A][3];	// lsu.scala:210:16
        ldq_21_bits_uop_xcpt_ae_if = _RANDOM[10'h17A][4];	// lsu.scala:210:16
        ldq_21_bits_uop_xcpt_ma_if = _RANDOM[10'h17A][5];	// lsu.scala:210:16
        ldq_21_bits_uop_bp_debug_if = _RANDOM[10'h17A][6];	// lsu.scala:210:16
        ldq_21_bits_uop_bp_xcpt_if = _RANDOM[10'h17A][7];	// lsu.scala:210:16
        ldq_21_bits_uop_debug_fsrc = _RANDOM[10'h17A][9:8];	// lsu.scala:210:16
        ldq_21_bits_uop_debug_tsrc = _RANDOM[10'h17A][11:10];	// lsu.scala:210:16
        ldq_21_bits_addr_valid = _RANDOM[10'h17A][12];	// lsu.scala:210:16
        ldq_21_bits_addr_bits = {_RANDOM[10'h17A][31:13], _RANDOM[10'h17B][20:0]};	// lsu.scala:210:16
        ldq_21_bits_addr_is_virtual = _RANDOM[10'h17B][21];	// lsu.scala:210:16
        ldq_21_bits_addr_is_uncacheable = _RANDOM[10'h17B][22];	// lsu.scala:210:16
        ldq_21_bits_executed = _RANDOM[10'h17B][23];	// lsu.scala:210:16
        ldq_21_bits_succeeded = _RANDOM[10'h17B][24];	// lsu.scala:210:16
        ldq_21_bits_order_fail = _RANDOM[10'h17B][25];	// lsu.scala:210:16
        ldq_21_bits_observed = _RANDOM[10'h17B][26];	// lsu.scala:210:16
        ldq_21_bits_st_dep_mask = {_RANDOM[10'h17B][31:27], _RANDOM[10'h17C][18:0]};	// lsu.scala:210:16
        ldq_21_bits_youngest_stq_idx = _RANDOM[10'h17C][23:19];	// lsu.scala:210:16
        ldq_21_bits_forward_std_val = _RANDOM[10'h17C][24];	// lsu.scala:210:16
        ldq_21_bits_forward_stq_idx = _RANDOM[10'h17C][29:25];	// lsu.scala:210:16
        ldq_22_valid = _RANDOM[10'h17E][30];	// lsu.scala:210:16
        ldq_22_bits_uop_uopc = {_RANDOM[10'h17E][31], _RANDOM[10'h17F][5:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_inst = {_RANDOM[10'h17F][31:6], _RANDOM[10'h180][5:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_debug_inst = {_RANDOM[10'h180][31:6], _RANDOM[10'h181][5:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_is_rvc = _RANDOM[10'h181][6];	// lsu.scala:210:16
        ldq_22_bits_uop_debug_pc = {_RANDOM[10'h181][31:7], _RANDOM[10'h182][14:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_iq_type = _RANDOM[10'h182][17:15];	// lsu.scala:210:16
        ldq_22_bits_uop_fu_code = _RANDOM[10'h182][27:18];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_br_type = _RANDOM[10'h182][31:28];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_op1_sel = _RANDOM[10'h183][1:0];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_op2_sel = _RANDOM[10'h183][4:2];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_imm_sel = _RANDOM[10'h183][7:5];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_op_fcn = _RANDOM[10'h183][11:8];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_fcn_dw = _RANDOM[10'h183][12];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_csr_cmd = _RANDOM[10'h183][15:13];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_is_load = _RANDOM[10'h183][16];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_is_sta = _RANDOM[10'h183][17];	// lsu.scala:210:16
        ldq_22_bits_uop_ctrl_is_std = _RANDOM[10'h183][18];	// lsu.scala:210:16
        ldq_22_bits_uop_iw_state = _RANDOM[10'h183][20:19];	// lsu.scala:210:16
        ldq_22_bits_uop_iw_p1_poisoned = _RANDOM[10'h183][21];	// lsu.scala:210:16
        ldq_22_bits_uop_iw_p2_poisoned = _RANDOM[10'h183][22];	// lsu.scala:210:16
        ldq_22_bits_uop_is_br = _RANDOM[10'h183][23];	// lsu.scala:210:16
        ldq_22_bits_uop_is_jalr = _RANDOM[10'h183][24];	// lsu.scala:210:16
        ldq_22_bits_uop_is_jal = _RANDOM[10'h183][25];	// lsu.scala:210:16
        ldq_22_bits_uop_is_sfb = _RANDOM[10'h183][26];	// lsu.scala:210:16
        ldq_22_bits_uop_br_mask = {_RANDOM[10'h183][31:27], _RANDOM[10'h184][10:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_br_tag = _RANDOM[10'h184][14:11];	// lsu.scala:210:16
        ldq_22_bits_uop_ftq_idx = _RANDOM[10'h184][19:15];	// lsu.scala:210:16
        ldq_22_bits_uop_edge_inst = _RANDOM[10'h184][20];	// lsu.scala:210:16
        ldq_22_bits_uop_pc_lob = _RANDOM[10'h184][26:21];	// lsu.scala:210:16
        ldq_22_bits_uop_taken = _RANDOM[10'h184][27];	// lsu.scala:210:16
        ldq_22_bits_uop_imm_packed = {_RANDOM[10'h184][31:28], _RANDOM[10'h185][15:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_csr_addr = _RANDOM[10'h185][27:16];	// lsu.scala:210:16
        ldq_22_bits_uop_rob_idx = {_RANDOM[10'h185][31:28], _RANDOM[10'h186][2:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_ldq_idx = _RANDOM[10'h186][7:3];	// lsu.scala:210:16
        ldq_22_bits_uop_stq_idx = _RANDOM[10'h186][12:8];	// lsu.scala:210:16
        ldq_22_bits_uop_rxq_idx = _RANDOM[10'h186][14:13];	// lsu.scala:210:16
        ldq_22_bits_uop_pdst = _RANDOM[10'h186][21:15];	// lsu.scala:210:16
        ldq_22_bits_uop_prs1 = _RANDOM[10'h186][28:22];	// lsu.scala:210:16
        ldq_22_bits_uop_prs2 = {_RANDOM[10'h186][31:29], _RANDOM[10'h187][3:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_prs3 = _RANDOM[10'h187][10:4];	// lsu.scala:210:16
        ldq_22_bits_uop_ppred = _RANDOM[10'h187][15:11];	// lsu.scala:210:16
        ldq_22_bits_uop_prs1_busy = _RANDOM[10'h187][16];	// lsu.scala:210:16
        ldq_22_bits_uop_prs2_busy = _RANDOM[10'h187][17];	// lsu.scala:210:16
        ldq_22_bits_uop_prs3_busy = _RANDOM[10'h187][18];	// lsu.scala:210:16
        ldq_22_bits_uop_ppred_busy = _RANDOM[10'h187][19];	// lsu.scala:210:16
        ldq_22_bits_uop_stale_pdst = _RANDOM[10'h187][26:20];	// lsu.scala:210:16
        ldq_22_bits_uop_exception = _RANDOM[10'h187][27];	// lsu.scala:210:16
        ldq_22_bits_uop_exc_cause =
          {_RANDOM[10'h187][31:28], _RANDOM[10'h188], _RANDOM[10'h189][27:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_bypassable = _RANDOM[10'h189][28];	// lsu.scala:210:16
        ldq_22_bits_uop_mem_cmd = {_RANDOM[10'h189][31:29], _RANDOM[10'h18A][1:0]};	// lsu.scala:210:16
        ldq_22_bits_uop_mem_size = _RANDOM[10'h18A][3:2];	// lsu.scala:210:16
        ldq_22_bits_uop_mem_signed = _RANDOM[10'h18A][4];	// lsu.scala:210:16
        ldq_22_bits_uop_is_fence = _RANDOM[10'h18A][5];	// lsu.scala:210:16
        ldq_22_bits_uop_is_fencei = _RANDOM[10'h18A][6];	// lsu.scala:210:16
        ldq_22_bits_uop_is_amo = _RANDOM[10'h18A][7];	// lsu.scala:210:16
        ldq_22_bits_uop_uses_ldq = _RANDOM[10'h18A][8];	// lsu.scala:210:16
        ldq_22_bits_uop_uses_stq = _RANDOM[10'h18A][9];	// lsu.scala:210:16
        ldq_22_bits_uop_is_sys_pc2epc = _RANDOM[10'h18A][10];	// lsu.scala:210:16
        ldq_22_bits_uop_is_unique = _RANDOM[10'h18A][11];	// lsu.scala:210:16
        ldq_22_bits_uop_flush_on_commit = _RANDOM[10'h18A][12];	// lsu.scala:210:16
        ldq_22_bits_uop_ldst_is_rs1 = _RANDOM[10'h18A][13];	// lsu.scala:210:16
        ldq_22_bits_uop_ldst = _RANDOM[10'h18A][19:14];	// lsu.scala:210:16
        ldq_22_bits_uop_lrs1 = _RANDOM[10'h18A][25:20];	// lsu.scala:210:16
        ldq_22_bits_uop_lrs2 = _RANDOM[10'h18A][31:26];	// lsu.scala:210:16
        ldq_22_bits_uop_lrs3 = _RANDOM[10'h18B][5:0];	// lsu.scala:210:16
        ldq_22_bits_uop_ldst_val = _RANDOM[10'h18B][6];	// lsu.scala:210:16
        ldq_22_bits_uop_dst_rtype = _RANDOM[10'h18B][8:7];	// lsu.scala:210:16
        ldq_22_bits_uop_lrs1_rtype = _RANDOM[10'h18B][10:9];	// lsu.scala:210:16
        ldq_22_bits_uop_lrs2_rtype = _RANDOM[10'h18B][12:11];	// lsu.scala:210:16
        ldq_22_bits_uop_frs3_en = _RANDOM[10'h18B][13];	// lsu.scala:210:16
        ldq_22_bits_uop_fp_val = _RANDOM[10'h18B][14];	// lsu.scala:210:16
        ldq_22_bits_uop_fp_single = _RANDOM[10'h18B][15];	// lsu.scala:210:16
        ldq_22_bits_uop_xcpt_pf_if = _RANDOM[10'h18B][16];	// lsu.scala:210:16
        ldq_22_bits_uop_xcpt_ae_if = _RANDOM[10'h18B][17];	// lsu.scala:210:16
        ldq_22_bits_uop_xcpt_ma_if = _RANDOM[10'h18B][18];	// lsu.scala:210:16
        ldq_22_bits_uop_bp_debug_if = _RANDOM[10'h18B][19];	// lsu.scala:210:16
        ldq_22_bits_uop_bp_xcpt_if = _RANDOM[10'h18B][20];	// lsu.scala:210:16
        ldq_22_bits_uop_debug_fsrc = _RANDOM[10'h18B][22:21];	// lsu.scala:210:16
        ldq_22_bits_uop_debug_tsrc = _RANDOM[10'h18B][24:23];	// lsu.scala:210:16
        ldq_22_bits_addr_valid = _RANDOM[10'h18B][25];	// lsu.scala:210:16
        ldq_22_bits_addr_bits =
          {_RANDOM[10'h18B][31:26], _RANDOM[10'h18C], _RANDOM[10'h18D][1:0]};	// lsu.scala:210:16
        ldq_22_bits_addr_is_virtual = _RANDOM[10'h18D][2];	// lsu.scala:210:16
        ldq_22_bits_addr_is_uncacheable = _RANDOM[10'h18D][3];	// lsu.scala:210:16
        ldq_22_bits_executed = _RANDOM[10'h18D][4];	// lsu.scala:210:16
        ldq_22_bits_succeeded = _RANDOM[10'h18D][5];	// lsu.scala:210:16
        ldq_22_bits_order_fail = _RANDOM[10'h18D][6];	// lsu.scala:210:16
        ldq_22_bits_observed = _RANDOM[10'h18D][7];	// lsu.scala:210:16
        ldq_22_bits_st_dep_mask = _RANDOM[10'h18D][31:8];	// lsu.scala:210:16
        ldq_22_bits_youngest_stq_idx = _RANDOM[10'h18E][4:0];	// lsu.scala:210:16
        ldq_22_bits_forward_std_val = _RANDOM[10'h18E][5];	// lsu.scala:210:16
        ldq_22_bits_forward_stq_idx = _RANDOM[10'h18E][10:6];	// lsu.scala:210:16
        ldq_23_valid = _RANDOM[10'h190][11];	// lsu.scala:210:16
        ldq_23_bits_uop_uopc = _RANDOM[10'h190][18:12];	// lsu.scala:210:16
        ldq_23_bits_uop_inst = {_RANDOM[10'h190][31:19], _RANDOM[10'h191][18:0]};	// lsu.scala:210:16
        ldq_23_bits_uop_debug_inst = {_RANDOM[10'h191][31:19], _RANDOM[10'h192][18:0]};	// lsu.scala:210:16
        ldq_23_bits_uop_is_rvc = _RANDOM[10'h192][19];	// lsu.scala:210:16
        ldq_23_bits_uop_debug_pc = {_RANDOM[10'h192][31:20], _RANDOM[10'h193][27:0]};	// lsu.scala:210:16
        ldq_23_bits_uop_iq_type = _RANDOM[10'h193][30:28];	// lsu.scala:210:16
        ldq_23_bits_uop_fu_code = {_RANDOM[10'h193][31], _RANDOM[10'h194][8:0]};	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_br_type = _RANDOM[10'h194][12:9];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_op1_sel = _RANDOM[10'h194][14:13];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_op2_sel = _RANDOM[10'h194][17:15];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_imm_sel = _RANDOM[10'h194][20:18];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_op_fcn = _RANDOM[10'h194][24:21];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_fcn_dw = _RANDOM[10'h194][25];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_csr_cmd = _RANDOM[10'h194][28:26];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_is_load = _RANDOM[10'h194][29];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_is_sta = _RANDOM[10'h194][30];	// lsu.scala:210:16
        ldq_23_bits_uop_ctrl_is_std = _RANDOM[10'h194][31];	// lsu.scala:210:16
        ldq_23_bits_uop_iw_state = _RANDOM[10'h195][1:0];	// lsu.scala:210:16
        ldq_23_bits_uop_iw_p1_poisoned = _RANDOM[10'h195][2];	// lsu.scala:210:16
        ldq_23_bits_uop_iw_p2_poisoned = _RANDOM[10'h195][3];	// lsu.scala:210:16
        ldq_23_bits_uop_is_br = _RANDOM[10'h195][4];	// lsu.scala:210:16
        ldq_23_bits_uop_is_jalr = _RANDOM[10'h195][5];	// lsu.scala:210:16
        ldq_23_bits_uop_is_jal = _RANDOM[10'h195][6];	// lsu.scala:210:16
        ldq_23_bits_uop_is_sfb = _RANDOM[10'h195][7];	// lsu.scala:210:16
        ldq_23_bits_uop_br_mask = _RANDOM[10'h195][23:8];	// lsu.scala:210:16
        ldq_23_bits_uop_br_tag = _RANDOM[10'h195][27:24];	// lsu.scala:210:16
        ldq_23_bits_uop_ftq_idx = {_RANDOM[10'h195][31:28], _RANDOM[10'h196][0]};	// lsu.scala:210:16
        ldq_23_bits_uop_edge_inst = _RANDOM[10'h196][1];	// lsu.scala:210:16
        ldq_23_bits_uop_pc_lob = _RANDOM[10'h196][7:2];	// lsu.scala:210:16
        ldq_23_bits_uop_taken = _RANDOM[10'h196][8];	// lsu.scala:210:16
        ldq_23_bits_uop_imm_packed = _RANDOM[10'h196][28:9];	// lsu.scala:210:16
        ldq_23_bits_uop_csr_addr = {_RANDOM[10'h196][31:29], _RANDOM[10'h197][8:0]};	// lsu.scala:210:16
        ldq_23_bits_uop_rob_idx = _RANDOM[10'h197][15:9];	// lsu.scala:210:16
        ldq_23_bits_uop_ldq_idx = _RANDOM[10'h197][20:16];	// lsu.scala:210:16
        ldq_23_bits_uop_stq_idx = _RANDOM[10'h197][25:21];	// lsu.scala:210:16
        ldq_23_bits_uop_rxq_idx = _RANDOM[10'h197][27:26];	// lsu.scala:210:16
        ldq_23_bits_uop_pdst = {_RANDOM[10'h197][31:28], _RANDOM[10'h198][2:0]};	// lsu.scala:210:16
        ldq_23_bits_uop_prs1 = _RANDOM[10'h198][9:3];	// lsu.scala:210:16
        ldq_23_bits_uop_prs2 = _RANDOM[10'h198][16:10];	// lsu.scala:210:16
        ldq_23_bits_uop_prs3 = _RANDOM[10'h198][23:17];	// lsu.scala:210:16
        ldq_23_bits_uop_ppred = _RANDOM[10'h198][28:24];	// lsu.scala:210:16
        ldq_23_bits_uop_prs1_busy = _RANDOM[10'h198][29];	// lsu.scala:210:16
        ldq_23_bits_uop_prs2_busy = _RANDOM[10'h198][30];	// lsu.scala:210:16
        ldq_23_bits_uop_prs3_busy = _RANDOM[10'h198][31];	// lsu.scala:210:16
        ldq_23_bits_uop_ppred_busy = _RANDOM[10'h199][0];	// lsu.scala:210:16
        ldq_23_bits_uop_stale_pdst = _RANDOM[10'h199][7:1];	// lsu.scala:210:16
        ldq_23_bits_uop_exception = _RANDOM[10'h199][8];	// lsu.scala:210:16
        ldq_23_bits_uop_exc_cause =
          {_RANDOM[10'h199][31:9], _RANDOM[10'h19A], _RANDOM[10'h19B][8:0]};	// lsu.scala:210:16
        ldq_23_bits_uop_bypassable = _RANDOM[10'h19B][9];	// lsu.scala:210:16
        ldq_23_bits_uop_mem_cmd = _RANDOM[10'h19B][14:10];	// lsu.scala:210:16
        ldq_23_bits_uop_mem_size = _RANDOM[10'h19B][16:15];	// lsu.scala:210:16
        ldq_23_bits_uop_mem_signed = _RANDOM[10'h19B][17];	// lsu.scala:210:16
        ldq_23_bits_uop_is_fence = _RANDOM[10'h19B][18];	// lsu.scala:210:16
        ldq_23_bits_uop_is_fencei = _RANDOM[10'h19B][19];	// lsu.scala:210:16
        ldq_23_bits_uop_is_amo = _RANDOM[10'h19B][20];	// lsu.scala:210:16
        ldq_23_bits_uop_uses_ldq = _RANDOM[10'h19B][21];	// lsu.scala:210:16
        ldq_23_bits_uop_uses_stq = _RANDOM[10'h19B][22];	// lsu.scala:210:16
        ldq_23_bits_uop_is_sys_pc2epc = _RANDOM[10'h19B][23];	// lsu.scala:210:16
        ldq_23_bits_uop_is_unique = _RANDOM[10'h19B][24];	// lsu.scala:210:16
        ldq_23_bits_uop_flush_on_commit = _RANDOM[10'h19B][25];	// lsu.scala:210:16
        ldq_23_bits_uop_ldst_is_rs1 = _RANDOM[10'h19B][26];	// lsu.scala:210:16
        ldq_23_bits_uop_ldst = {_RANDOM[10'h19B][31:27], _RANDOM[10'h19C][0]};	// lsu.scala:210:16
        ldq_23_bits_uop_lrs1 = _RANDOM[10'h19C][6:1];	// lsu.scala:210:16
        ldq_23_bits_uop_lrs2 = _RANDOM[10'h19C][12:7];	// lsu.scala:210:16
        ldq_23_bits_uop_lrs3 = _RANDOM[10'h19C][18:13];	// lsu.scala:210:16
        ldq_23_bits_uop_ldst_val = _RANDOM[10'h19C][19];	// lsu.scala:210:16
        ldq_23_bits_uop_dst_rtype = _RANDOM[10'h19C][21:20];	// lsu.scala:210:16
        ldq_23_bits_uop_lrs1_rtype = _RANDOM[10'h19C][23:22];	// lsu.scala:210:16
        ldq_23_bits_uop_lrs2_rtype = _RANDOM[10'h19C][25:24];	// lsu.scala:210:16
        ldq_23_bits_uop_frs3_en = _RANDOM[10'h19C][26];	// lsu.scala:210:16
        ldq_23_bits_uop_fp_val = _RANDOM[10'h19C][27];	// lsu.scala:210:16
        ldq_23_bits_uop_fp_single = _RANDOM[10'h19C][28];	// lsu.scala:210:16
        ldq_23_bits_uop_xcpt_pf_if = _RANDOM[10'h19C][29];	// lsu.scala:210:16
        ldq_23_bits_uop_xcpt_ae_if = _RANDOM[10'h19C][30];	// lsu.scala:210:16
        ldq_23_bits_uop_xcpt_ma_if = _RANDOM[10'h19C][31];	// lsu.scala:210:16
        ldq_23_bits_uop_bp_debug_if = _RANDOM[10'h19D][0];	// lsu.scala:210:16
        ldq_23_bits_uop_bp_xcpt_if = _RANDOM[10'h19D][1];	// lsu.scala:210:16
        ldq_23_bits_uop_debug_fsrc = _RANDOM[10'h19D][3:2];	// lsu.scala:210:16
        ldq_23_bits_uop_debug_tsrc = _RANDOM[10'h19D][5:4];	// lsu.scala:210:16
        ldq_23_bits_addr_valid = _RANDOM[10'h19D][6];	// lsu.scala:210:16
        ldq_23_bits_addr_bits = {_RANDOM[10'h19D][31:7], _RANDOM[10'h19E][14:0]};	// lsu.scala:210:16
        ldq_23_bits_addr_is_virtual = _RANDOM[10'h19E][15];	// lsu.scala:210:16
        ldq_23_bits_addr_is_uncacheable = _RANDOM[10'h19E][16];	// lsu.scala:210:16
        ldq_23_bits_executed = _RANDOM[10'h19E][17];	// lsu.scala:210:16
        ldq_23_bits_succeeded = _RANDOM[10'h19E][18];	// lsu.scala:210:16
        ldq_23_bits_order_fail = _RANDOM[10'h19E][19];	// lsu.scala:210:16
        ldq_23_bits_observed = _RANDOM[10'h19E][20];	// lsu.scala:210:16
        ldq_23_bits_st_dep_mask = {_RANDOM[10'h19E][31:21], _RANDOM[10'h19F][12:0]};	// lsu.scala:210:16
        ldq_23_bits_youngest_stq_idx = _RANDOM[10'h19F][17:13];	// lsu.scala:210:16
        ldq_23_bits_forward_std_val = _RANDOM[10'h19F][18];	// lsu.scala:210:16
        ldq_23_bits_forward_stq_idx = _RANDOM[10'h19F][23:19];	// lsu.scala:210:16
        stq_0_valid = _RANDOM[10'h1A1][24];	// lsu.scala:211:16
        stq_0_bits_uop_uopc = _RANDOM[10'h1A1][31:25];	// lsu.scala:211:16
        stq_0_bits_uop_inst = _RANDOM[10'h1A2];	// lsu.scala:211:16
        stq_0_bits_uop_debug_inst = _RANDOM[10'h1A3];	// lsu.scala:211:16
        stq_0_bits_uop_is_rvc = _RANDOM[10'h1A4][0];	// lsu.scala:211:16
        stq_0_bits_uop_debug_pc = {_RANDOM[10'h1A4][31:1], _RANDOM[10'h1A5][8:0]};	// lsu.scala:211:16
        stq_0_bits_uop_iq_type = _RANDOM[10'h1A5][11:9];	// lsu.scala:211:16
        stq_0_bits_uop_fu_code = _RANDOM[10'h1A5][21:12];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_br_type = _RANDOM[10'h1A5][25:22];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op1_sel = _RANDOM[10'h1A5][27:26];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op2_sel = _RANDOM[10'h1A5][30:28];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_imm_sel = {_RANDOM[10'h1A5][31], _RANDOM[10'h1A6][1:0]};	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op_fcn = _RANDOM[10'h1A6][5:2];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1A6][6];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1A6][9:7];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_is_load = _RANDOM[10'h1A6][10];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_is_sta = _RANDOM[10'h1A6][11];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_is_std = _RANDOM[10'h1A6][12];	// lsu.scala:211:16
        stq_0_bits_uop_iw_state = _RANDOM[10'h1A6][14:13];	// lsu.scala:211:16
        stq_0_bits_uop_iw_p1_poisoned = _RANDOM[10'h1A6][15];	// lsu.scala:211:16
        stq_0_bits_uop_iw_p2_poisoned = _RANDOM[10'h1A6][16];	// lsu.scala:211:16
        stq_0_bits_uop_is_br = _RANDOM[10'h1A6][17];	// lsu.scala:211:16
        stq_0_bits_uop_is_jalr = _RANDOM[10'h1A6][18];	// lsu.scala:211:16
        stq_0_bits_uop_is_jal = _RANDOM[10'h1A6][19];	// lsu.scala:211:16
        stq_0_bits_uop_is_sfb = _RANDOM[10'h1A6][20];	// lsu.scala:211:16
        stq_0_bits_uop_br_mask = {_RANDOM[10'h1A6][31:21], _RANDOM[10'h1A7][4:0]};	// lsu.scala:211:16
        stq_0_bits_uop_br_tag = _RANDOM[10'h1A7][8:5];	// lsu.scala:211:16
        stq_0_bits_uop_ftq_idx = _RANDOM[10'h1A7][13:9];	// lsu.scala:211:16
        stq_0_bits_uop_edge_inst = _RANDOM[10'h1A7][14];	// lsu.scala:211:16
        stq_0_bits_uop_pc_lob = _RANDOM[10'h1A7][20:15];	// lsu.scala:211:16
        stq_0_bits_uop_taken = _RANDOM[10'h1A7][21];	// lsu.scala:211:16
        stq_0_bits_uop_imm_packed = {_RANDOM[10'h1A7][31:22], _RANDOM[10'h1A8][9:0]};	// lsu.scala:211:16
        stq_0_bits_uop_csr_addr = _RANDOM[10'h1A8][21:10];	// lsu.scala:211:16
        stq_0_bits_uop_rob_idx = _RANDOM[10'h1A8][28:22];	// lsu.scala:211:16
        stq_0_bits_uop_ldq_idx = {_RANDOM[10'h1A8][31:29], _RANDOM[10'h1A9][1:0]};	// lsu.scala:211:16
        stq_0_bits_uop_stq_idx = _RANDOM[10'h1A9][6:2];	// lsu.scala:211:16
        stq_0_bits_uop_rxq_idx = _RANDOM[10'h1A9][8:7];	// lsu.scala:211:16
        stq_0_bits_uop_pdst = _RANDOM[10'h1A9][15:9];	// lsu.scala:211:16
        stq_0_bits_uop_prs1 = _RANDOM[10'h1A9][22:16];	// lsu.scala:211:16
        stq_0_bits_uop_prs2 = _RANDOM[10'h1A9][29:23];	// lsu.scala:211:16
        stq_0_bits_uop_prs3 = {_RANDOM[10'h1A9][31:30], _RANDOM[10'h1AA][4:0]};	// lsu.scala:211:16
        stq_0_bits_uop_ppred = _RANDOM[10'h1AA][9:5];	// lsu.scala:211:16
        stq_0_bits_uop_prs1_busy = _RANDOM[10'h1AA][10];	// lsu.scala:211:16
        stq_0_bits_uop_prs2_busy = _RANDOM[10'h1AA][11];	// lsu.scala:211:16
        stq_0_bits_uop_prs3_busy = _RANDOM[10'h1AA][12];	// lsu.scala:211:16
        stq_0_bits_uop_ppred_busy = _RANDOM[10'h1AA][13];	// lsu.scala:211:16
        stq_0_bits_uop_stale_pdst = _RANDOM[10'h1AA][20:14];	// lsu.scala:211:16
        stq_0_bits_uop_exception = _RANDOM[10'h1AA][21];	// lsu.scala:211:16
        stq_0_bits_uop_exc_cause =
          {_RANDOM[10'h1AA][31:22], _RANDOM[10'h1AB], _RANDOM[10'h1AC][21:0]};	// lsu.scala:211:16
        stq_0_bits_uop_bypassable = _RANDOM[10'h1AC][22];	// lsu.scala:211:16
        stq_0_bits_uop_mem_cmd = _RANDOM[10'h1AC][27:23];	// lsu.scala:211:16
        stq_0_bits_uop_mem_size = _RANDOM[10'h1AC][29:28];	// lsu.scala:211:16
        stq_0_bits_uop_mem_signed = _RANDOM[10'h1AC][30];	// lsu.scala:211:16
        stq_0_bits_uop_is_fence = _RANDOM[10'h1AC][31];	// lsu.scala:211:16
        stq_0_bits_uop_is_fencei = _RANDOM[10'h1AD][0];	// lsu.scala:211:16
        stq_0_bits_uop_is_amo = _RANDOM[10'h1AD][1];	// lsu.scala:211:16
        stq_0_bits_uop_uses_ldq = _RANDOM[10'h1AD][2];	// lsu.scala:211:16
        stq_0_bits_uop_uses_stq = _RANDOM[10'h1AD][3];	// lsu.scala:211:16
        stq_0_bits_uop_is_sys_pc2epc = _RANDOM[10'h1AD][4];	// lsu.scala:211:16
        stq_0_bits_uop_is_unique = _RANDOM[10'h1AD][5];	// lsu.scala:211:16
        stq_0_bits_uop_flush_on_commit = _RANDOM[10'h1AD][6];	// lsu.scala:211:16
        stq_0_bits_uop_ldst_is_rs1 = _RANDOM[10'h1AD][7];	// lsu.scala:211:16
        stq_0_bits_uop_ldst = _RANDOM[10'h1AD][13:8];	// lsu.scala:211:16
        stq_0_bits_uop_lrs1 = _RANDOM[10'h1AD][19:14];	// lsu.scala:211:16
        stq_0_bits_uop_lrs2 = _RANDOM[10'h1AD][25:20];	// lsu.scala:211:16
        stq_0_bits_uop_lrs3 = _RANDOM[10'h1AD][31:26];	// lsu.scala:211:16
        stq_0_bits_uop_ldst_val = _RANDOM[10'h1AE][0];	// lsu.scala:211:16
        stq_0_bits_uop_dst_rtype = _RANDOM[10'h1AE][2:1];	// lsu.scala:211:16
        stq_0_bits_uop_lrs1_rtype = _RANDOM[10'h1AE][4:3];	// lsu.scala:211:16
        stq_0_bits_uop_lrs2_rtype = _RANDOM[10'h1AE][6:5];	// lsu.scala:211:16
        stq_0_bits_uop_frs3_en = _RANDOM[10'h1AE][7];	// lsu.scala:211:16
        stq_0_bits_uop_fp_val = _RANDOM[10'h1AE][8];	// lsu.scala:211:16
        stq_0_bits_uop_fp_single = _RANDOM[10'h1AE][9];	// lsu.scala:211:16
        stq_0_bits_uop_xcpt_pf_if = _RANDOM[10'h1AE][10];	// lsu.scala:211:16
        stq_0_bits_uop_xcpt_ae_if = _RANDOM[10'h1AE][11];	// lsu.scala:211:16
        stq_0_bits_uop_xcpt_ma_if = _RANDOM[10'h1AE][12];	// lsu.scala:211:16
        stq_0_bits_uop_bp_debug_if = _RANDOM[10'h1AE][13];	// lsu.scala:211:16
        stq_0_bits_uop_bp_xcpt_if = _RANDOM[10'h1AE][14];	// lsu.scala:211:16
        stq_0_bits_uop_debug_fsrc = _RANDOM[10'h1AE][16:15];	// lsu.scala:211:16
        stq_0_bits_uop_debug_tsrc = _RANDOM[10'h1AE][18:17];	// lsu.scala:211:16
        stq_0_bits_addr_valid = _RANDOM[10'h1AE][19];	// lsu.scala:211:16
        stq_0_bits_addr_bits = {_RANDOM[10'h1AE][31:20], _RANDOM[10'h1AF][27:0]};	// lsu.scala:211:16
        stq_0_bits_addr_is_virtual = _RANDOM[10'h1AF][28];	// lsu.scala:211:16
        stq_0_bits_data_valid = _RANDOM[10'h1AF][29];	// lsu.scala:211:16
        stq_0_bits_data_bits =
          {_RANDOM[10'h1AF][31:30], _RANDOM[10'h1B0], _RANDOM[10'h1B1][29:0]};	// lsu.scala:211:16
        stq_0_bits_committed = _RANDOM[10'h1B1][30];	// lsu.scala:211:16
        stq_0_bits_succeeded = _RANDOM[10'h1B1][31];	// lsu.scala:211:16
        stq_1_valid = _RANDOM[10'h1B4][0];	// lsu.scala:211:16
        stq_1_bits_uop_uopc = _RANDOM[10'h1B4][7:1];	// lsu.scala:211:16
        stq_1_bits_uop_inst = {_RANDOM[10'h1B4][31:8], _RANDOM[10'h1B5][7:0]};	// lsu.scala:211:16
        stq_1_bits_uop_debug_inst = {_RANDOM[10'h1B5][31:8], _RANDOM[10'h1B6][7:0]};	// lsu.scala:211:16
        stq_1_bits_uop_is_rvc = _RANDOM[10'h1B6][8];	// lsu.scala:211:16
        stq_1_bits_uop_debug_pc = {_RANDOM[10'h1B6][31:9], _RANDOM[10'h1B7][16:0]};	// lsu.scala:211:16
        stq_1_bits_uop_iq_type = _RANDOM[10'h1B7][19:17];	// lsu.scala:211:16
        stq_1_bits_uop_fu_code = _RANDOM[10'h1B7][29:20];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_br_type = {_RANDOM[10'h1B7][31:30], _RANDOM[10'h1B8][1:0]};	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op1_sel = _RANDOM[10'h1B8][3:2];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op2_sel = _RANDOM[10'h1B8][6:4];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_imm_sel = _RANDOM[10'h1B8][9:7];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op_fcn = _RANDOM[10'h1B8][13:10];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1B8][14];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1B8][17:15];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_is_load = _RANDOM[10'h1B8][18];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_is_sta = _RANDOM[10'h1B8][19];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_is_std = _RANDOM[10'h1B8][20];	// lsu.scala:211:16
        stq_1_bits_uop_iw_state = _RANDOM[10'h1B8][22:21];	// lsu.scala:211:16
        stq_1_bits_uop_iw_p1_poisoned = _RANDOM[10'h1B8][23];	// lsu.scala:211:16
        stq_1_bits_uop_iw_p2_poisoned = _RANDOM[10'h1B8][24];	// lsu.scala:211:16
        stq_1_bits_uop_is_br = _RANDOM[10'h1B8][25];	// lsu.scala:211:16
        stq_1_bits_uop_is_jalr = _RANDOM[10'h1B8][26];	// lsu.scala:211:16
        stq_1_bits_uop_is_jal = _RANDOM[10'h1B8][27];	// lsu.scala:211:16
        stq_1_bits_uop_is_sfb = _RANDOM[10'h1B8][28];	// lsu.scala:211:16
        stq_1_bits_uop_br_mask = {_RANDOM[10'h1B8][31:29], _RANDOM[10'h1B9][12:0]};	// lsu.scala:211:16
        stq_1_bits_uop_br_tag = _RANDOM[10'h1B9][16:13];	// lsu.scala:211:16
        stq_1_bits_uop_ftq_idx = _RANDOM[10'h1B9][21:17];	// lsu.scala:211:16
        stq_1_bits_uop_edge_inst = _RANDOM[10'h1B9][22];	// lsu.scala:211:16
        stq_1_bits_uop_pc_lob = _RANDOM[10'h1B9][28:23];	// lsu.scala:211:16
        stq_1_bits_uop_taken = _RANDOM[10'h1B9][29];	// lsu.scala:211:16
        stq_1_bits_uop_imm_packed = {_RANDOM[10'h1B9][31:30], _RANDOM[10'h1BA][17:0]};	// lsu.scala:211:16
        stq_1_bits_uop_csr_addr = _RANDOM[10'h1BA][29:18];	// lsu.scala:211:16
        stq_1_bits_uop_rob_idx = {_RANDOM[10'h1BA][31:30], _RANDOM[10'h1BB][4:0]};	// lsu.scala:211:16
        stq_1_bits_uop_ldq_idx = _RANDOM[10'h1BB][9:5];	// lsu.scala:211:16
        stq_1_bits_uop_stq_idx = _RANDOM[10'h1BB][14:10];	// lsu.scala:211:16
        stq_1_bits_uop_rxq_idx = _RANDOM[10'h1BB][16:15];	// lsu.scala:211:16
        stq_1_bits_uop_pdst = _RANDOM[10'h1BB][23:17];	// lsu.scala:211:16
        stq_1_bits_uop_prs1 = _RANDOM[10'h1BB][30:24];	// lsu.scala:211:16
        stq_1_bits_uop_prs2 = {_RANDOM[10'h1BB][31], _RANDOM[10'h1BC][5:0]};	// lsu.scala:211:16
        stq_1_bits_uop_prs3 = _RANDOM[10'h1BC][12:6];	// lsu.scala:211:16
        stq_1_bits_uop_ppred = _RANDOM[10'h1BC][17:13];	// lsu.scala:211:16
        stq_1_bits_uop_prs1_busy = _RANDOM[10'h1BC][18];	// lsu.scala:211:16
        stq_1_bits_uop_prs2_busy = _RANDOM[10'h1BC][19];	// lsu.scala:211:16
        stq_1_bits_uop_prs3_busy = _RANDOM[10'h1BC][20];	// lsu.scala:211:16
        stq_1_bits_uop_ppred_busy = _RANDOM[10'h1BC][21];	// lsu.scala:211:16
        stq_1_bits_uop_stale_pdst = _RANDOM[10'h1BC][28:22];	// lsu.scala:211:16
        stq_1_bits_uop_exception = _RANDOM[10'h1BC][29];	// lsu.scala:211:16
        stq_1_bits_uop_exc_cause =
          {_RANDOM[10'h1BC][31:30], _RANDOM[10'h1BD], _RANDOM[10'h1BE][29:0]};	// lsu.scala:211:16
        stq_1_bits_uop_bypassable = _RANDOM[10'h1BE][30];	// lsu.scala:211:16
        stq_1_bits_uop_mem_cmd = {_RANDOM[10'h1BE][31], _RANDOM[10'h1BF][3:0]};	// lsu.scala:211:16
        stq_1_bits_uop_mem_size = _RANDOM[10'h1BF][5:4];	// lsu.scala:211:16
        stq_1_bits_uop_mem_signed = _RANDOM[10'h1BF][6];	// lsu.scala:211:16
        stq_1_bits_uop_is_fence = _RANDOM[10'h1BF][7];	// lsu.scala:211:16
        stq_1_bits_uop_is_fencei = _RANDOM[10'h1BF][8];	// lsu.scala:211:16
        stq_1_bits_uop_is_amo = _RANDOM[10'h1BF][9];	// lsu.scala:211:16
        stq_1_bits_uop_uses_ldq = _RANDOM[10'h1BF][10];	// lsu.scala:211:16
        stq_1_bits_uop_uses_stq = _RANDOM[10'h1BF][11];	// lsu.scala:211:16
        stq_1_bits_uop_is_sys_pc2epc = _RANDOM[10'h1BF][12];	// lsu.scala:211:16
        stq_1_bits_uop_is_unique = _RANDOM[10'h1BF][13];	// lsu.scala:211:16
        stq_1_bits_uop_flush_on_commit = _RANDOM[10'h1BF][14];	// lsu.scala:211:16
        stq_1_bits_uop_ldst_is_rs1 = _RANDOM[10'h1BF][15];	// lsu.scala:211:16
        stq_1_bits_uop_ldst = _RANDOM[10'h1BF][21:16];	// lsu.scala:211:16
        stq_1_bits_uop_lrs1 = _RANDOM[10'h1BF][27:22];	// lsu.scala:211:16
        stq_1_bits_uop_lrs2 = {_RANDOM[10'h1BF][31:28], _RANDOM[10'h1C0][1:0]};	// lsu.scala:211:16
        stq_1_bits_uop_lrs3 = _RANDOM[10'h1C0][7:2];	// lsu.scala:211:16
        stq_1_bits_uop_ldst_val = _RANDOM[10'h1C0][8];	// lsu.scala:211:16
        stq_1_bits_uop_dst_rtype = _RANDOM[10'h1C0][10:9];	// lsu.scala:211:16
        stq_1_bits_uop_lrs1_rtype = _RANDOM[10'h1C0][12:11];	// lsu.scala:211:16
        stq_1_bits_uop_lrs2_rtype = _RANDOM[10'h1C0][14:13];	// lsu.scala:211:16
        stq_1_bits_uop_frs3_en = _RANDOM[10'h1C0][15];	// lsu.scala:211:16
        stq_1_bits_uop_fp_val = _RANDOM[10'h1C0][16];	// lsu.scala:211:16
        stq_1_bits_uop_fp_single = _RANDOM[10'h1C0][17];	// lsu.scala:211:16
        stq_1_bits_uop_xcpt_pf_if = _RANDOM[10'h1C0][18];	// lsu.scala:211:16
        stq_1_bits_uop_xcpt_ae_if = _RANDOM[10'h1C0][19];	// lsu.scala:211:16
        stq_1_bits_uop_xcpt_ma_if = _RANDOM[10'h1C0][20];	// lsu.scala:211:16
        stq_1_bits_uop_bp_debug_if = _RANDOM[10'h1C0][21];	// lsu.scala:211:16
        stq_1_bits_uop_bp_xcpt_if = _RANDOM[10'h1C0][22];	// lsu.scala:211:16
        stq_1_bits_uop_debug_fsrc = _RANDOM[10'h1C0][24:23];	// lsu.scala:211:16
        stq_1_bits_uop_debug_tsrc = _RANDOM[10'h1C0][26:25];	// lsu.scala:211:16
        stq_1_bits_addr_valid = _RANDOM[10'h1C0][27];	// lsu.scala:211:16
        stq_1_bits_addr_bits =
          {_RANDOM[10'h1C0][31:28], _RANDOM[10'h1C1], _RANDOM[10'h1C2][3:0]};	// lsu.scala:211:16
        stq_1_bits_addr_is_virtual = _RANDOM[10'h1C2][4];	// lsu.scala:211:16
        stq_1_bits_data_valid = _RANDOM[10'h1C2][5];	// lsu.scala:211:16
        stq_1_bits_data_bits =
          {_RANDOM[10'h1C2][31:6], _RANDOM[10'h1C3], _RANDOM[10'h1C4][5:0]};	// lsu.scala:211:16
        stq_1_bits_committed = _RANDOM[10'h1C4][6];	// lsu.scala:211:16
        stq_1_bits_succeeded = _RANDOM[10'h1C4][7];	// lsu.scala:211:16
        stq_2_valid = _RANDOM[10'h1C6][8];	// lsu.scala:211:16
        stq_2_bits_uop_uopc = _RANDOM[10'h1C6][15:9];	// lsu.scala:211:16
        stq_2_bits_uop_inst = {_RANDOM[10'h1C6][31:16], _RANDOM[10'h1C7][15:0]};	// lsu.scala:211:16
        stq_2_bits_uop_debug_inst = {_RANDOM[10'h1C7][31:16], _RANDOM[10'h1C8][15:0]};	// lsu.scala:211:16
        stq_2_bits_uop_is_rvc = _RANDOM[10'h1C8][16];	// lsu.scala:211:16
        stq_2_bits_uop_debug_pc = {_RANDOM[10'h1C8][31:17], _RANDOM[10'h1C9][24:0]};	// lsu.scala:211:16
        stq_2_bits_uop_iq_type = _RANDOM[10'h1C9][27:25];	// lsu.scala:211:16
        stq_2_bits_uop_fu_code = {_RANDOM[10'h1C9][31:28], _RANDOM[10'h1CA][5:0]};	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_br_type = _RANDOM[10'h1CA][9:6];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op1_sel = _RANDOM[10'h1CA][11:10];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op2_sel = _RANDOM[10'h1CA][14:12];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_imm_sel = _RANDOM[10'h1CA][17:15];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op_fcn = _RANDOM[10'h1CA][21:18];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1CA][22];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1CA][25:23];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_is_load = _RANDOM[10'h1CA][26];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_is_sta = _RANDOM[10'h1CA][27];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_is_std = _RANDOM[10'h1CA][28];	// lsu.scala:211:16
        stq_2_bits_uop_iw_state = _RANDOM[10'h1CA][30:29];	// lsu.scala:211:16
        stq_2_bits_uop_iw_p1_poisoned = _RANDOM[10'h1CA][31];	// lsu.scala:211:16
        stq_2_bits_uop_iw_p2_poisoned = _RANDOM[10'h1CB][0];	// lsu.scala:211:16
        stq_2_bits_uop_is_br = _RANDOM[10'h1CB][1];	// lsu.scala:211:16
        stq_2_bits_uop_is_jalr = _RANDOM[10'h1CB][2];	// lsu.scala:211:16
        stq_2_bits_uop_is_jal = _RANDOM[10'h1CB][3];	// lsu.scala:211:16
        stq_2_bits_uop_is_sfb = _RANDOM[10'h1CB][4];	// lsu.scala:211:16
        stq_2_bits_uop_br_mask = _RANDOM[10'h1CB][20:5];	// lsu.scala:211:16
        stq_2_bits_uop_br_tag = _RANDOM[10'h1CB][24:21];	// lsu.scala:211:16
        stq_2_bits_uop_ftq_idx = _RANDOM[10'h1CB][29:25];	// lsu.scala:211:16
        stq_2_bits_uop_edge_inst = _RANDOM[10'h1CB][30];	// lsu.scala:211:16
        stq_2_bits_uop_pc_lob = {_RANDOM[10'h1CB][31], _RANDOM[10'h1CC][4:0]};	// lsu.scala:211:16
        stq_2_bits_uop_taken = _RANDOM[10'h1CC][5];	// lsu.scala:211:16
        stq_2_bits_uop_imm_packed = _RANDOM[10'h1CC][25:6];	// lsu.scala:211:16
        stq_2_bits_uop_csr_addr = {_RANDOM[10'h1CC][31:26], _RANDOM[10'h1CD][5:0]};	// lsu.scala:211:16
        stq_2_bits_uop_rob_idx = _RANDOM[10'h1CD][12:6];	// lsu.scala:211:16
        stq_2_bits_uop_ldq_idx = _RANDOM[10'h1CD][17:13];	// lsu.scala:211:16
        stq_2_bits_uop_stq_idx = _RANDOM[10'h1CD][22:18];	// lsu.scala:211:16
        stq_2_bits_uop_rxq_idx = _RANDOM[10'h1CD][24:23];	// lsu.scala:211:16
        stq_2_bits_uop_pdst = _RANDOM[10'h1CD][31:25];	// lsu.scala:211:16
        stq_2_bits_uop_prs1 = _RANDOM[10'h1CE][6:0];	// lsu.scala:211:16
        stq_2_bits_uop_prs2 = _RANDOM[10'h1CE][13:7];	// lsu.scala:211:16
        stq_2_bits_uop_prs3 = _RANDOM[10'h1CE][20:14];	// lsu.scala:211:16
        stq_2_bits_uop_ppred = _RANDOM[10'h1CE][25:21];	// lsu.scala:211:16
        stq_2_bits_uop_prs1_busy = _RANDOM[10'h1CE][26];	// lsu.scala:211:16
        stq_2_bits_uop_prs2_busy = _RANDOM[10'h1CE][27];	// lsu.scala:211:16
        stq_2_bits_uop_prs3_busy = _RANDOM[10'h1CE][28];	// lsu.scala:211:16
        stq_2_bits_uop_ppred_busy = _RANDOM[10'h1CE][29];	// lsu.scala:211:16
        stq_2_bits_uop_stale_pdst = {_RANDOM[10'h1CE][31:30], _RANDOM[10'h1CF][4:0]};	// lsu.scala:211:16
        stq_2_bits_uop_exception = _RANDOM[10'h1CF][5];	// lsu.scala:211:16
        stq_2_bits_uop_exc_cause =
          {_RANDOM[10'h1CF][31:6], _RANDOM[10'h1D0], _RANDOM[10'h1D1][5:0]};	// lsu.scala:211:16
        stq_2_bits_uop_bypassable = _RANDOM[10'h1D1][6];	// lsu.scala:211:16
        stq_2_bits_uop_mem_cmd = _RANDOM[10'h1D1][11:7];	// lsu.scala:211:16
        stq_2_bits_uop_mem_size = _RANDOM[10'h1D1][13:12];	// lsu.scala:211:16
        stq_2_bits_uop_mem_signed = _RANDOM[10'h1D1][14];	// lsu.scala:211:16
        stq_2_bits_uop_is_fence = _RANDOM[10'h1D1][15];	// lsu.scala:211:16
        stq_2_bits_uop_is_fencei = _RANDOM[10'h1D1][16];	// lsu.scala:211:16
        stq_2_bits_uop_is_amo = _RANDOM[10'h1D1][17];	// lsu.scala:211:16
        stq_2_bits_uop_uses_ldq = _RANDOM[10'h1D1][18];	// lsu.scala:211:16
        stq_2_bits_uop_uses_stq = _RANDOM[10'h1D1][19];	// lsu.scala:211:16
        stq_2_bits_uop_is_sys_pc2epc = _RANDOM[10'h1D1][20];	// lsu.scala:211:16
        stq_2_bits_uop_is_unique = _RANDOM[10'h1D1][21];	// lsu.scala:211:16
        stq_2_bits_uop_flush_on_commit = _RANDOM[10'h1D1][22];	// lsu.scala:211:16
        stq_2_bits_uop_ldst_is_rs1 = _RANDOM[10'h1D1][23];	// lsu.scala:211:16
        stq_2_bits_uop_ldst = _RANDOM[10'h1D1][29:24];	// lsu.scala:211:16
        stq_2_bits_uop_lrs1 = {_RANDOM[10'h1D1][31:30], _RANDOM[10'h1D2][3:0]};	// lsu.scala:211:16
        stq_2_bits_uop_lrs2 = _RANDOM[10'h1D2][9:4];	// lsu.scala:211:16
        stq_2_bits_uop_lrs3 = _RANDOM[10'h1D2][15:10];	// lsu.scala:211:16
        stq_2_bits_uop_ldst_val = _RANDOM[10'h1D2][16];	// lsu.scala:211:16
        stq_2_bits_uop_dst_rtype = _RANDOM[10'h1D2][18:17];	// lsu.scala:211:16
        stq_2_bits_uop_lrs1_rtype = _RANDOM[10'h1D2][20:19];	// lsu.scala:211:16
        stq_2_bits_uop_lrs2_rtype = _RANDOM[10'h1D2][22:21];	// lsu.scala:211:16
        stq_2_bits_uop_frs3_en = _RANDOM[10'h1D2][23];	// lsu.scala:211:16
        stq_2_bits_uop_fp_val = _RANDOM[10'h1D2][24];	// lsu.scala:211:16
        stq_2_bits_uop_fp_single = _RANDOM[10'h1D2][25];	// lsu.scala:211:16
        stq_2_bits_uop_xcpt_pf_if = _RANDOM[10'h1D2][26];	// lsu.scala:211:16
        stq_2_bits_uop_xcpt_ae_if = _RANDOM[10'h1D2][27];	// lsu.scala:211:16
        stq_2_bits_uop_xcpt_ma_if = _RANDOM[10'h1D2][28];	// lsu.scala:211:16
        stq_2_bits_uop_bp_debug_if = _RANDOM[10'h1D2][29];	// lsu.scala:211:16
        stq_2_bits_uop_bp_xcpt_if = _RANDOM[10'h1D2][30];	// lsu.scala:211:16
        stq_2_bits_uop_debug_fsrc = {_RANDOM[10'h1D2][31], _RANDOM[10'h1D3][0]};	// lsu.scala:211:16
        stq_2_bits_uop_debug_tsrc = _RANDOM[10'h1D3][2:1];	// lsu.scala:211:16
        stq_2_bits_addr_valid = _RANDOM[10'h1D3][3];	// lsu.scala:211:16
        stq_2_bits_addr_bits = {_RANDOM[10'h1D3][31:4], _RANDOM[10'h1D4][11:0]};	// lsu.scala:211:16
        stq_2_bits_addr_is_virtual = _RANDOM[10'h1D4][12];	// lsu.scala:211:16
        stq_2_bits_data_valid = _RANDOM[10'h1D4][13];	// lsu.scala:211:16
        stq_2_bits_data_bits =
          {_RANDOM[10'h1D4][31:14], _RANDOM[10'h1D5], _RANDOM[10'h1D6][13:0]};	// lsu.scala:211:16
        stq_2_bits_committed = _RANDOM[10'h1D6][14];	// lsu.scala:211:16
        stq_2_bits_succeeded = _RANDOM[10'h1D6][15];	// lsu.scala:211:16
        stq_3_valid = _RANDOM[10'h1D8][16];	// lsu.scala:211:16
        stq_3_bits_uop_uopc = _RANDOM[10'h1D8][23:17];	// lsu.scala:211:16
        stq_3_bits_uop_inst = {_RANDOM[10'h1D8][31:24], _RANDOM[10'h1D9][23:0]};	// lsu.scala:211:16
        stq_3_bits_uop_debug_inst = {_RANDOM[10'h1D9][31:24], _RANDOM[10'h1DA][23:0]};	// lsu.scala:211:16
        stq_3_bits_uop_is_rvc = _RANDOM[10'h1DA][24];	// lsu.scala:211:16
        stq_3_bits_uop_debug_pc =
          {_RANDOM[10'h1DA][31:25], _RANDOM[10'h1DB], _RANDOM[10'h1DC][0]};	// lsu.scala:211:16
        stq_3_bits_uop_iq_type = _RANDOM[10'h1DC][3:1];	// lsu.scala:211:16
        stq_3_bits_uop_fu_code = _RANDOM[10'h1DC][13:4];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_br_type = _RANDOM[10'h1DC][17:14];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op1_sel = _RANDOM[10'h1DC][19:18];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op2_sel = _RANDOM[10'h1DC][22:20];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_imm_sel = _RANDOM[10'h1DC][25:23];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op_fcn = _RANDOM[10'h1DC][29:26];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1DC][30];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h1DC][31], _RANDOM[10'h1DD][1:0]};	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_is_load = _RANDOM[10'h1DD][2];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_is_sta = _RANDOM[10'h1DD][3];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_is_std = _RANDOM[10'h1DD][4];	// lsu.scala:211:16
        stq_3_bits_uop_iw_state = _RANDOM[10'h1DD][6:5];	// lsu.scala:211:16
        stq_3_bits_uop_iw_p1_poisoned = _RANDOM[10'h1DD][7];	// lsu.scala:211:16
        stq_3_bits_uop_iw_p2_poisoned = _RANDOM[10'h1DD][8];	// lsu.scala:211:16
        stq_3_bits_uop_is_br = _RANDOM[10'h1DD][9];	// lsu.scala:211:16
        stq_3_bits_uop_is_jalr = _RANDOM[10'h1DD][10];	// lsu.scala:211:16
        stq_3_bits_uop_is_jal = _RANDOM[10'h1DD][11];	// lsu.scala:211:16
        stq_3_bits_uop_is_sfb = _RANDOM[10'h1DD][12];	// lsu.scala:211:16
        stq_3_bits_uop_br_mask = _RANDOM[10'h1DD][28:13];	// lsu.scala:211:16
        stq_3_bits_uop_br_tag = {_RANDOM[10'h1DD][31:29], _RANDOM[10'h1DE][0]};	// lsu.scala:211:16
        stq_3_bits_uop_ftq_idx = _RANDOM[10'h1DE][5:1];	// lsu.scala:211:16
        stq_3_bits_uop_edge_inst = _RANDOM[10'h1DE][6];	// lsu.scala:211:16
        stq_3_bits_uop_pc_lob = _RANDOM[10'h1DE][12:7];	// lsu.scala:211:16
        stq_3_bits_uop_taken = _RANDOM[10'h1DE][13];	// lsu.scala:211:16
        stq_3_bits_uop_imm_packed = {_RANDOM[10'h1DE][31:14], _RANDOM[10'h1DF][1:0]};	// lsu.scala:211:16
        stq_3_bits_uop_csr_addr = _RANDOM[10'h1DF][13:2];	// lsu.scala:211:16
        stq_3_bits_uop_rob_idx = _RANDOM[10'h1DF][20:14];	// lsu.scala:211:16
        stq_3_bits_uop_ldq_idx = _RANDOM[10'h1DF][25:21];	// lsu.scala:211:16
        stq_3_bits_uop_stq_idx = _RANDOM[10'h1DF][30:26];	// lsu.scala:211:16
        stq_3_bits_uop_rxq_idx = {_RANDOM[10'h1DF][31], _RANDOM[10'h1E0][0]};	// lsu.scala:211:16
        stq_3_bits_uop_pdst = _RANDOM[10'h1E0][7:1];	// lsu.scala:211:16
        stq_3_bits_uop_prs1 = _RANDOM[10'h1E0][14:8];	// lsu.scala:211:16
        stq_3_bits_uop_prs2 = _RANDOM[10'h1E0][21:15];	// lsu.scala:211:16
        stq_3_bits_uop_prs3 = _RANDOM[10'h1E0][28:22];	// lsu.scala:211:16
        stq_3_bits_uop_ppred = {_RANDOM[10'h1E0][31:29], _RANDOM[10'h1E1][1:0]};	// lsu.scala:211:16
        stq_3_bits_uop_prs1_busy = _RANDOM[10'h1E1][2];	// lsu.scala:211:16
        stq_3_bits_uop_prs2_busy = _RANDOM[10'h1E1][3];	// lsu.scala:211:16
        stq_3_bits_uop_prs3_busy = _RANDOM[10'h1E1][4];	// lsu.scala:211:16
        stq_3_bits_uop_ppred_busy = _RANDOM[10'h1E1][5];	// lsu.scala:211:16
        stq_3_bits_uop_stale_pdst = _RANDOM[10'h1E1][12:6];	// lsu.scala:211:16
        stq_3_bits_uop_exception = _RANDOM[10'h1E1][13];	// lsu.scala:211:16
        stq_3_bits_uop_exc_cause =
          {_RANDOM[10'h1E1][31:14], _RANDOM[10'h1E2], _RANDOM[10'h1E3][13:0]};	// lsu.scala:211:16
        stq_3_bits_uop_bypassable = _RANDOM[10'h1E3][14];	// lsu.scala:211:16
        stq_3_bits_uop_mem_cmd = _RANDOM[10'h1E3][19:15];	// lsu.scala:211:16
        stq_3_bits_uop_mem_size = _RANDOM[10'h1E3][21:20];	// lsu.scala:211:16
        stq_3_bits_uop_mem_signed = _RANDOM[10'h1E3][22];	// lsu.scala:211:16
        stq_3_bits_uop_is_fence = _RANDOM[10'h1E3][23];	// lsu.scala:211:16
        stq_3_bits_uop_is_fencei = _RANDOM[10'h1E3][24];	// lsu.scala:211:16
        stq_3_bits_uop_is_amo = _RANDOM[10'h1E3][25];	// lsu.scala:211:16
        stq_3_bits_uop_uses_ldq = _RANDOM[10'h1E3][26];	// lsu.scala:211:16
        stq_3_bits_uop_uses_stq = _RANDOM[10'h1E3][27];	// lsu.scala:211:16
        stq_3_bits_uop_is_sys_pc2epc = _RANDOM[10'h1E3][28];	// lsu.scala:211:16
        stq_3_bits_uop_is_unique = _RANDOM[10'h1E3][29];	// lsu.scala:211:16
        stq_3_bits_uop_flush_on_commit = _RANDOM[10'h1E3][30];	// lsu.scala:211:16
        stq_3_bits_uop_ldst_is_rs1 = _RANDOM[10'h1E3][31];	// lsu.scala:211:16
        stq_3_bits_uop_ldst = _RANDOM[10'h1E4][5:0];	// lsu.scala:211:16
        stq_3_bits_uop_lrs1 = _RANDOM[10'h1E4][11:6];	// lsu.scala:211:16
        stq_3_bits_uop_lrs2 = _RANDOM[10'h1E4][17:12];	// lsu.scala:211:16
        stq_3_bits_uop_lrs3 = _RANDOM[10'h1E4][23:18];	// lsu.scala:211:16
        stq_3_bits_uop_ldst_val = _RANDOM[10'h1E4][24];	// lsu.scala:211:16
        stq_3_bits_uop_dst_rtype = _RANDOM[10'h1E4][26:25];	// lsu.scala:211:16
        stq_3_bits_uop_lrs1_rtype = _RANDOM[10'h1E4][28:27];	// lsu.scala:211:16
        stq_3_bits_uop_lrs2_rtype = _RANDOM[10'h1E4][30:29];	// lsu.scala:211:16
        stq_3_bits_uop_frs3_en = _RANDOM[10'h1E4][31];	// lsu.scala:211:16
        stq_3_bits_uop_fp_val = _RANDOM[10'h1E5][0];	// lsu.scala:211:16
        stq_3_bits_uop_fp_single = _RANDOM[10'h1E5][1];	// lsu.scala:211:16
        stq_3_bits_uop_xcpt_pf_if = _RANDOM[10'h1E5][2];	// lsu.scala:211:16
        stq_3_bits_uop_xcpt_ae_if = _RANDOM[10'h1E5][3];	// lsu.scala:211:16
        stq_3_bits_uop_xcpt_ma_if = _RANDOM[10'h1E5][4];	// lsu.scala:211:16
        stq_3_bits_uop_bp_debug_if = _RANDOM[10'h1E5][5];	// lsu.scala:211:16
        stq_3_bits_uop_bp_xcpt_if = _RANDOM[10'h1E5][6];	// lsu.scala:211:16
        stq_3_bits_uop_debug_fsrc = _RANDOM[10'h1E5][8:7];	// lsu.scala:211:16
        stq_3_bits_uop_debug_tsrc = _RANDOM[10'h1E5][10:9];	// lsu.scala:211:16
        stq_3_bits_addr_valid = _RANDOM[10'h1E5][11];	// lsu.scala:211:16
        stq_3_bits_addr_bits = {_RANDOM[10'h1E5][31:12], _RANDOM[10'h1E6][19:0]};	// lsu.scala:211:16
        stq_3_bits_addr_is_virtual = _RANDOM[10'h1E6][20];	// lsu.scala:211:16
        stq_3_bits_data_valid = _RANDOM[10'h1E6][21];	// lsu.scala:211:16
        stq_3_bits_data_bits =
          {_RANDOM[10'h1E6][31:22], _RANDOM[10'h1E7], _RANDOM[10'h1E8][21:0]};	// lsu.scala:211:16
        stq_3_bits_committed = _RANDOM[10'h1E8][22];	// lsu.scala:211:16
        stq_3_bits_succeeded = _RANDOM[10'h1E8][23];	// lsu.scala:211:16
        stq_4_valid = _RANDOM[10'h1EA][24];	// lsu.scala:211:16
        stq_4_bits_uop_uopc = _RANDOM[10'h1EA][31:25];	// lsu.scala:211:16
        stq_4_bits_uop_inst = _RANDOM[10'h1EB];	// lsu.scala:211:16
        stq_4_bits_uop_debug_inst = _RANDOM[10'h1EC];	// lsu.scala:211:16
        stq_4_bits_uop_is_rvc = _RANDOM[10'h1ED][0];	// lsu.scala:211:16
        stq_4_bits_uop_debug_pc = {_RANDOM[10'h1ED][31:1], _RANDOM[10'h1EE][8:0]};	// lsu.scala:211:16
        stq_4_bits_uop_iq_type = _RANDOM[10'h1EE][11:9];	// lsu.scala:211:16
        stq_4_bits_uop_fu_code = _RANDOM[10'h1EE][21:12];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_br_type = _RANDOM[10'h1EE][25:22];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op1_sel = _RANDOM[10'h1EE][27:26];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op2_sel = _RANDOM[10'h1EE][30:28];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_imm_sel = {_RANDOM[10'h1EE][31], _RANDOM[10'h1EF][1:0]};	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op_fcn = _RANDOM[10'h1EF][5:2];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1EF][6];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1EF][9:7];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_is_load = _RANDOM[10'h1EF][10];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_is_sta = _RANDOM[10'h1EF][11];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_is_std = _RANDOM[10'h1EF][12];	// lsu.scala:211:16
        stq_4_bits_uop_iw_state = _RANDOM[10'h1EF][14:13];	// lsu.scala:211:16
        stq_4_bits_uop_iw_p1_poisoned = _RANDOM[10'h1EF][15];	// lsu.scala:211:16
        stq_4_bits_uop_iw_p2_poisoned = _RANDOM[10'h1EF][16];	// lsu.scala:211:16
        stq_4_bits_uop_is_br = _RANDOM[10'h1EF][17];	// lsu.scala:211:16
        stq_4_bits_uop_is_jalr = _RANDOM[10'h1EF][18];	// lsu.scala:211:16
        stq_4_bits_uop_is_jal = _RANDOM[10'h1EF][19];	// lsu.scala:211:16
        stq_4_bits_uop_is_sfb = _RANDOM[10'h1EF][20];	// lsu.scala:211:16
        stq_4_bits_uop_br_mask = {_RANDOM[10'h1EF][31:21], _RANDOM[10'h1F0][4:0]};	// lsu.scala:211:16
        stq_4_bits_uop_br_tag = _RANDOM[10'h1F0][8:5];	// lsu.scala:211:16
        stq_4_bits_uop_ftq_idx = _RANDOM[10'h1F0][13:9];	// lsu.scala:211:16
        stq_4_bits_uop_edge_inst = _RANDOM[10'h1F0][14];	// lsu.scala:211:16
        stq_4_bits_uop_pc_lob = _RANDOM[10'h1F0][20:15];	// lsu.scala:211:16
        stq_4_bits_uop_taken = _RANDOM[10'h1F0][21];	// lsu.scala:211:16
        stq_4_bits_uop_imm_packed = {_RANDOM[10'h1F0][31:22], _RANDOM[10'h1F1][9:0]};	// lsu.scala:211:16
        stq_4_bits_uop_csr_addr = _RANDOM[10'h1F1][21:10];	// lsu.scala:211:16
        stq_4_bits_uop_rob_idx = _RANDOM[10'h1F1][28:22];	// lsu.scala:211:16
        stq_4_bits_uop_ldq_idx = {_RANDOM[10'h1F1][31:29], _RANDOM[10'h1F2][1:0]};	// lsu.scala:211:16
        stq_4_bits_uop_stq_idx = _RANDOM[10'h1F2][6:2];	// lsu.scala:211:16
        stq_4_bits_uop_rxq_idx = _RANDOM[10'h1F2][8:7];	// lsu.scala:211:16
        stq_4_bits_uop_pdst = _RANDOM[10'h1F2][15:9];	// lsu.scala:211:16
        stq_4_bits_uop_prs1 = _RANDOM[10'h1F2][22:16];	// lsu.scala:211:16
        stq_4_bits_uop_prs2 = _RANDOM[10'h1F2][29:23];	// lsu.scala:211:16
        stq_4_bits_uop_prs3 = {_RANDOM[10'h1F2][31:30], _RANDOM[10'h1F3][4:0]};	// lsu.scala:211:16
        stq_4_bits_uop_ppred = _RANDOM[10'h1F3][9:5];	// lsu.scala:211:16
        stq_4_bits_uop_prs1_busy = _RANDOM[10'h1F3][10];	// lsu.scala:211:16
        stq_4_bits_uop_prs2_busy = _RANDOM[10'h1F3][11];	// lsu.scala:211:16
        stq_4_bits_uop_prs3_busy = _RANDOM[10'h1F3][12];	// lsu.scala:211:16
        stq_4_bits_uop_ppred_busy = _RANDOM[10'h1F3][13];	// lsu.scala:211:16
        stq_4_bits_uop_stale_pdst = _RANDOM[10'h1F3][20:14];	// lsu.scala:211:16
        stq_4_bits_uop_exception = _RANDOM[10'h1F3][21];	// lsu.scala:211:16
        stq_4_bits_uop_exc_cause =
          {_RANDOM[10'h1F3][31:22], _RANDOM[10'h1F4], _RANDOM[10'h1F5][21:0]};	// lsu.scala:211:16
        stq_4_bits_uop_bypassable = _RANDOM[10'h1F5][22];	// lsu.scala:211:16
        stq_4_bits_uop_mem_cmd = _RANDOM[10'h1F5][27:23];	// lsu.scala:211:16
        stq_4_bits_uop_mem_size = _RANDOM[10'h1F5][29:28];	// lsu.scala:211:16
        stq_4_bits_uop_mem_signed = _RANDOM[10'h1F5][30];	// lsu.scala:211:16
        stq_4_bits_uop_is_fence = _RANDOM[10'h1F5][31];	// lsu.scala:211:16
        stq_4_bits_uop_is_fencei = _RANDOM[10'h1F6][0];	// lsu.scala:211:16
        stq_4_bits_uop_is_amo = _RANDOM[10'h1F6][1];	// lsu.scala:211:16
        stq_4_bits_uop_uses_ldq = _RANDOM[10'h1F6][2];	// lsu.scala:211:16
        stq_4_bits_uop_uses_stq = _RANDOM[10'h1F6][3];	// lsu.scala:211:16
        stq_4_bits_uop_is_sys_pc2epc = _RANDOM[10'h1F6][4];	// lsu.scala:211:16
        stq_4_bits_uop_is_unique = _RANDOM[10'h1F6][5];	// lsu.scala:211:16
        stq_4_bits_uop_flush_on_commit = _RANDOM[10'h1F6][6];	// lsu.scala:211:16
        stq_4_bits_uop_ldst_is_rs1 = _RANDOM[10'h1F6][7];	// lsu.scala:211:16
        stq_4_bits_uop_ldst = _RANDOM[10'h1F6][13:8];	// lsu.scala:211:16
        stq_4_bits_uop_lrs1 = _RANDOM[10'h1F6][19:14];	// lsu.scala:211:16
        stq_4_bits_uop_lrs2 = _RANDOM[10'h1F6][25:20];	// lsu.scala:211:16
        stq_4_bits_uop_lrs3 = _RANDOM[10'h1F6][31:26];	// lsu.scala:211:16
        stq_4_bits_uop_ldst_val = _RANDOM[10'h1F7][0];	// lsu.scala:211:16
        stq_4_bits_uop_dst_rtype = _RANDOM[10'h1F7][2:1];	// lsu.scala:211:16
        stq_4_bits_uop_lrs1_rtype = _RANDOM[10'h1F7][4:3];	// lsu.scala:211:16
        stq_4_bits_uop_lrs2_rtype = _RANDOM[10'h1F7][6:5];	// lsu.scala:211:16
        stq_4_bits_uop_frs3_en = _RANDOM[10'h1F7][7];	// lsu.scala:211:16
        stq_4_bits_uop_fp_val = _RANDOM[10'h1F7][8];	// lsu.scala:211:16
        stq_4_bits_uop_fp_single = _RANDOM[10'h1F7][9];	// lsu.scala:211:16
        stq_4_bits_uop_xcpt_pf_if = _RANDOM[10'h1F7][10];	// lsu.scala:211:16
        stq_4_bits_uop_xcpt_ae_if = _RANDOM[10'h1F7][11];	// lsu.scala:211:16
        stq_4_bits_uop_xcpt_ma_if = _RANDOM[10'h1F7][12];	// lsu.scala:211:16
        stq_4_bits_uop_bp_debug_if = _RANDOM[10'h1F7][13];	// lsu.scala:211:16
        stq_4_bits_uop_bp_xcpt_if = _RANDOM[10'h1F7][14];	// lsu.scala:211:16
        stq_4_bits_uop_debug_fsrc = _RANDOM[10'h1F7][16:15];	// lsu.scala:211:16
        stq_4_bits_uop_debug_tsrc = _RANDOM[10'h1F7][18:17];	// lsu.scala:211:16
        stq_4_bits_addr_valid = _RANDOM[10'h1F7][19];	// lsu.scala:211:16
        stq_4_bits_addr_bits = {_RANDOM[10'h1F7][31:20], _RANDOM[10'h1F8][27:0]};	// lsu.scala:211:16
        stq_4_bits_addr_is_virtual = _RANDOM[10'h1F8][28];	// lsu.scala:211:16
        stq_4_bits_data_valid = _RANDOM[10'h1F8][29];	// lsu.scala:211:16
        stq_4_bits_data_bits =
          {_RANDOM[10'h1F8][31:30], _RANDOM[10'h1F9], _RANDOM[10'h1FA][29:0]};	// lsu.scala:211:16
        stq_4_bits_committed = _RANDOM[10'h1FA][30];	// lsu.scala:211:16
        stq_4_bits_succeeded = _RANDOM[10'h1FA][31];	// lsu.scala:211:16
        stq_5_valid = _RANDOM[10'h1FD][0];	// lsu.scala:211:16
        stq_5_bits_uop_uopc = _RANDOM[10'h1FD][7:1];	// lsu.scala:211:16
        stq_5_bits_uop_inst = {_RANDOM[10'h1FD][31:8], _RANDOM[10'h1FE][7:0]};	// lsu.scala:211:16
        stq_5_bits_uop_debug_inst = {_RANDOM[10'h1FE][31:8], _RANDOM[10'h1FF][7:0]};	// lsu.scala:211:16
        stq_5_bits_uop_is_rvc = _RANDOM[10'h1FF][8];	// lsu.scala:211:16
        stq_5_bits_uop_debug_pc = {_RANDOM[10'h1FF][31:9], _RANDOM[10'h200][16:0]};	// lsu.scala:211:16
        stq_5_bits_uop_iq_type = _RANDOM[10'h200][19:17];	// lsu.scala:211:16
        stq_5_bits_uop_fu_code = _RANDOM[10'h200][29:20];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_br_type = {_RANDOM[10'h200][31:30], _RANDOM[10'h201][1:0]};	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op1_sel = _RANDOM[10'h201][3:2];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op2_sel = _RANDOM[10'h201][6:4];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_imm_sel = _RANDOM[10'h201][9:7];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op_fcn = _RANDOM[10'h201][13:10];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_fcn_dw = _RANDOM[10'h201][14];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_csr_cmd = _RANDOM[10'h201][17:15];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_is_load = _RANDOM[10'h201][18];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_is_sta = _RANDOM[10'h201][19];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_is_std = _RANDOM[10'h201][20];	// lsu.scala:211:16
        stq_5_bits_uop_iw_state = _RANDOM[10'h201][22:21];	// lsu.scala:211:16
        stq_5_bits_uop_iw_p1_poisoned = _RANDOM[10'h201][23];	// lsu.scala:211:16
        stq_5_bits_uop_iw_p2_poisoned = _RANDOM[10'h201][24];	// lsu.scala:211:16
        stq_5_bits_uop_is_br = _RANDOM[10'h201][25];	// lsu.scala:211:16
        stq_5_bits_uop_is_jalr = _RANDOM[10'h201][26];	// lsu.scala:211:16
        stq_5_bits_uop_is_jal = _RANDOM[10'h201][27];	// lsu.scala:211:16
        stq_5_bits_uop_is_sfb = _RANDOM[10'h201][28];	// lsu.scala:211:16
        stq_5_bits_uop_br_mask = {_RANDOM[10'h201][31:29], _RANDOM[10'h202][12:0]};	// lsu.scala:211:16
        stq_5_bits_uop_br_tag = _RANDOM[10'h202][16:13];	// lsu.scala:211:16
        stq_5_bits_uop_ftq_idx = _RANDOM[10'h202][21:17];	// lsu.scala:211:16
        stq_5_bits_uop_edge_inst = _RANDOM[10'h202][22];	// lsu.scala:211:16
        stq_5_bits_uop_pc_lob = _RANDOM[10'h202][28:23];	// lsu.scala:211:16
        stq_5_bits_uop_taken = _RANDOM[10'h202][29];	// lsu.scala:211:16
        stq_5_bits_uop_imm_packed = {_RANDOM[10'h202][31:30], _RANDOM[10'h203][17:0]};	// lsu.scala:211:16
        stq_5_bits_uop_csr_addr = _RANDOM[10'h203][29:18];	// lsu.scala:211:16
        stq_5_bits_uop_rob_idx = {_RANDOM[10'h203][31:30], _RANDOM[10'h204][4:0]};	// lsu.scala:211:16
        stq_5_bits_uop_ldq_idx = _RANDOM[10'h204][9:5];	// lsu.scala:211:16
        stq_5_bits_uop_stq_idx = _RANDOM[10'h204][14:10];	// lsu.scala:211:16
        stq_5_bits_uop_rxq_idx = _RANDOM[10'h204][16:15];	// lsu.scala:211:16
        stq_5_bits_uop_pdst = _RANDOM[10'h204][23:17];	// lsu.scala:211:16
        stq_5_bits_uop_prs1 = _RANDOM[10'h204][30:24];	// lsu.scala:211:16
        stq_5_bits_uop_prs2 = {_RANDOM[10'h204][31], _RANDOM[10'h205][5:0]};	// lsu.scala:211:16
        stq_5_bits_uop_prs3 = _RANDOM[10'h205][12:6];	// lsu.scala:211:16
        stq_5_bits_uop_ppred = _RANDOM[10'h205][17:13];	// lsu.scala:211:16
        stq_5_bits_uop_prs1_busy = _RANDOM[10'h205][18];	// lsu.scala:211:16
        stq_5_bits_uop_prs2_busy = _RANDOM[10'h205][19];	// lsu.scala:211:16
        stq_5_bits_uop_prs3_busy = _RANDOM[10'h205][20];	// lsu.scala:211:16
        stq_5_bits_uop_ppred_busy = _RANDOM[10'h205][21];	// lsu.scala:211:16
        stq_5_bits_uop_stale_pdst = _RANDOM[10'h205][28:22];	// lsu.scala:211:16
        stq_5_bits_uop_exception = _RANDOM[10'h205][29];	// lsu.scala:211:16
        stq_5_bits_uop_exc_cause =
          {_RANDOM[10'h205][31:30], _RANDOM[10'h206], _RANDOM[10'h207][29:0]};	// lsu.scala:211:16
        stq_5_bits_uop_bypassable = _RANDOM[10'h207][30];	// lsu.scala:211:16
        stq_5_bits_uop_mem_cmd = {_RANDOM[10'h207][31], _RANDOM[10'h208][3:0]};	// lsu.scala:211:16
        stq_5_bits_uop_mem_size = _RANDOM[10'h208][5:4];	// lsu.scala:211:16
        stq_5_bits_uop_mem_signed = _RANDOM[10'h208][6];	// lsu.scala:211:16
        stq_5_bits_uop_is_fence = _RANDOM[10'h208][7];	// lsu.scala:211:16
        stq_5_bits_uop_is_fencei = _RANDOM[10'h208][8];	// lsu.scala:211:16
        stq_5_bits_uop_is_amo = _RANDOM[10'h208][9];	// lsu.scala:211:16
        stq_5_bits_uop_uses_ldq = _RANDOM[10'h208][10];	// lsu.scala:211:16
        stq_5_bits_uop_uses_stq = _RANDOM[10'h208][11];	// lsu.scala:211:16
        stq_5_bits_uop_is_sys_pc2epc = _RANDOM[10'h208][12];	// lsu.scala:211:16
        stq_5_bits_uop_is_unique = _RANDOM[10'h208][13];	// lsu.scala:211:16
        stq_5_bits_uop_flush_on_commit = _RANDOM[10'h208][14];	// lsu.scala:211:16
        stq_5_bits_uop_ldst_is_rs1 = _RANDOM[10'h208][15];	// lsu.scala:211:16
        stq_5_bits_uop_ldst = _RANDOM[10'h208][21:16];	// lsu.scala:211:16
        stq_5_bits_uop_lrs1 = _RANDOM[10'h208][27:22];	// lsu.scala:211:16
        stq_5_bits_uop_lrs2 = {_RANDOM[10'h208][31:28], _RANDOM[10'h209][1:0]};	// lsu.scala:211:16
        stq_5_bits_uop_lrs3 = _RANDOM[10'h209][7:2];	// lsu.scala:211:16
        stq_5_bits_uop_ldst_val = _RANDOM[10'h209][8];	// lsu.scala:211:16
        stq_5_bits_uop_dst_rtype = _RANDOM[10'h209][10:9];	// lsu.scala:211:16
        stq_5_bits_uop_lrs1_rtype = _RANDOM[10'h209][12:11];	// lsu.scala:211:16
        stq_5_bits_uop_lrs2_rtype = _RANDOM[10'h209][14:13];	// lsu.scala:211:16
        stq_5_bits_uop_frs3_en = _RANDOM[10'h209][15];	// lsu.scala:211:16
        stq_5_bits_uop_fp_val = _RANDOM[10'h209][16];	// lsu.scala:211:16
        stq_5_bits_uop_fp_single = _RANDOM[10'h209][17];	// lsu.scala:211:16
        stq_5_bits_uop_xcpt_pf_if = _RANDOM[10'h209][18];	// lsu.scala:211:16
        stq_5_bits_uop_xcpt_ae_if = _RANDOM[10'h209][19];	// lsu.scala:211:16
        stq_5_bits_uop_xcpt_ma_if = _RANDOM[10'h209][20];	// lsu.scala:211:16
        stq_5_bits_uop_bp_debug_if = _RANDOM[10'h209][21];	// lsu.scala:211:16
        stq_5_bits_uop_bp_xcpt_if = _RANDOM[10'h209][22];	// lsu.scala:211:16
        stq_5_bits_uop_debug_fsrc = _RANDOM[10'h209][24:23];	// lsu.scala:211:16
        stq_5_bits_uop_debug_tsrc = _RANDOM[10'h209][26:25];	// lsu.scala:211:16
        stq_5_bits_addr_valid = _RANDOM[10'h209][27];	// lsu.scala:211:16
        stq_5_bits_addr_bits =
          {_RANDOM[10'h209][31:28], _RANDOM[10'h20A], _RANDOM[10'h20B][3:0]};	// lsu.scala:211:16
        stq_5_bits_addr_is_virtual = _RANDOM[10'h20B][4];	// lsu.scala:211:16
        stq_5_bits_data_valid = _RANDOM[10'h20B][5];	// lsu.scala:211:16
        stq_5_bits_data_bits =
          {_RANDOM[10'h20B][31:6], _RANDOM[10'h20C], _RANDOM[10'h20D][5:0]};	// lsu.scala:211:16
        stq_5_bits_committed = _RANDOM[10'h20D][6];	// lsu.scala:211:16
        stq_5_bits_succeeded = _RANDOM[10'h20D][7];	// lsu.scala:211:16
        stq_6_valid = _RANDOM[10'h20F][8];	// lsu.scala:211:16
        stq_6_bits_uop_uopc = _RANDOM[10'h20F][15:9];	// lsu.scala:211:16
        stq_6_bits_uop_inst = {_RANDOM[10'h20F][31:16], _RANDOM[10'h210][15:0]};	// lsu.scala:211:16
        stq_6_bits_uop_debug_inst = {_RANDOM[10'h210][31:16], _RANDOM[10'h211][15:0]};	// lsu.scala:211:16
        stq_6_bits_uop_is_rvc = _RANDOM[10'h211][16];	// lsu.scala:211:16
        stq_6_bits_uop_debug_pc = {_RANDOM[10'h211][31:17], _RANDOM[10'h212][24:0]};	// lsu.scala:211:16
        stq_6_bits_uop_iq_type = _RANDOM[10'h212][27:25];	// lsu.scala:211:16
        stq_6_bits_uop_fu_code = {_RANDOM[10'h212][31:28], _RANDOM[10'h213][5:0]};	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_br_type = _RANDOM[10'h213][9:6];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op1_sel = _RANDOM[10'h213][11:10];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op2_sel = _RANDOM[10'h213][14:12];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_imm_sel = _RANDOM[10'h213][17:15];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op_fcn = _RANDOM[10'h213][21:18];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_fcn_dw = _RANDOM[10'h213][22];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_csr_cmd = _RANDOM[10'h213][25:23];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_is_load = _RANDOM[10'h213][26];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_is_sta = _RANDOM[10'h213][27];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_is_std = _RANDOM[10'h213][28];	// lsu.scala:211:16
        stq_6_bits_uop_iw_state = _RANDOM[10'h213][30:29];	// lsu.scala:211:16
        stq_6_bits_uop_iw_p1_poisoned = _RANDOM[10'h213][31];	// lsu.scala:211:16
        stq_6_bits_uop_iw_p2_poisoned = _RANDOM[10'h214][0];	// lsu.scala:211:16
        stq_6_bits_uop_is_br = _RANDOM[10'h214][1];	// lsu.scala:211:16
        stq_6_bits_uop_is_jalr = _RANDOM[10'h214][2];	// lsu.scala:211:16
        stq_6_bits_uop_is_jal = _RANDOM[10'h214][3];	// lsu.scala:211:16
        stq_6_bits_uop_is_sfb = _RANDOM[10'h214][4];	// lsu.scala:211:16
        stq_6_bits_uop_br_mask = _RANDOM[10'h214][20:5];	// lsu.scala:211:16
        stq_6_bits_uop_br_tag = _RANDOM[10'h214][24:21];	// lsu.scala:211:16
        stq_6_bits_uop_ftq_idx = _RANDOM[10'h214][29:25];	// lsu.scala:211:16
        stq_6_bits_uop_edge_inst = _RANDOM[10'h214][30];	// lsu.scala:211:16
        stq_6_bits_uop_pc_lob = {_RANDOM[10'h214][31], _RANDOM[10'h215][4:0]};	// lsu.scala:211:16
        stq_6_bits_uop_taken = _RANDOM[10'h215][5];	// lsu.scala:211:16
        stq_6_bits_uop_imm_packed = _RANDOM[10'h215][25:6];	// lsu.scala:211:16
        stq_6_bits_uop_csr_addr = {_RANDOM[10'h215][31:26], _RANDOM[10'h216][5:0]};	// lsu.scala:211:16
        stq_6_bits_uop_rob_idx = _RANDOM[10'h216][12:6];	// lsu.scala:211:16
        stq_6_bits_uop_ldq_idx = _RANDOM[10'h216][17:13];	// lsu.scala:211:16
        stq_6_bits_uop_stq_idx = _RANDOM[10'h216][22:18];	// lsu.scala:211:16
        stq_6_bits_uop_rxq_idx = _RANDOM[10'h216][24:23];	// lsu.scala:211:16
        stq_6_bits_uop_pdst = _RANDOM[10'h216][31:25];	// lsu.scala:211:16
        stq_6_bits_uop_prs1 = _RANDOM[10'h217][6:0];	// lsu.scala:211:16
        stq_6_bits_uop_prs2 = _RANDOM[10'h217][13:7];	// lsu.scala:211:16
        stq_6_bits_uop_prs3 = _RANDOM[10'h217][20:14];	// lsu.scala:211:16
        stq_6_bits_uop_ppred = _RANDOM[10'h217][25:21];	// lsu.scala:211:16
        stq_6_bits_uop_prs1_busy = _RANDOM[10'h217][26];	// lsu.scala:211:16
        stq_6_bits_uop_prs2_busy = _RANDOM[10'h217][27];	// lsu.scala:211:16
        stq_6_bits_uop_prs3_busy = _RANDOM[10'h217][28];	// lsu.scala:211:16
        stq_6_bits_uop_ppred_busy = _RANDOM[10'h217][29];	// lsu.scala:211:16
        stq_6_bits_uop_stale_pdst = {_RANDOM[10'h217][31:30], _RANDOM[10'h218][4:0]};	// lsu.scala:211:16
        stq_6_bits_uop_exception = _RANDOM[10'h218][5];	// lsu.scala:211:16
        stq_6_bits_uop_exc_cause =
          {_RANDOM[10'h218][31:6], _RANDOM[10'h219], _RANDOM[10'h21A][5:0]};	// lsu.scala:211:16
        stq_6_bits_uop_bypassable = _RANDOM[10'h21A][6];	// lsu.scala:211:16
        stq_6_bits_uop_mem_cmd = _RANDOM[10'h21A][11:7];	// lsu.scala:211:16
        stq_6_bits_uop_mem_size = _RANDOM[10'h21A][13:12];	// lsu.scala:211:16
        stq_6_bits_uop_mem_signed = _RANDOM[10'h21A][14];	// lsu.scala:211:16
        stq_6_bits_uop_is_fence = _RANDOM[10'h21A][15];	// lsu.scala:211:16
        stq_6_bits_uop_is_fencei = _RANDOM[10'h21A][16];	// lsu.scala:211:16
        stq_6_bits_uop_is_amo = _RANDOM[10'h21A][17];	// lsu.scala:211:16
        stq_6_bits_uop_uses_ldq = _RANDOM[10'h21A][18];	// lsu.scala:211:16
        stq_6_bits_uop_uses_stq = _RANDOM[10'h21A][19];	// lsu.scala:211:16
        stq_6_bits_uop_is_sys_pc2epc = _RANDOM[10'h21A][20];	// lsu.scala:211:16
        stq_6_bits_uop_is_unique = _RANDOM[10'h21A][21];	// lsu.scala:211:16
        stq_6_bits_uop_flush_on_commit = _RANDOM[10'h21A][22];	// lsu.scala:211:16
        stq_6_bits_uop_ldst_is_rs1 = _RANDOM[10'h21A][23];	// lsu.scala:211:16
        stq_6_bits_uop_ldst = _RANDOM[10'h21A][29:24];	// lsu.scala:211:16
        stq_6_bits_uop_lrs1 = {_RANDOM[10'h21A][31:30], _RANDOM[10'h21B][3:0]};	// lsu.scala:211:16
        stq_6_bits_uop_lrs2 = _RANDOM[10'h21B][9:4];	// lsu.scala:211:16
        stq_6_bits_uop_lrs3 = _RANDOM[10'h21B][15:10];	// lsu.scala:211:16
        stq_6_bits_uop_ldst_val = _RANDOM[10'h21B][16];	// lsu.scala:211:16
        stq_6_bits_uop_dst_rtype = _RANDOM[10'h21B][18:17];	// lsu.scala:211:16
        stq_6_bits_uop_lrs1_rtype = _RANDOM[10'h21B][20:19];	// lsu.scala:211:16
        stq_6_bits_uop_lrs2_rtype = _RANDOM[10'h21B][22:21];	// lsu.scala:211:16
        stq_6_bits_uop_frs3_en = _RANDOM[10'h21B][23];	// lsu.scala:211:16
        stq_6_bits_uop_fp_val = _RANDOM[10'h21B][24];	// lsu.scala:211:16
        stq_6_bits_uop_fp_single = _RANDOM[10'h21B][25];	// lsu.scala:211:16
        stq_6_bits_uop_xcpt_pf_if = _RANDOM[10'h21B][26];	// lsu.scala:211:16
        stq_6_bits_uop_xcpt_ae_if = _RANDOM[10'h21B][27];	// lsu.scala:211:16
        stq_6_bits_uop_xcpt_ma_if = _RANDOM[10'h21B][28];	// lsu.scala:211:16
        stq_6_bits_uop_bp_debug_if = _RANDOM[10'h21B][29];	// lsu.scala:211:16
        stq_6_bits_uop_bp_xcpt_if = _RANDOM[10'h21B][30];	// lsu.scala:211:16
        stq_6_bits_uop_debug_fsrc = {_RANDOM[10'h21B][31], _RANDOM[10'h21C][0]};	// lsu.scala:211:16
        stq_6_bits_uop_debug_tsrc = _RANDOM[10'h21C][2:1];	// lsu.scala:211:16
        stq_6_bits_addr_valid = _RANDOM[10'h21C][3];	// lsu.scala:211:16
        stq_6_bits_addr_bits = {_RANDOM[10'h21C][31:4], _RANDOM[10'h21D][11:0]};	// lsu.scala:211:16
        stq_6_bits_addr_is_virtual = _RANDOM[10'h21D][12];	// lsu.scala:211:16
        stq_6_bits_data_valid = _RANDOM[10'h21D][13];	// lsu.scala:211:16
        stq_6_bits_data_bits =
          {_RANDOM[10'h21D][31:14], _RANDOM[10'h21E], _RANDOM[10'h21F][13:0]};	// lsu.scala:211:16
        stq_6_bits_committed = _RANDOM[10'h21F][14];	// lsu.scala:211:16
        stq_6_bits_succeeded = _RANDOM[10'h21F][15];	// lsu.scala:211:16
        stq_7_valid = _RANDOM[10'h221][16];	// lsu.scala:211:16
        stq_7_bits_uop_uopc = _RANDOM[10'h221][23:17];	// lsu.scala:211:16
        stq_7_bits_uop_inst = {_RANDOM[10'h221][31:24], _RANDOM[10'h222][23:0]};	// lsu.scala:211:16
        stq_7_bits_uop_debug_inst = {_RANDOM[10'h222][31:24], _RANDOM[10'h223][23:0]};	// lsu.scala:211:16
        stq_7_bits_uop_is_rvc = _RANDOM[10'h223][24];	// lsu.scala:211:16
        stq_7_bits_uop_debug_pc =
          {_RANDOM[10'h223][31:25], _RANDOM[10'h224], _RANDOM[10'h225][0]};	// lsu.scala:211:16
        stq_7_bits_uop_iq_type = _RANDOM[10'h225][3:1];	// lsu.scala:211:16
        stq_7_bits_uop_fu_code = _RANDOM[10'h225][13:4];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_br_type = _RANDOM[10'h225][17:14];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op1_sel = _RANDOM[10'h225][19:18];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op2_sel = _RANDOM[10'h225][22:20];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_imm_sel = _RANDOM[10'h225][25:23];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op_fcn = _RANDOM[10'h225][29:26];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_fcn_dw = _RANDOM[10'h225][30];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h225][31], _RANDOM[10'h226][1:0]};	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_is_load = _RANDOM[10'h226][2];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_is_sta = _RANDOM[10'h226][3];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_is_std = _RANDOM[10'h226][4];	// lsu.scala:211:16
        stq_7_bits_uop_iw_state = _RANDOM[10'h226][6:5];	// lsu.scala:211:16
        stq_7_bits_uop_iw_p1_poisoned = _RANDOM[10'h226][7];	// lsu.scala:211:16
        stq_7_bits_uop_iw_p2_poisoned = _RANDOM[10'h226][8];	// lsu.scala:211:16
        stq_7_bits_uop_is_br = _RANDOM[10'h226][9];	// lsu.scala:211:16
        stq_7_bits_uop_is_jalr = _RANDOM[10'h226][10];	// lsu.scala:211:16
        stq_7_bits_uop_is_jal = _RANDOM[10'h226][11];	// lsu.scala:211:16
        stq_7_bits_uop_is_sfb = _RANDOM[10'h226][12];	// lsu.scala:211:16
        stq_7_bits_uop_br_mask = _RANDOM[10'h226][28:13];	// lsu.scala:211:16
        stq_7_bits_uop_br_tag = {_RANDOM[10'h226][31:29], _RANDOM[10'h227][0]};	// lsu.scala:211:16
        stq_7_bits_uop_ftq_idx = _RANDOM[10'h227][5:1];	// lsu.scala:211:16
        stq_7_bits_uop_edge_inst = _RANDOM[10'h227][6];	// lsu.scala:211:16
        stq_7_bits_uop_pc_lob = _RANDOM[10'h227][12:7];	// lsu.scala:211:16
        stq_7_bits_uop_taken = _RANDOM[10'h227][13];	// lsu.scala:211:16
        stq_7_bits_uop_imm_packed = {_RANDOM[10'h227][31:14], _RANDOM[10'h228][1:0]};	// lsu.scala:211:16
        stq_7_bits_uop_csr_addr = _RANDOM[10'h228][13:2];	// lsu.scala:211:16
        stq_7_bits_uop_rob_idx = _RANDOM[10'h228][20:14];	// lsu.scala:211:16
        stq_7_bits_uop_ldq_idx = _RANDOM[10'h228][25:21];	// lsu.scala:211:16
        stq_7_bits_uop_stq_idx = _RANDOM[10'h228][30:26];	// lsu.scala:211:16
        stq_7_bits_uop_rxq_idx = {_RANDOM[10'h228][31], _RANDOM[10'h229][0]};	// lsu.scala:211:16
        stq_7_bits_uop_pdst = _RANDOM[10'h229][7:1];	// lsu.scala:211:16
        stq_7_bits_uop_prs1 = _RANDOM[10'h229][14:8];	// lsu.scala:211:16
        stq_7_bits_uop_prs2 = _RANDOM[10'h229][21:15];	// lsu.scala:211:16
        stq_7_bits_uop_prs3 = _RANDOM[10'h229][28:22];	// lsu.scala:211:16
        stq_7_bits_uop_ppred = {_RANDOM[10'h229][31:29], _RANDOM[10'h22A][1:0]};	// lsu.scala:211:16
        stq_7_bits_uop_prs1_busy = _RANDOM[10'h22A][2];	// lsu.scala:211:16
        stq_7_bits_uop_prs2_busy = _RANDOM[10'h22A][3];	// lsu.scala:211:16
        stq_7_bits_uop_prs3_busy = _RANDOM[10'h22A][4];	// lsu.scala:211:16
        stq_7_bits_uop_ppred_busy = _RANDOM[10'h22A][5];	// lsu.scala:211:16
        stq_7_bits_uop_stale_pdst = _RANDOM[10'h22A][12:6];	// lsu.scala:211:16
        stq_7_bits_uop_exception = _RANDOM[10'h22A][13];	// lsu.scala:211:16
        stq_7_bits_uop_exc_cause =
          {_RANDOM[10'h22A][31:14], _RANDOM[10'h22B], _RANDOM[10'h22C][13:0]};	// lsu.scala:211:16
        stq_7_bits_uop_bypassable = _RANDOM[10'h22C][14];	// lsu.scala:211:16
        stq_7_bits_uop_mem_cmd = _RANDOM[10'h22C][19:15];	// lsu.scala:211:16
        stq_7_bits_uop_mem_size = _RANDOM[10'h22C][21:20];	// lsu.scala:211:16
        stq_7_bits_uop_mem_signed = _RANDOM[10'h22C][22];	// lsu.scala:211:16
        stq_7_bits_uop_is_fence = _RANDOM[10'h22C][23];	// lsu.scala:211:16
        stq_7_bits_uop_is_fencei = _RANDOM[10'h22C][24];	// lsu.scala:211:16
        stq_7_bits_uop_is_amo = _RANDOM[10'h22C][25];	// lsu.scala:211:16
        stq_7_bits_uop_uses_ldq = _RANDOM[10'h22C][26];	// lsu.scala:211:16
        stq_7_bits_uop_uses_stq = _RANDOM[10'h22C][27];	// lsu.scala:211:16
        stq_7_bits_uop_is_sys_pc2epc = _RANDOM[10'h22C][28];	// lsu.scala:211:16
        stq_7_bits_uop_is_unique = _RANDOM[10'h22C][29];	// lsu.scala:211:16
        stq_7_bits_uop_flush_on_commit = _RANDOM[10'h22C][30];	// lsu.scala:211:16
        stq_7_bits_uop_ldst_is_rs1 = _RANDOM[10'h22C][31];	// lsu.scala:211:16
        stq_7_bits_uop_ldst = _RANDOM[10'h22D][5:0];	// lsu.scala:211:16
        stq_7_bits_uop_lrs1 = _RANDOM[10'h22D][11:6];	// lsu.scala:211:16
        stq_7_bits_uop_lrs2 = _RANDOM[10'h22D][17:12];	// lsu.scala:211:16
        stq_7_bits_uop_lrs3 = _RANDOM[10'h22D][23:18];	// lsu.scala:211:16
        stq_7_bits_uop_ldst_val = _RANDOM[10'h22D][24];	// lsu.scala:211:16
        stq_7_bits_uop_dst_rtype = _RANDOM[10'h22D][26:25];	// lsu.scala:211:16
        stq_7_bits_uop_lrs1_rtype = _RANDOM[10'h22D][28:27];	// lsu.scala:211:16
        stq_7_bits_uop_lrs2_rtype = _RANDOM[10'h22D][30:29];	// lsu.scala:211:16
        stq_7_bits_uop_frs3_en = _RANDOM[10'h22D][31];	// lsu.scala:211:16
        stq_7_bits_uop_fp_val = _RANDOM[10'h22E][0];	// lsu.scala:211:16
        stq_7_bits_uop_fp_single = _RANDOM[10'h22E][1];	// lsu.scala:211:16
        stq_7_bits_uop_xcpt_pf_if = _RANDOM[10'h22E][2];	// lsu.scala:211:16
        stq_7_bits_uop_xcpt_ae_if = _RANDOM[10'h22E][3];	// lsu.scala:211:16
        stq_7_bits_uop_xcpt_ma_if = _RANDOM[10'h22E][4];	// lsu.scala:211:16
        stq_7_bits_uop_bp_debug_if = _RANDOM[10'h22E][5];	// lsu.scala:211:16
        stq_7_bits_uop_bp_xcpt_if = _RANDOM[10'h22E][6];	// lsu.scala:211:16
        stq_7_bits_uop_debug_fsrc = _RANDOM[10'h22E][8:7];	// lsu.scala:211:16
        stq_7_bits_uop_debug_tsrc = _RANDOM[10'h22E][10:9];	// lsu.scala:211:16
        stq_7_bits_addr_valid = _RANDOM[10'h22E][11];	// lsu.scala:211:16
        stq_7_bits_addr_bits = {_RANDOM[10'h22E][31:12], _RANDOM[10'h22F][19:0]};	// lsu.scala:211:16
        stq_7_bits_addr_is_virtual = _RANDOM[10'h22F][20];	// lsu.scala:211:16
        stq_7_bits_data_valid = _RANDOM[10'h22F][21];	// lsu.scala:211:16
        stq_7_bits_data_bits =
          {_RANDOM[10'h22F][31:22], _RANDOM[10'h230], _RANDOM[10'h231][21:0]};	// lsu.scala:211:16
        stq_7_bits_committed = _RANDOM[10'h231][22];	// lsu.scala:211:16
        stq_7_bits_succeeded = _RANDOM[10'h231][23];	// lsu.scala:211:16
        stq_8_valid = _RANDOM[10'h233][24];	// lsu.scala:211:16
        stq_8_bits_uop_uopc = _RANDOM[10'h233][31:25];	// lsu.scala:211:16
        stq_8_bits_uop_inst = _RANDOM[10'h234];	// lsu.scala:211:16
        stq_8_bits_uop_debug_inst = _RANDOM[10'h235];	// lsu.scala:211:16
        stq_8_bits_uop_is_rvc = _RANDOM[10'h236][0];	// lsu.scala:211:16
        stq_8_bits_uop_debug_pc = {_RANDOM[10'h236][31:1], _RANDOM[10'h237][8:0]};	// lsu.scala:211:16
        stq_8_bits_uop_iq_type = _RANDOM[10'h237][11:9];	// lsu.scala:211:16
        stq_8_bits_uop_fu_code = _RANDOM[10'h237][21:12];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_br_type = _RANDOM[10'h237][25:22];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op1_sel = _RANDOM[10'h237][27:26];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op2_sel = _RANDOM[10'h237][30:28];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_imm_sel = {_RANDOM[10'h237][31], _RANDOM[10'h238][1:0]};	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op_fcn = _RANDOM[10'h238][5:2];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_fcn_dw = _RANDOM[10'h238][6];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_csr_cmd = _RANDOM[10'h238][9:7];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_is_load = _RANDOM[10'h238][10];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_is_sta = _RANDOM[10'h238][11];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_is_std = _RANDOM[10'h238][12];	// lsu.scala:211:16
        stq_8_bits_uop_iw_state = _RANDOM[10'h238][14:13];	// lsu.scala:211:16
        stq_8_bits_uop_iw_p1_poisoned = _RANDOM[10'h238][15];	// lsu.scala:211:16
        stq_8_bits_uop_iw_p2_poisoned = _RANDOM[10'h238][16];	// lsu.scala:211:16
        stq_8_bits_uop_is_br = _RANDOM[10'h238][17];	// lsu.scala:211:16
        stq_8_bits_uop_is_jalr = _RANDOM[10'h238][18];	// lsu.scala:211:16
        stq_8_bits_uop_is_jal = _RANDOM[10'h238][19];	// lsu.scala:211:16
        stq_8_bits_uop_is_sfb = _RANDOM[10'h238][20];	// lsu.scala:211:16
        stq_8_bits_uop_br_mask = {_RANDOM[10'h238][31:21], _RANDOM[10'h239][4:0]};	// lsu.scala:211:16
        stq_8_bits_uop_br_tag = _RANDOM[10'h239][8:5];	// lsu.scala:211:16
        stq_8_bits_uop_ftq_idx = _RANDOM[10'h239][13:9];	// lsu.scala:211:16
        stq_8_bits_uop_edge_inst = _RANDOM[10'h239][14];	// lsu.scala:211:16
        stq_8_bits_uop_pc_lob = _RANDOM[10'h239][20:15];	// lsu.scala:211:16
        stq_8_bits_uop_taken = _RANDOM[10'h239][21];	// lsu.scala:211:16
        stq_8_bits_uop_imm_packed = {_RANDOM[10'h239][31:22], _RANDOM[10'h23A][9:0]};	// lsu.scala:211:16
        stq_8_bits_uop_csr_addr = _RANDOM[10'h23A][21:10];	// lsu.scala:211:16
        stq_8_bits_uop_rob_idx = _RANDOM[10'h23A][28:22];	// lsu.scala:211:16
        stq_8_bits_uop_ldq_idx = {_RANDOM[10'h23A][31:29], _RANDOM[10'h23B][1:0]};	// lsu.scala:211:16
        stq_8_bits_uop_stq_idx = _RANDOM[10'h23B][6:2];	// lsu.scala:211:16
        stq_8_bits_uop_rxq_idx = _RANDOM[10'h23B][8:7];	// lsu.scala:211:16
        stq_8_bits_uop_pdst = _RANDOM[10'h23B][15:9];	// lsu.scala:211:16
        stq_8_bits_uop_prs1 = _RANDOM[10'h23B][22:16];	// lsu.scala:211:16
        stq_8_bits_uop_prs2 = _RANDOM[10'h23B][29:23];	// lsu.scala:211:16
        stq_8_bits_uop_prs3 = {_RANDOM[10'h23B][31:30], _RANDOM[10'h23C][4:0]};	// lsu.scala:211:16
        stq_8_bits_uop_ppred = _RANDOM[10'h23C][9:5];	// lsu.scala:211:16
        stq_8_bits_uop_prs1_busy = _RANDOM[10'h23C][10];	// lsu.scala:211:16
        stq_8_bits_uop_prs2_busy = _RANDOM[10'h23C][11];	// lsu.scala:211:16
        stq_8_bits_uop_prs3_busy = _RANDOM[10'h23C][12];	// lsu.scala:211:16
        stq_8_bits_uop_ppred_busy = _RANDOM[10'h23C][13];	// lsu.scala:211:16
        stq_8_bits_uop_stale_pdst = _RANDOM[10'h23C][20:14];	// lsu.scala:211:16
        stq_8_bits_uop_exception = _RANDOM[10'h23C][21];	// lsu.scala:211:16
        stq_8_bits_uop_exc_cause =
          {_RANDOM[10'h23C][31:22], _RANDOM[10'h23D], _RANDOM[10'h23E][21:0]};	// lsu.scala:211:16
        stq_8_bits_uop_bypassable = _RANDOM[10'h23E][22];	// lsu.scala:211:16
        stq_8_bits_uop_mem_cmd = _RANDOM[10'h23E][27:23];	// lsu.scala:211:16
        stq_8_bits_uop_mem_size = _RANDOM[10'h23E][29:28];	// lsu.scala:211:16
        stq_8_bits_uop_mem_signed = _RANDOM[10'h23E][30];	// lsu.scala:211:16
        stq_8_bits_uop_is_fence = _RANDOM[10'h23E][31];	// lsu.scala:211:16
        stq_8_bits_uop_is_fencei = _RANDOM[10'h23F][0];	// lsu.scala:211:16
        stq_8_bits_uop_is_amo = _RANDOM[10'h23F][1];	// lsu.scala:211:16
        stq_8_bits_uop_uses_ldq = _RANDOM[10'h23F][2];	// lsu.scala:211:16
        stq_8_bits_uop_uses_stq = _RANDOM[10'h23F][3];	// lsu.scala:211:16
        stq_8_bits_uop_is_sys_pc2epc = _RANDOM[10'h23F][4];	// lsu.scala:211:16
        stq_8_bits_uop_is_unique = _RANDOM[10'h23F][5];	// lsu.scala:211:16
        stq_8_bits_uop_flush_on_commit = _RANDOM[10'h23F][6];	// lsu.scala:211:16
        stq_8_bits_uop_ldst_is_rs1 = _RANDOM[10'h23F][7];	// lsu.scala:211:16
        stq_8_bits_uop_ldst = _RANDOM[10'h23F][13:8];	// lsu.scala:211:16
        stq_8_bits_uop_lrs1 = _RANDOM[10'h23F][19:14];	// lsu.scala:211:16
        stq_8_bits_uop_lrs2 = _RANDOM[10'h23F][25:20];	// lsu.scala:211:16
        stq_8_bits_uop_lrs3 = _RANDOM[10'h23F][31:26];	// lsu.scala:211:16
        stq_8_bits_uop_ldst_val = _RANDOM[10'h240][0];	// lsu.scala:211:16
        stq_8_bits_uop_dst_rtype = _RANDOM[10'h240][2:1];	// lsu.scala:211:16
        stq_8_bits_uop_lrs1_rtype = _RANDOM[10'h240][4:3];	// lsu.scala:211:16
        stq_8_bits_uop_lrs2_rtype = _RANDOM[10'h240][6:5];	// lsu.scala:211:16
        stq_8_bits_uop_frs3_en = _RANDOM[10'h240][7];	// lsu.scala:211:16
        stq_8_bits_uop_fp_val = _RANDOM[10'h240][8];	// lsu.scala:211:16
        stq_8_bits_uop_fp_single = _RANDOM[10'h240][9];	// lsu.scala:211:16
        stq_8_bits_uop_xcpt_pf_if = _RANDOM[10'h240][10];	// lsu.scala:211:16
        stq_8_bits_uop_xcpt_ae_if = _RANDOM[10'h240][11];	// lsu.scala:211:16
        stq_8_bits_uop_xcpt_ma_if = _RANDOM[10'h240][12];	// lsu.scala:211:16
        stq_8_bits_uop_bp_debug_if = _RANDOM[10'h240][13];	// lsu.scala:211:16
        stq_8_bits_uop_bp_xcpt_if = _RANDOM[10'h240][14];	// lsu.scala:211:16
        stq_8_bits_uop_debug_fsrc = _RANDOM[10'h240][16:15];	// lsu.scala:211:16
        stq_8_bits_uop_debug_tsrc = _RANDOM[10'h240][18:17];	// lsu.scala:211:16
        stq_8_bits_addr_valid = _RANDOM[10'h240][19];	// lsu.scala:211:16
        stq_8_bits_addr_bits = {_RANDOM[10'h240][31:20], _RANDOM[10'h241][27:0]};	// lsu.scala:211:16
        stq_8_bits_addr_is_virtual = _RANDOM[10'h241][28];	// lsu.scala:211:16
        stq_8_bits_data_valid = _RANDOM[10'h241][29];	// lsu.scala:211:16
        stq_8_bits_data_bits =
          {_RANDOM[10'h241][31:30], _RANDOM[10'h242], _RANDOM[10'h243][29:0]};	// lsu.scala:211:16
        stq_8_bits_committed = _RANDOM[10'h243][30];	// lsu.scala:211:16
        stq_8_bits_succeeded = _RANDOM[10'h243][31];	// lsu.scala:211:16
        stq_9_valid = _RANDOM[10'h246][0];	// lsu.scala:211:16
        stq_9_bits_uop_uopc = _RANDOM[10'h246][7:1];	// lsu.scala:211:16
        stq_9_bits_uop_inst = {_RANDOM[10'h246][31:8], _RANDOM[10'h247][7:0]};	// lsu.scala:211:16
        stq_9_bits_uop_debug_inst = {_RANDOM[10'h247][31:8], _RANDOM[10'h248][7:0]};	// lsu.scala:211:16
        stq_9_bits_uop_is_rvc = _RANDOM[10'h248][8];	// lsu.scala:211:16
        stq_9_bits_uop_debug_pc = {_RANDOM[10'h248][31:9], _RANDOM[10'h249][16:0]};	// lsu.scala:211:16
        stq_9_bits_uop_iq_type = _RANDOM[10'h249][19:17];	// lsu.scala:211:16
        stq_9_bits_uop_fu_code = _RANDOM[10'h249][29:20];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_br_type = {_RANDOM[10'h249][31:30], _RANDOM[10'h24A][1:0]};	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op1_sel = _RANDOM[10'h24A][3:2];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op2_sel = _RANDOM[10'h24A][6:4];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_imm_sel = _RANDOM[10'h24A][9:7];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op_fcn = _RANDOM[10'h24A][13:10];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_fcn_dw = _RANDOM[10'h24A][14];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_csr_cmd = _RANDOM[10'h24A][17:15];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_is_load = _RANDOM[10'h24A][18];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_is_sta = _RANDOM[10'h24A][19];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_is_std = _RANDOM[10'h24A][20];	// lsu.scala:211:16
        stq_9_bits_uop_iw_state = _RANDOM[10'h24A][22:21];	// lsu.scala:211:16
        stq_9_bits_uop_iw_p1_poisoned = _RANDOM[10'h24A][23];	// lsu.scala:211:16
        stq_9_bits_uop_iw_p2_poisoned = _RANDOM[10'h24A][24];	// lsu.scala:211:16
        stq_9_bits_uop_is_br = _RANDOM[10'h24A][25];	// lsu.scala:211:16
        stq_9_bits_uop_is_jalr = _RANDOM[10'h24A][26];	// lsu.scala:211:16
        stq_9_bits_uop_is_jal = _RANDOM[10'h24A][27];	// lsu.scala:211:16
        stq_9_bits_uop_is_sfb = _RANDOM[10'h24A][28];	// lsu.scala:211:16
        stq_9_bits_uop_br_mask = {_RANDOM[10'h24A][31:29], _RANDOM[10'h24B][12:0]};	// lsu.scala:211:16
        stq_9_bits_uop_br_tag = _RANDOM[10'h24B][16:13];	// lsu.scala:211:16
        stq_9_bits_uop_ftq_idx = _RANDOM[10'h24B][21:17];	// lsu.scala:211:16
        stq_9_bits_uop_edge_inst = _RANDOM[10'h24B][22];	// lsu.scala:211:16
        stq_9_bits_uop_pc_lob = _RANDOM[10'h24B][28:23];	// lsu.scala:211:16
        stq_9_bits_uop_taken = _RANDOM[10'h24B][29];	// lsu.scala:211:16
        stq_9_bits_uop_imm_packed = {_RANDOM[10'h24B][31:30], _RANDOM[10'h24C][17:0]};	// lsu.scala:211:16
        stq_9_bits_uop_csr_addr = _RANDOM[10'h24C][29:18];	// lsu.scala:211:16
        stq_9_bits_uop_rob_idx = {_RANDOM[10'h24C][31:30], _RANDOM[10'h24D][4:0]};	// lsu.scala:211:16
        stq_9_bits_uop_ldq_idx = _RANDOM[10'h24D][9:5];	// lsu.scala:211:16
        stq_9_bits_uop_stq_idx = _RANDOM[10'h24D][14:10];	// lsu.scala:211:16
        stq_9_bits_uop_rxq_idx = _RANDOM[10'h24D][16:15];	// lsu.scala:211:16
        stq_9_bits_uop_pdst = _RANDOM[10'h24D][23:17];	// lsu.scala:211:16
        stq_9_bits_uop_prs1 = _RANDOM[10'h24D][30:24];	// lsu.scala:211:16
        stq_9_bits_uop_prs2 = {_RANDOM[10'h24D][31], _RANDOM[10'h24E][5:0]};	// lsu.scala:211:16
        stq_9_bits_uop_prs3 = _RANDOM[10'h24E][12:6];	// lsu.scala:211:16
        stq_9_bits_uop_ppred = _RANDOM[10'h24E][17:13];	// lsu.scala:211:16
        stq_9_bits_uop_prs1_busy = _RANDOM[10'h24E][18];	// lsu.scala:211:16
        stq_9_bits_uop_prs2_busy = _RANDOM[10'h24E][19];	// lsu.scala:211:16
        stq_9_bits_uop_prs3_busy = _RANDOM[10'h24E][20];	// lsu.scala:211:16
        stq_9_bits_uop_ppred_busy = _RANDOM[10'h24E][21];	// lsu.scala:211:16
        stq_9_bits_uop_stale_pdst = _RANDOM[10'h24E][28:22];	// lsu.scala:211:16
        stq_9_bits_uop_exception = _RANDOM[10'h24E][29];	// lsu.scala:211:16
        stq_9_bits_uop_exc_cause =
          {_RANDOM[10'h24E][31:30], _RANDOM[10'h24F], _RANDOM[10'h250][29:0]};	// lsu.scala:211:16
        stq_9_bits_uop_bypassable = _RANDOM[10'h250][30];	// lsu.scala:211:16
        stq_9_bits_uop_mem_cmd = {_RANDOM[10'h250][31], _RANDOM[10'h251][3:0]};	// lsu.scala:211:16
        stq_9_bits_uop_mem_size = _RANDOM[10'h251][5:4];	// lsu.scala:211:16
        stq_9_bits_uop_mem_signed = _RANDOM[10'h251][6];	// lsu.scala:211:16
        stq_9_bits_uop_is_fence = _RANDOM[10'h251][7];	// lsu.scala:211:16
        stq_9_bits_uop_is_fencei = _RANDOM[10'h251][8];	// lsu.scala:211:16
        stq_9_bits_uop_is_amo = _RANDOM[10'h251][9];	// lsu.scala:211:16
        stq_9_bits_uop_uses_ldq = _RANDOM[10'h251][10];	// lsu.scala:211:16
        stq_9_bits_uop_uses_stq = _RANDOM[10'h251][11];	// lsu.scala:211:16
        stq_9_bits_uop_is_sys_pc2epc = _RANDOM[10'h251][12];	// lsu.scala:211:16
        stq_9_bits_uop_is_unique = _RANDOM[10'h251][13];	// lsu.scala:211:16
        stq_9_bits_uop_flush_on_commit = _RANDOM[10'h251][14];	// lsu.scala:211:16
        stq_9_bits_uop_ldst_is_rs1 = _RANDOM[10'h251][15];	// lsu.scala:211:16
        stq_9_bits_uop_ldst = _RANDOM[10'h251][21:16];	// lsu.scala:211:16
        stq_9_bits_uop_lrs1 = _RANDOM[10'h251][27:22];	// lsu.scala:211:16
        stq_9_bits_uop_lrs2 = {_RANDOM[10'h251][31:28], _RANDOM[10'h252][1:0]};	// lsu.scala:211:16
        stq_9_bits_uop_lrs3 = _RANDOM[10'h252][7:2];	// lsu.scala:211:16
        stq_9_bits_uop_ldst_val = _RANDOM[10'h252][8];	// lsu.scala:211:16
        stq_9_bits_uop_dst_rtype = _RANDOM[10'h252][10:9];	// lsu.scala:211:16
        stq_9_bits_uop_lrs1_rtype = _RANDOM[10'h252][12:11];	// lsu.scala:211:16
        stq_9_bits_uop_lrs2_rtype = _RANDOM[10'h252][14:13];	// lsu.scala:211:16
        stq_9_bits_uop_frs3_en = _RANDOM[10'h252][15];	// lsu.scala:211:16
        stq_9_bits_uop_fp_val = _RANDOM[10'h252][16];	// lsu.scala:211:16
        stq_9_bits_uop_fp_single = _RANDOM[10'h252][17];	// lsu.scala:211:16
        stq_9_bits_uop_xcpt_pf_if = _RANDOM[10'h252][18];	// lsu.scala:211:16
        stq_9_bits_uop_xcpt_ae_if = _RANDOM[10'h252][19];	// lsu.scala:211:16
        stq_9_bits_uop_xcpt_ma_if = _RANDOM[10'h252][20];	// lsu.scala:211:16
        stq_9_bits_uop_bp_debug_if = _RANDOM[10'h252][21];	// lsu.scala:211:16
        stq_9_bits_uop_bp_xcpt_if = _RANDOM[10'h252][22];	// lsu.scala:211:16
        stq_9_bits_uop_debug_fsrc = _RANDOM[10'h252][24:23];	// lsu.scala:211:16
        stq_9_bits_uop_debug_tsrc = _RANDOM[10'h252][26:25];	// lsu.scala:211:16
        stq_9_bits_addr_valid = _RANDOM[10'h252][27];	// lsu.scala:211:16
        stq_9_bits_addr_bits =
          {_RANDOM[10'h252][31:28], _RANDOM[10'h253], _RANDOM[10'h254][3:0]};	// lsu.scala:211:16
        stq_9_bits_addr_is_virtual = _RANDOM[10'h254][4];	// lsu.scala:211:16
        stq_9_bits_data_valid = _RANDOM[10'h254][5];	// lsu.scala:211:16
        stq_9_bits_data_bits =
          {_RANDOM[10'h254][31:6], _RANDOM[10'h255], _RANDOM[10'h256][5:0]};	// lsu.scala:211:16
        stq_9_bits_committed = _RANDOM[10'h256][6];	// lsu.scala:211:16
        stq_9_bits_succeeded = _RANDOM[10'h256][7];	// lsu.scala:211:16
        stq_10_valid = _RANDOM[10'h258][8];	// lsu.scala:211:16
        stq_10_bits_uop_uopc = _RANDOM[10'h258][15:9];	// lsu.scala:211:16
        stq_10_bits_uop_inst = {_RANDOM[10'h258][31:16], _RANDOM[10'h259][15:0]};	// lsu.scala:211:16
        stq_10_bits_uop_debug_inst = {_RANDOM[10'h259][31:16], _RANDOM[10'h25A][15:0]};	// lsu.scala:211:16
        stq_10_bits_uop_is_rvc = _RANDOM[10'h25A][16];	// lsu.scala:211:16
        stq_10_bits_uop_debug_pc = {_RANDOM[10'h25A][31:17], _RANDOM[10'h25B][24:0]};	// lsu.scala:211:16
        stq_10_bits_uop_iq_type = _RANDOM[10'h25B][27:25];	// lsu.scala:211:16
        stq_10_bits_uop_fu_code = {_RANDOM[10'h25B][31:28], _RANDOM[10'h25C][5:0]};	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_br_type = _RANDOM[10'h25C][9:6];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op1_sel = _RANDOM[10'h25C][11:10];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op2_sel = _RANDOM[10'h25C][14:12];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_imm_sel = _RANDOM[10'h25C][17:15];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op_fcn = _RANDOM[10'h25C][21:18];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_fcn_dw = _RANDOM[10'h25C][22];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_csr_cmd = _RANDOM[10'h25C][25:23];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_is_load = _RANDOM[10'h25C][26];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_is_sta = _RANDOM[10'h25C][27];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_is_std = _RANDOM[10'h25C][28];	// lsu.scala:211:16
        stq_10_bits_uop_iw_state = _RANDOM[10'h25C][30:29];	// lsu.scala:211:16
        stq_10_bits_uop_iw_p1_poisoned = _RANDOM[10'h25C][31];	// lsu.scala:211:16
        stq_10_bits_uop_iw_p2_poisoned = _RANDOM[10'h25D][0];	// lsu.scala:211:16
        stq_10_bits_uop_is_br = _RANDOM[10'h25D][1];	// lsu.scala:211:16
        stq_10_bits_uop_is_jalr = _RANDOM[10'h25D][2];	// lsu.scala:211:16
        stq_10_bits_uop_is_jal = _RANDOM[10'h25D][3];	// lsu.scala:211:16
        stq_10_bits_uop_is_sfb = _RANDOM[10'h25D][4];	// lsu.scala:211:16
        stq_10_bits_uop_br_mask = _RANDOM[10'h25D][20:5];	// lsu.scala:211:16
        stq_10_bits_uop_br_tag = _RANDOM[10'h25D][24:21];	// lsu.scala:211:16
        stq_10_bits_uop_ftq_idx = _RANDOM[10'h25D][29:25];	// lsu.scala:211:16
        stq_10_bits_uop_edge_inst = _RANDOM[10'h25D][30];	// lsu.scala:211:16
        stq_10_bits_uop_pc_lob = {_RANDOM[10'h25D][31], _RANDOM[10'h25E][4:0]};	// lsu.scala:211:16
        stq_10_bits_uop_taken = _RANDOM[10'h25E][5];	// lsu.scala:211:16
        stq_10_bits_uop_imm_packed = _RANDOM[10'h25E][25:6];	// lsu.scala:211:16
        stq_10_bits_uop_csr_addr = {_RANDOM[10'h25E][31:26], _RANDOM[10'h25F][5:0]};	// lsu.scala:211:16
        stq_10_bits_uop_rob_idx = _RANDOM[10'h25F][12:6];	// lsu.scala:211:16
        stq_10_bits_uop_ldq_idx = _RANDOM[10'h25F][17:13];	// lsu.scala:211:16
        stq_10_bits_uop_stq_idx = _RANDOM[10'h25F][22:18];	// lsu.scala:211:16
        stq_10_bits_uop_rxq_idx = _RANDOM[10'h25F][24:23];	// lsu.scala:211:16
        stq_10_bits_uop_pdst = _RANDOM[10'h25F][31:25];	// lsu.scala:211:16
        stq_10_bits_uop_prs1 = _RANDOM[10'h260][6:0];	// lsu.scala:211:16
        stq_10_bits_uop_prs2 = _RANDOM[10'h260][13:7];	// lsu.scala:211:16
        stq_10_bits_uop_prs3 = _RANDOM[10'h260][20:14];	// lsu.scala:211:16
        stq_10_bits_uop_ppred = _RANDOM[10'h260][25:21];	// lsu.scala:211:16
        stq_10_bits_uop_prs1_busy = _RANDOM[10'h260][26];	// lsu.scala:211:16
        stq_10_bits_uop_prs2_busy = _RANDOM[10'h260][27];	// lsu.scala:211:16
        stq_10_bits_uop_prs3_busy = _RANDOM[10'h260][28];	// lsu.scala:211:16
        stq_10_bits_uop_ppred_busy = _RANDOM[10'h260][29];	// lsu.scala:211:16
        stq_10_bits_uop_stale_pdst = {_RANDOM[10'h260][31:30], _RANDOM[10'h261][4:0]};	// lsu.scala:211:16
        stq_10_bits_uop_exception = _RANDOM[10'h261][5];	// lsu.scala:211:16
        stq_10_bits_uop_exc_cause =
          {_RANDOM[10'h261][31:6], _RANDOM[10'h262], _RANDOM[10'h263][5:0]};	// lsu.scala:211:16
        stq_10_bits_uop_bypassable = _RANDOM[10'h263][6];	// lsu.scala:211:16
        stq_10_bits_uop_mem_cmd = _RANDOM[10'h263][11:7];	// lsu.scala:211:16
        stq_10_bits_uop_mem_size = _RANDOM[10'h263][13:12];	// lsu.scala:211:16
        stq_10_bits_uop_mem_signed = _RANDOM[10'h263][14];	// lsu.scala:211:16
        stq_10_bits_uop_is_fence = _RANDOM[10'h263][15];	// lsu.scala:211:16
        stq_10_bits_uop_is_fencei = _RANDOM[10'h263][16];	// lsu.scala:211:16
        stq_10_bits_uop_is_amo = _RANDOM[10'h263][17];	// lsu.scala:211:16
        stq_10_bits_uop_uses_ldq = _RANDOM[10'h263][18];	// lsu.scala:211:16
        stq_10_bits_uop_uses_stq = _RANDOM[10'h263][19];	// lsu.scala:211:16
        stq_10_bits_uop_is_sys_pc2epc = _RANDOM[10'h263][20];	// lsu.scala:211:16
        stq_10_bits_uop_is_unique = _RANDOM[10'h263][21];	// lsu.scala:211:16
        stq_10_bits_uop_flush_on_commit = _RANDOM[10'h263][22];	// lsu.scala:211:16
        stq_10_bits_uop_ldst_is_rs1 = _RANDOM[10'h263][23];	// lsu.scala:211:16
        stq_10_bits_uop_ldst = _RANDOM[10'h263][29:24];	// lsu.scala:211:16
        stq_10_bits_uop_lrs1 = {_RANDOM[10'h263][31:30], _RANDOM[10'h264][3:0]};	// lsu.scala:211:16
        stq_10_bits_uop_lrs2 = _RANDOM[10'h264][9:4];	// lsu.scala:211:16
        stq_10_bits_uop_lrs3 = _RANDOM[10'h264][15:10];	// lsu.scala:211:16
        stq_10_bits_uop_ldst_val = _RANDOM[10'h264][16];	// lsu.scala:211:16
        stq_10_bits_uop_dst_rtype = _RANDOM[10'h264][18:17];	// lsu.scala:211:16
        stq_10_bits_uop_lrs1_rtype = _RANDOM[10'h264][20:19];	// lsu.scala:211:16
        stq_10_bits_uop_lrs2_rtype = _RANDOM[10'h264][22:21];	// lsu.scala:211:16
        stq_10_bits_uop_frs3_en = _RANDOM[10'h264][23];	// lsu.scala:211:16
        stq_10_bits_uop_fp_val = _RANDOM[10'h264][24];	// lsu.scala:211:16
        stq_10_bits_uop_fp_single = _RANDOM[10'h264][25];	// lsu.scala:211:16
        stq_10_bits_uop_xcpt_pf_if = _RANDOM[10'h264][26];	// lsu.scala:211:16
        stq_10_bits_uop_xcpt_ae_if = _RANDOM[10'h264][27];	// lsu.scala:211:16
        stq_10_bits_uop_xcpt_ma_if = _RANDOM[10'h264][28];	// lsu.scala:211:16
        stq_10_bits_uop_bp_debug_if = _RANDOM[10'h264][29];	// lsu.scala:211:16
        stq_10_bits_uop_bp_xcpt_if = _RANDOM[10'h264][30];	// lsu.scala:211:16
        stq_10_bits_uop_debug_fsrc = {_RANDOM[10'h264][31], _RANDOM[10'h265][0]};	// lsu.scala:211:16
        stq_10_bits_uop_debug_tsrc = _RANDOM[10'h265][2:1];	// lsu.scala:211:16
        stq_10_bits_addr_valid = _RANDOM[10'h265][3];	// lsu.scala:211:16
        stq_10_bits_addr_bits = {_RANDOM[10'h265][31:4], _RANDOM[10'h266][11:0]};	// lsu.scala:211:16
        stq_10_bits_addr_is_virtual = _RANDOM[10'h266][12];	// lsu.scala:211:16
        stq_10_bits_data_valid = _RANDOM[10'h266][13];	// lsu.scala:211:16
        stq_10_bits_data_bits =
          {_RANDOM[10'h266][31:14], _RANDOM[10'h267], _RANDOM[10'h268][13:0]};	// lsu.scala:211:16
        stq_10_bits_committed = _RANDOM[10'h268][14];	// lsu.scala:211:16
        stq_10_bits_succeeded = _RANDOM[10'h268][15];	// lsu.scala:211:16
        stq_11_valid = _RANDOM[10'h26A][16];	// lsu.scala:211:16
        stq_11_bits_uop_uopc = _RANDOM[10'h26A][23:17];	// lsu.scala:211:16
        stq_11_bits_uop_inst = {_RANDOM[10'h26A][31:24], _RANDOM[10'h26B][23:0]};	// lsu.scala:211:16
        stq_11_bits_uop_debug_inst = {_RANDOM[10'h26B][31:24], _RANDOM[10'h26C][23:0]};	// lsu.scala:211:16
        stq_11_bits_uop_is_rvc = _RANDOM[10'h26C][24];	// lsu.scala:211:16
        stq_11_bits_uop_debug_pc =
          {_RANDOM[10'h26C][31:25], _RANDOM[10'h26D], _RANDOM[10'h26E][0]};	// lsu.scala:211:16
        stq_11_bits_uop_iq_type = _RANDOM[10'h26E][3:1];	// lsu.scala:211:16
        stq_11_bits_uop_fu_code = _RANDOM[10'h26E][13:4];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_br_type = _RANDOM[10'h26E][17:14];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op1_sel = _RANDOM[10'h26E][19:18];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op2_sel = _RANDOM[10'h26E][22:20];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_imm_sel = _RANDOM[10'h26E][25:23];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op_fcn = _RANDOM[10'h26E][29:26];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_fcn_dw = _RANDOM[10'h26E][30];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h26E][31], _RANDOM[10'h26F][1:0]};	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_is_load = _RANDOM[10'h26F][2];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_is_sta = _RANDOM[10'h26F][3];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_is_std = _RANDOM[10'h26F][4];	// lsu.scala:211:16
        stq_11_bits_uop_iw_state = _RANDOM[10'h26F][6:5];	// lsu.scala:211:16
        stq_11_bits_uop_iw_p1_poisoned = _RANDOM[10'h26F][7];	// lsu.scala:211:16
        stq_11_bits_uop_iw_p2_poisoned = _RANDOM[10'h26F][8];	// lsu.scala:211:16
        stq_11_bits_uop_is_br = _RANDOM[10'h26F][9];	// lsu.scala:211:16
        stq_11_bits_uop_is_jalr = _RANDOM[10'h26F][10];	// lsu.scala:211:16
        stq_11_bits_uop_is_jal = _RANDOM[10'h26F][11];	// lsu.scala:211:16
        stq_11_bits_uop_is_sfb = _RANDOM[10'h26F][12];	// lsu.scala:211:16
        stq_11_bits_uop_br_mask = _RANDOM[10'h26F][28:13];	// lsu.scala:211:16
        stq_11_bits_uop_br_tag = {_RANDOM[10'h26F][31:29], _RANDOM[10'h270][0]};	// lsu.scala:211:16
        stq_11_bits_uop_ftq_idx = _RANDOM[10'h270][5:1];	// lsu.scala:211:16
        stq_11_bits_uop_edge_inst = _RANDOM[10'h270][6];	// lsu.scala:211:16
        stq_11_bits_uop_pc_lob = _RANDOM[10'h270][12:7];	// lsu.scala:211:16
        stq_11_bits_uop_taken = _RANDOM[10'h270][13];	// lsu.scala:211:16
        stq_11_bits_uop_imm_packed = {_RANDOM[10'h270][31:14], _RANDOM[10'h271][1:0]};	// lsu.scala:211:16
        stq_11_bits_uop_csr_addr = _RANDOM[10'h271][13:2];	// lsu.scala:211:16
        stq_11_bits_uop_rob_idx = _RANDOM[10'h271][20:14];	// lsu.scala:211:16
        stq_11_bits_uop_ldq_idx = _RANDOM[10'h271][25:21];	// lsu.scala:211:16
        stq_11_bits_uop_stq_idx = _RANDOM[10'h271][30:26];	// lsu.scala:211:16
        stq_11_bits_uop_rxq_idx = {_RANDOM[10'h271][31], _RANDOM[10'h272][0]};	// lsu.scala:211:16
        stq_11_bits_uop_pdst = _RANDOM[10'h272][7:1];	// lsu.scala:211:16
        stq_11_bits_uop_prs1 = _RANDOM[10'h272][14:8];	// lsu.scala:211:16
        stq_11_bits_uop_prs2 = _RANDOM[10'h272][21:15];	// lsu.scala:211:16
        stq_11_bits_uop_prs3 = _RANDOM[10'h272][28:22];	// lsu.scala:211:16
        stq_11_bits_uop_ppred = {_RANDOM[10'h272][31:29], _RANDOM[10'h273][1:0]};	// lsu.scala:211:16
        stq_11_bits_uop_prs1_busy = _RANDOM[10'h273][2];	// lsu.scala:211:16
        stq_11_bits_uop_prs2_busy = _RANDOM[10'h273][3];	// lsu.scala:211:16
        stq_11_bits_uop_prs3_busy = _RANDOM[10'h273][4];	// lsu.scala:211:16
        stq_11_bits_uop_ppred_busy = _RANDOM[10'h273][5];	// lsu.scala:211:16
        stq_11_bits_uop_stale_pdst = _RANDOM[10'h273][12:6];	// lsu.scala:211:16
        stq_11_bits_uop_exception = _RANDOM[10'h273][13];	// lsu.scala:211:16
        stq_11_bits_uop_exc_cause =
          {_RANDOM[10'h273][31:14], _RANDOM[10'h274], _RANDOM[10'h275][13:0]};	// lsu.scala:211:16
        stq_11_bits_uop_bypassable = _RANDOM[10'h275][14];	// lsu.scala:211:16
        stq_11_bits_uop_mem_cmd = _RANDOM[10'h275][19:15];	// lsu.scala:211:16
        stq_11_bits_uop_mem_size = _RANDOM[10'h275][21:20];	// lsu.scala:211:16
        stq_11_bits_uop_mem_signed = _RANDOM[10'h275][22];	// lsu.scala:211:16
        stq_11_bits_uop_is_fence = _RANDOM[10'h275][23];	// lsu.scala:211:16
        stq_11_bits_uop_is_fencei = _RANDOM[10'h275][24];	// lsu.scala:211:16
        stq_11_bits_uop_is_amo = _RANDOM[10'h275][25];	// lsu.scala:211:16
        stq_11_bits_uop_uses_ldq = _RANDOM[10'h275][26];	// lsu.scala:211:16
        stq_11_bits_uop_uses_stq = _RANDOM[10'h275][27];	// lsu.scala:211:16
        stq_11_bits_uop_is_sys_pc2epc = _RANDOM[10'h275][28];	// lsu.scala:211:16
        stq_11_bits_uop_is_unique = _RANDOM[10'h275][29];	// lsu.scala:211:16
        stq_11_bits_uop_flush_on_commit = _RANDOM[10'h275][30];	// lsu.scala:211:16
        stq_11_bits_uop_ldst_is_rs1 = _RANDOM[10'h275][31];	// lsu.scala:211:16
        stq_11_bits_uop_ldst = _RANDOM[10'h276][5:0];	// lsu.scala:211:16
        stq_11_bits_uop_lrs1 = _RANDOM[10'h276][11:6];	// lsu.scala:211:16
        stq_11_bits_uop_lrs2 = _RANDOM[10'h276][17:12];	// lsu.scala:211:16
        stq_11_bits_uop_lrs3 = _RANDOM[10'h276][23:18];	// lsu.scala:211:16
        stq_11_bits_uop_ldst_val = _RANDOM[10'h276][24];	// lsu.scala:211:16
        stq_11_bits_uop_dst_rtype = _RANDOM[10'h276][26:25];	// lsu.scala:211:16
        stq_11_bits_uop_lrs1_rtype = _RANDOM[10'h276][28:27];	// lsu.scala:211:16
        stq_11_bits_uop_lrs2_rtype = _RANDOM[10'h276][30:29];	// lsu.scala:211:16
        stq_11_bits_uop_frs3_en = _RANDOM[10'h276][31];	// lsu.scala:211:16
        stq_11_bits_uop_fp_val = _RANDOM[10'h277][0];	// lsu.scala:211:16
        stq_11_bits_uop_fp_single = _RANDOM[10'h277][1];	// lsu.scala:211:16
        stq_11_bits_uop_xcpt_pf_if = _RANDOM[10'h277][2];	// lsu.scala:211:16
        stq_11_bits_uop_xcpt_ae_if = _RANDOM[10'h277][3];	// lsu.scala:211:16
        stq_11_bits_uop_xcpt_ma_if = _RANDOM[10'h277][4];	// lsu.scala:211:16
        stq_11_bits_uop_bp_debug_if = _RANDOM[10'h277][5];	// lsu.scala:211:16
        stq_11_bits_uop_bp_xcpt_if = _RANDOM[10'h277][6];	// lsu.scala:211:16
        stq_11_bits_uop_debug_fsrc = _RANDOM[10'h277][8:7];	// lsu.scala:211:16
        stq_11_bits_uop_debug_tsrc = _RANDOM[10'h277][10:9];	// lsu.scala:211:16
        stq_11_bits_addr_valid = _RANDOM[10'h277][11];	// lsu.scala:211:16
        stq_11_bits_addr_bits = {_RANDOM[10'h277][31:12], _RANDOM[10'h278][19:0]};	// lsu.scala:211:16
        stq_11_bits_addr_is_virtual = _RANDOM[10'h278][20];	// lsu.scala:211:16
        stq_11_bits_data_valid = _RANDOM[10'h278][21];	// lsu.scala:211:16
        stq_11_bits_data_bits =
          {_RANDOM[10'h278][31:22], _RANDOM[10'h279], _RANDOM[10'h27A][21:0]};	// lsu.scala:211:16
        stq_11_bits_committed = _RANDOM[10'h27A][22];	// lsu.scala:211:16
        stq_11_bits_succeeded = _RANDOM[10'h27A][23];	// lsu.scala:211:16
        stq_12_valid = _RANDOM[10'h27C][24];	// lsu.scala:211:16
        stq_12_bits_uop_uopc = _RANDOM[10'h27C][31:25];	// lsu.scala:211:16
        stq_12_bits_uop_inst = _RANDOM[10'h27D];	// lsu.scala:211:16
        stq_12_bits_uop_debug_inst = _RANDOM[10'h27E];	// lsu.scala:211:16
        stq_12_bits_uop_is_rvc = _RANDOM[10'h27F][0];	// lsu.scala:211:16
        stq_12_bits_uop_debug_pc = {_RANDOM[10'h27F][31:1], _RANDOM[10'h280][8:0]};	// lsu.scala:211:16
        stq_12_bits_uop_iq_type = _RANDOM[10'h280][11:9];	// lsu.scala:211:16
        stq_12_bits_uop_fu_code = _RANDOM[10'h280][21:12];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_br_type = _RANDOM[10'h280][25:22];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op1_sel = _RANDOM[10'h280][27:26];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op2_sel = _RANDOM[10'h280][30:28];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_imm_sel = {_RANDOM[10'h280][31], _RANDOM[10'h281][1:0]};	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op_fcn = _RANDOM[10'h281][5:2];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_fcn_dw = _RANDOM[10'h281][6];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_csr_cmd = _RANDOM[10'h281][9:7];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_is_load = _RANDOM[10'h281][10];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_is_sta = _RANDOM[10'h281][11];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_is_std = _RANDOM[10'h281][12];	// lsu.scala:211:16
        stq_12_bits_uop_iw_state = _RANDOM[10'h281][14:13];	// lsu.scala:211:16
        stq_12_bits_uop_iw_p1_poisoned = _RANDOM[10'h281][15];	// lsu.scala:211:16
        stq_12_bits_uop_iw_p2_poisoned = _RANDOM[10'h281][16];	// lsu.scala:211:16
        stq_12_bits_uop_is_br = _RANDOM[10'h281][17];	// lsu.scala:211:16
        stq_12_bits_uop_is_jalr = _RANDOM[10'h281][18];	// lsu.scala:211:16
        stq_12_bits_uop_is_jal = _RANDOM[10'h281][19];	// lsu.scala:211:16
        stq_12_bits_uop_is_sfb = _RANDOM[10'h281][20];	// lsu.scala:211:16
        stq_12_bits_uop_br_mask = {_RANDOM[10'h281][31:21], _RANDOM[10'h282][4:0]};	// lsu.scala:211:16
        stq_12_bits_uop_br_tag = _RANDOM[10'h282][8:5];	// lsu.scala:211:16
        stq_12_bits_uop_ftq_idx = _RANDOM[10'h282][13:9];	// lsu.scala:211:16
        stq_12_bits_uop_edge_inst = _RANDOM[10'h282][14];	// lsu.scala:211:16
        stq_12_bits_uop_pc_lob = _RANDOM[10'h282][20:15];	// lsu.scala:211:16
        stq_12_bits_uop_taken = _RANDOM[10'h282][21];	// lsu.scala:211:16
        stq_12_bits_uop_imm_packed = {_RANDOM[10'h282][31:22], _RANDOM[10'h283][9:0]};	// lsu.scala:211:16
        stq_12_bits_uop_csr_addr = _RANDOM[10'h283][21:10];	// lsu.scala:211:16
        stq_12_bits_uop_rob_idx = _RANDOM[10'h283][28:22];	// lsu.scala:211:16
        stq_12_bits_uop_ldq_idx = {_RANDOM[10'h283][31:29], _RANDOM[10'h284][1:0]};	// lsu.scala:211:16
        stq_12_bits_uop_stq_idx = _RANDOM[10'h284][6:2];	// lsu.scala:211:16
        stq_12_bits_uop_rxq_idx = _RANDOM[10'h284][8:7];	// lsu.scala:211:16
        stq_12_bits_uop_pdst = _RANDOM[10'h284][15:9];	// lsu.scala:211:16
        stq_12_bits_uop_prs1 = _RANDOM[10'h284][22:16];	// lsu.scala:211:16
        stq_12_bits_uop_prs2 = _RANDOM[10'h284][29:23];	// lsu.scala:211:16
        stq_12_bits_uop_prs3 = {_RANDOM[10'h284][31:30], _RANDOM[10'h285][4:0]};	// lsu.scala:211:16
        stq_12_bits_uop_ppred = _RANDOM[10'h285][9:5];	// lsu.scala:211:16
        stq_12_bits_uop_prs1_busy = _RANDOM[10'h285][10];	// lsu.scala:211:16
        stq_12_bits_uop_prs2_busy = _RANDOM[10'h285][11];	// lsu.scala:211:16
        stq_12_bits_uop_prs3_busy = _RANDOM[10'h285][12];	// lsu.scala:211:16
        stq_12_bits_uop_ppred_busy = _RANDOM[10'h285][13];	// lsu.scala:211:16
        stq_12_bits_uop_stale_pdst = _RANDOM[10'h285][20:14];	// lsu.scala:211:16
        stq_12_bits_uop_exception = _RANDOM[10'h285][21];	// lsu.scala:211:16
        stq_12_bits_uop_exc_cause =
          {_RANDOM[10'h285][31:22], _RANDOM[10'h286], _RANDOM[10'h287][21:0]};	// lsu.scala:211:16
        stq_12_bits_uop_bypassable = _RANDOM[10'h287][22];	// lsu.scala:211:16
        stq_12_bits_uop_mem_cmd = _RANDOM[10'h287][27:23];	// lsu.scala:211:16
        stq_12_bits_uop_mem_size = _RANDOM[10'h287][29:28];	// lsu.scala:211:16
        stq_12_bits_uop_mem_signed = _RANDOM[10'h287][30];	// lsu.scala:211:16
        stq_12_bits_uop_is_fence = _RANDOM[10'h287][31];	// lsu.scala:211:16
        stq_12_bits_uop_is_fencei = _RANDOM[10'h288][0];	// lsu.scala:211:16
        stq_12_bits_uop_is_amo = _RANDOM[10'h288][1];	// lsu.scala:211:16
        stq_12_bits_uop_uses_ldq = _RANDOM[10'h288][2];	// lsu.scala:211:16
        stq_12_bits_uop_uses_stq = _RANDOM[10'h288][3];	// lsu.scala:211:16
        stq_12_bits_uop_is_sys_pc2epc = _RANDOM[10'h288][4];	// lsu.scala:211:16
        stq_12_bits_uop_is_unique = _RANDOM[10'h288][5];	// lsu.scala:211:16
        stq_12_bits_uop_flush_on_commit = _RANDOM[10'h288][6];	// lsu.scala:211:16
        stq_12_bits_uop_ldst_is_rs1 = _RANDOM[10'h288][7];	// lsu.scala:211:16
        stq_12_bits_uop_ldst = _RANDOM[10'h288][13:8];	// lsu.scala:211:16
        stq_12_bits_uop_lrs1 = _RANDOM[10'h288][19:14];	// lsu.scala:211:16
        stq_12_bits_uop_lrs2 = _RANDOM[10'h288][25:20];	// lsu.scala:211:16
        stq_12_bits_uop_lrs3 = _RANDOM[10'h288][31:26];	// lsu.scala:211:16
        stq_12_bits_uop_ldst_val = _RANDOM[10'h289][0];	// lsu.scala:211:16
        stq_12_bits_uop_dst_rtype = _RANDOM[10'h289][2:1];	// lsu.scala:211:16
        stq_12_bits_uop_lrs1_rtype = _RANDOM[10'h289][4:3];	// lsu.scala:211:16
        stq_12_bits_uop_lrs2_rtype = _RANDOM[10'h289][6:5];	// lsu.scala:211:16
        stq_12_bits_uop_frs3_en = _RANDOM[10'h289][7];	// lsu.scala:211:16
        stq_12_bits_uop_fp_val = _RANDOM[10'h289][8];	// lsu.scala:211:16
        stq_12_bits_uop_fp_single = _RANDOM[10'h289][9];	// lsu.scala:211:16
        stq_12_bits_uop_xcpt_pf_if = _RANDOM[10'h289][10];	// lsu.scala:211:16
        stq_12_bits_uop_xcpt_ae_if = _RANDOM[10'h289][11];	// lsu.scala:211:16
        stq_12_bits_uop_xcpt_ma_if = _RANDOM[10'h289][12];	// lsu.scala:211:16
        stq_12_bits_uop_bp_debug_if = _RANDOM[10'h289][13];	// lsu.scala:211:16
        stq_12_bits_uop_bp_xcpt_if = _RANDOM[10'h289][14];	// lsu.scala:211:16
        stq_12_bits_uop_debug_fsrc = _RANDOM[10'h289][16:15];	// lsu.scala:211:16
        stq_12_bits_uop_debug_tsrc = _RANDOM[10'h289][18:17];	// lsu.scala:211:16
        stq_12_bits_addr_valid = _RANDOM[10'h289][19];	// lsu.scala:211:16
        stq_12_bits_addr_bits = {_RANDOM[10'h289][31:20], _RANDOM[10'h28A][27:0]};	// lsu.scala:211:16
        stq_12_bits_addr_is_virtual = _RANDOM[10'h28A][28];	// lsu.scala:211:16
        stq_12_bits_data_valid = _RANDOM[10'h28A][29];	// lsu.scala:211:16
        stq_12_bits_data_bits =
          {_RANDOM[10'h28A][31:30], _RANDOM[10'h28B], _RANDOM[10'h28C][29:0]};	// lsu.scala:211:16
        stq_12_bits_committed = _RANDOM[10'h28C][30];	// lsu.scala:211:16
        stq_12_bits_succeeded = _RANDOM[10'h28C][31];	// lsu.scala:211:16
        stq_13_valid = _RANDOM[10'h28F][0];	// lsu.scala:211:16
        stq_13_bits_uop_uopc = _RANDOM[10'h28F][7:1];	// lsu.scala:211:16
        stq_13_bits_uop_inst = {_RANDOM[10'h28F][31:8], _RANDOM[10'h290][7:0]};	// lsu.scala:211:16
        stq_13_bits_uop_debug_inst = {_RANDOM[10'h290][31:8], _RANDOM[10'h291][7:0]};	// lsu.scala:211:16
        stq_13_bits_uop_is_rvc = _RANDOM[10'h291][8];	// lsu.scala:211:16
        stq_13_bits_uop_debug_pc = {_RANDOM[10'h291][31:9], _RANDOM[10'h292][16:0]};	// lsu.scala:211:16
        stq_13_bits_uop_iq_type = _RANDOM[10'h292][19:17];	// lsu.scala:211:16
        stq_13_bits_uop_fu_code = _RANDOM[10'h292][29:20];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_br_type = {_RANDOM[10'h292][31:30], _RANDOM[10'h293][1:0]};	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op1_sel = _RANDOM[10'h293][3:2];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op2_sel = _RANDOM[10'h293][6:4];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_imm_sel = _RANDOM[10'h293][9:7];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op_fcn = _RANDOM[10'h293][13:10];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_fcn_dw = _RANDOM[10'h293][14];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_csr_cmd = _RANDOM[10'h293][17:15];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_is_load = _RANDOM[10'h293][18];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_is_sta = _RANDOM[10'h293][19];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_is_std = _RANDOM[10'h293][20];	// lsu.scala:211:16
        stq_13_bits_uop_iw_state = _RANDOM[10'h293][22:21];	// lsu.scala:211:16
        stq_13_bits_uop_iw_p1_poisoned = _RANDOM[10'h293][23];	// lsu.scala:211:16
        stq_13_bits_uop_iw_p2_poisoned = _RANDOM[10'h293][24];	// lsu.scala:211:16
        stq_13_bits_uop_is_br = _RANDOM[10'h293][25];	// lsu.scala:211:16
        stq_13_bits_uop_is_jalr = _RANDOM[10'h293][26];	// lsu.scala:211:16
        stq_13_bits_uop_is_jal = _RANDOM[10'h293][27];	// lsu.scala:211:16
        stq_13_bits_uop_is_sfb = _RANDOM[10'h293][28];	// lsu.scala:211:16
        stq_13_bits_uop_br_mask = {_RANDOM[10'h293][31:29], _RANDOM[10'h294][12:0]};	// lsu.scala:211:16
        stq_13_bits_uop_br_tag = _RANDOM[10'h294][16:13];	// lsu.scala:211:16
        stq_13_bits_uop_ftq_idx = _RANDOM[10'h294][21:17];	// lsu.scala:211:16
        stq_13_bits_uop_edge_inst = _RANDOM[10'h294][22];	// lsu.scala:211:16
        stq_13_bits_uop_pc_lob = _RANDOM[10'h294][28:23];	// lsu.scala:211:16
        stq_13_bits_uop_taken = _RANDOM[10'h294][29];	// lsu.scala:211:16
        stq_13_bits_uop_imm_packed = {_RANDOM[10'h294][31:30], _RANDOM[10'h295][17:0]};	// lsu.scala:211:16
        stq_13_bits_uop_csr_addr = _RANDOM[10'h295][29:18];	// lsu.scala:211:16
        stq_13_bits_uop_rob_idx = {_RANDOM[10'h295][31:30], _RANDOM[10'h296][4:0]};	// lsu.scala:211:16
        stq_13_bits_uop_ldq_idx = _RANDOM[10'h296][9:5];	// lsu.scala:211:16
        stq_13_bits_uop_stq_idx = _RANDOM[10'h296][14:10];	// lsu.scala:211:16
        stq_13_bits_uop_rxq_idx = _RANDOM[10'h296][16:15];	// lsu.scala:211:16
        stq_13_bits_uop_pdst = _RANDOM[10'h296][23:17];	// lsu.scala:211:16
        stq_13_bits_uop_prs1 = _RANDOM[10'h296][30:24];	// lsu.scala:211:16
        stq_13_bits_uop_prs2 = {_RANDOM[10'h296][31], _RANDOM[10'h297][5:0]};	// lsu.scala:211:16
        stq_13_bits_uop_prs3 = _RANDOM[10'h297][12:6];	// lsu.scala:211:16
        stq_13_bits_uop_ppred = _RANDOM[10'h297][17:13];	// lsu.scala:211:16
        stq_13_bits_uop_prs1_busy = _RANDOM[10'h297][18];	// lsu.scala:211:16
        stq_13_bits_uop_prs2_busy = _RANDOM[10'h297][19];	// lsu.scala:211:16
        stq_13_bits_uop_prs3_busy = _RANDOM[10'h297][20];	// lsu.scala:211:16
        stq_13_bits_uop_ppred_busy = _RANDOM[10'h297][21];	// lsu.scala:211:16
        stq_13_bits_uop_stale_pdst = _RANDOM[10'h297][28:22];	// lsu.scala:211:16
        stq_13_bits_uop_exception = _RANDOM[10'h297][29];	// lsu.scala:211:16
        stq_13_bits_uop_exc_cause =
          {_RANDOM[10'h297][31:30], _RANDOM[10'h298], _RANDOM[10'h299][29:0]};	// lsu.scala:211:16
        stq_13_bits_uop_bypassable = _RANDOM[10'h299][30];	// lsu.scala:211:16
        stq_13_bits_uop_mem_cmd = {_RANDOM[10'h299][31], _RANDOM[10'h29A][3:0]};	// lsu.scala:211:16
        stq_13_bits_uop_mem_size = _RANDOM[10'h29A][5:4];	// lsu.scala:211:16
        stq_13_bits_uop_mem_signed = _RANDOM[10'h29A][6];	// lsu.scala:211:16
        stq_13_bits_uop_is_fence = _RANDOM[10'h29A][7];	// lsu.scala:211:16
        stq_13_bits_uop_is_fencei = _RANDOM[10'h29A][8];	// lsu.scala:211:16
        stq_13_bits_uop_is_amo = _RANDOM[10'h29A][9];	// lsu.scala:211:16
        stq_13_bits_uop_uses_ldq = _RANDOM[10'h29A][10];	// lsu.scala:211:16
        stq_13_bits_uop_uses_stq = _RANDOM[10'h29A][11];	// lsu.scala:211:16
        stq_13_bits_uop_is_sys_pc2epc = _RANDOM[10'h29A][12];	// lsu.scala:211:16
        stq_13_bits_uop_is_unique = _RANDOM[10'h29A][13];	// lsu.scala:211:16
        stq_13_bits_uop_flush_on_commit = _RANDOM[10'h29A][14];	// lsu.scala:211:16
        stq_13_bits_uop_ldst_is_rs1 = _RANDOM[10'h29A][15];	// lsu.scala:211:16
        stq_13_bits_uop_ldst = _RANDOM[10'h29A][21:16];	// lsu.scala:211:16
        stq_13_bits_uop_lrs1 = _RANDOM[10'h29A][27:22];	// lsu.scala:211:16
        stq_13_bits_uop_lrs2 = {_RANDOM[10'h29A][31:28], _RANDOM[10'h29B][1:0]};	// lsu.scala:211:16
        stq_13_bits_uop_lrs3 = _RANDOM[10'h29B][7:2];	// lsu.scala:211:16
        stq_13_bits_uop_ldst_val = _RANDOM[10'h29B][8];	// lsu.scala:211:16
        stq_13_bits_uop_dst_rtype = _RANDOM[10'h29B][10:9];	// lsu.scala:211:16
        stq_13_bits_uop_lrs1_rtype = _RANDOM[10'h29B][12:11];	// lsu.scala:211:16
        stq_13_bits_uop_lrs2_rtype = _RANDOM[10'h29B][14:13];	// lsu.scala:211:16
        stq_13_bits_uop_frs3_en = _RANDOM[10'h29B][15];	// lsu.scala:211:16
        stq_13_bits_uop_fp_val = _RANDOM[10'h29B][16];	// lsu.scala:211:16
        stq_13_bits_uop_fp_single = _RANDOM[10'h29B][17];	// lsu.scala:211:16
        stq_13_bits_uop_xcpt_pf_if = _RANDOM[10'h29B][18];	// lsu.scala:211:16
        stq_13_bits_uop_xcpt_ae_if = _RANDOM[10'h29B][19];	// lsu.scala:211:16
        stq_13_bits_uop_xcpt_ma_if = _RANDOM[10'h29B][20];	// lsu.scala:211:16
        stq_13_bits_uop_bp_debug_if = _RANDOM[10'h29B][21];	// lsu.scala:211:16
        stq_13_bits_uop_bp_xcpt_if = _RANDOM[10'h29B][22];	// lsu.scala:211:16
        stq_13_bits_uop_debug_fsrc = _RANDOM[10'h29B][24:23];	// lsu.scala:211:16
        stq_13_bits_uop_debug_tsrc = _RANDOM[10'h29B][26:25];	// lsu.scala:211:16
        stq_13_bits_addr_valid = _RANDOM[10'h29B][27];	// lsu.scala:211:16
        stq_13_bits_addr_bits =
          {_RANDOM[10'h29B][31:28], _RANDOM[10'h29C], _RANDOM[10'h29D][3:0]};	// lsu.scala:211:16
        stq_13_bits_addr_is_virtual = _RANDOM[10'h29D][4];	// lsu.scala:211:16
        stq_13_bits_data_valid = _RANDOM[10'h29D][5];	// lsu.scala:211:16
        stq_13_bits_data_bits =
          {_RANDOM[10'h29D][31:6], _RANDOM[10'h29E], _RANDOM[10'h29F][5:0]};	// lsu.scala:211:16
        stq_13_bits_committed = _RANDOM[10'h29F][6];	// lsu.scala:211:16
        stq_13_bits_succeeded = _RANDOM[10'h29F][7];	// lsu.scala:211:16
        stq_14_valid = _RANDOM[10'h2A1][8];	// lsu.scala:211:16
        stq_14_bits_uop_uopc = _RANDOM[10'h2A1][15:9];	// lsu.scala:211:16
        stq_14_bits_uop_inst = {_RANDOM[10'h2A1][31:16], _RANDOM[10'h2A2][15:0]};	// lsu.scala:211:16
        stq_14_bits_uop_debug_inst = {_RANDOM[10'h2A2][31:16], _RANDOM[10'h2A3][15:0]};	// lsu.scala:211:16
        stq_14_bits_uop_is_rvc = _RANDOM[10'h2A3][16];	// lsu.scala:211:16
        stq_14_bits_uop_debug_pc = {_RANDOM[10'h2A3][31:17], _RANDOM[10'h2A4][24:0]};	// lsu.scala:211:16
        stq_14_bits_uop_iq_type = _RANDOM[10'h2A4][27:25];	// lsu.scala:211:16
        stq_14_bits_uop_fu_code = {_RANDOM[10'h2A4][31:28], _RANDOM[10'h2A5][5:0]};	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_br_type = _RANDOM[10'h2A5][9:6];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op1_sel = _RANDOM[10'h2A5][11:10];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op2_sel = _RANDOM[10'h2A5][14:12];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_imm_sel = _RANDOM[10'h2A5][17:15];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op_fcn = _RANDOM[10'h2A5][21:18];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_fcn_dw = _RANDOM[10'h2A5][22];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_csr_cmd = _RANDOM[10'h2A5][25:23];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_is_load = _RANDOM[10'h2A5][26];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_is_sta = _RANDOM[10'h2A5][27];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_is_std = _RANDOM[10'h2A5][28];	// lsu.scala:211:16
        stq_14_bits_uop_iw_state = _RANDOM[10'h2A5][30:29];	// lsu.scala:211:16
        stq_14_bits_uop_iw_p1_poisoned = _RANDOM[10'h2A5][31];	// lsu.scala:211:16
        stq_14_bits_uop_iw_p2_poisoned = _RANDOM[10'h2A6][0];	// lsu.scala:211:16
        stq_14_bits_uop_is_br = _RANDOM[10'h2A6][1];	// lsu.scala:211:16
        stq_14_bits_uop_is_jalr = _RANDOM[10'h2A6][2];	// lsu.scala:211:16
        stq_14_bits_uop_is_jal = _RANDOM[10'h2A6][3];	// lsu.scala:211:16
        stq_14_bits_uop_is_sfb = _RANDOM[10'h2A6][4];	// lsu.scala:211:16
        stq_14_bits_uop_br_mask = _RANDOM[10'h2A6][20:5];	// lsu.scala:211:16
        stq_14_bits_uop_br_tag = _RANDOM[10'h2A6][24:21];	// lsu.scala:211:16
        stq_14_bits_uop_ftq_idx = _RANDOM[10'h2A6][29:25];	// lsu.scala:211:16
        stq_14_bits_uop_edge_inst = _RANDOM[10'h2A6][30];	// lsu.scala:211:16
        stq_14_bits_uop_pc_lob = {_RANDOM[10'h2A6][31], _RANDOM[10'h2A7][4:0]};	// lsu.scala:211:16
        stq_14_bits_uop_taken = _RANDOM[10'h2A7][5];	// lsu.scala:211:16
        stq_14_bits_uop_imm_packed = _RANDOM[10'h2A7][25:6];	// lsu.scala:211:16
        stq_14_bits_uop_csr_addr = {_RANDOM[10'h2A7][31:26], _RANDOM[10'h2A8][5:0]};	// lsu.scala:211:16
        stq_14_bits_uop_rob_idx = _RANDOM[10'h2A8][12:6];	// lsu.scala:211:16
        stq_14_bits_uop_ldq_idx = _RANDOM[10'h2A8][17:13];	// lsu.scala:211:16
        stq_14_bits_uop_stq_idx = _RANDOM[10'h2A8][22:18];	// lsu.scala:211:16
        stq_14_bits_uop_rxq_idx = _RANDOM[10'h2A8][24:23];	// lsu.scala:211:16
        stq_14_bits_uop_pdst = _RANDOM[10'h2A8][31:25];	// lsu.scala:211:16
        stq_14_bits_uop_prs1 = _RANDOM[10'h2A9][6:0];	// lsu.scala:211:16
        stq_14_bits_uop_prs2 = _RANDOM[10'h2A9][13:7];	// lsu.scala:211:16
        stq_14_bits_uop_prs3 = _RANDOM[10'h2A9][20:14];	// lsu.scala:211:16
        stq_14_bits_uop_ppred = _RANDOM[10'h2A9][25:21];	// lsu.scala:211:16
        stq_14_bits_uop_prs1_busy = _RANDOM[10'h2A9][26];	// lsu.scala:211:16
        stq_14_bits_uop_prs2_busy = _RANDOM[10'h2A9][27];	// lsu.scala:211:16
        stq_14_bits_uop_prs3_busy = _RANDOM[10'h2A9][28];	// lsu.scala:211:16
        stq_14_bits_uop_ppred_busy = _RANDOM[10'h2A9][29];	// lsu.scala:211:16
        stq_14_bits_uop_stale_pdst = {_RANDOM[10'h2A9][31:30], _RANDOM[10'h2AA][4:0]};	// lsu.scala:211:16
        stq_14_bits_uop_exception = _RANDOM[10'h2AA][5];	// lsu.scala:211:16
        stq_14_bits_uop_exc_cause =
          {_RANDOM[10'h2AA][31:6], _RANDOM[10'h2AB], _RANDOM[10'h2AC][5:0]};	// lsu.scala:211:16
        stq_14_bits_uop_bypassable = _RANDOM[10'h2AC][6];	// lsu.scala:211:16
        stq_14_bits_uop_mem_cmd = _RANDOM[10'h2AC][11:7];	// lsu.scala:211:16
        stq_14_bits_uop_mem_size = _RANDOM[10'h2AC][13:12];	// lsu.scala:211:16
        stq_14_bits_uop_mem_signed = _RANDOM[10'h2AC][14];	// lsu.scala:211:16
        stq_14_bits_uop_is_fence = _RANDOM[10'h2AC][15];	// lsu.scala:211:16
        stq_14_bits_uop_is_fencei = _RANDOM[10'h2AC][16];	// lsu.scala:211:16
        stq_14_bits_uop_is_amo = _RANDOM[10'h2AC][17];	// lsu.scala:211:16
        stq_14_bits_uop_uses_ldq = _RANDOM[10'h2AC][18];	// lsu.scala:211:16
        stq_14_bits_uop_uses_stq = _RANDOM[10'h2AC][19];	// lsu.scala:211:16
        stq_14_bits_uop_is_sys_pc2epc = _RANDOM[10'h2AC][20];	// lsu.scala:211:16
        stq_14_bits_uop_is_unique = _RANDOM[10'h2AC][21];	// lsu.scala:211:16
        stq_14_bits_uop_flush_on_commit = _RANDOM[10'h2AC][22];	// lsu.scala:211:16
        stq_14_bits_uop_ldst_is_rs1 = _RANDOM[10'h2AC][23];	// lsu.scala:211:16
        stq_14_bits_uop_ldst = _RANDOM[10'h2AC][29:24];	// lsu.scala:211:16
        stq_14_bits_uop_lrs1 = {_RANDOM[10'h2AC][31:30], _RANDOM[10'h2AD][3:0]};	// lsu.scala:211:16
        stq_14_bits_uop_lrs2 = _RANDOM[10'h2AD][9:4];	// lsu.scala:211:16
        stq_14_bits_uop_lrs3 = _RANDOM[10'h2AD][15:10];	// lsu.scala:211:16
        stq_14_bits_uop_ldst_val = _RANDOM[10'h2AD][16];	// lsu.scala:211:16
        stq_14_bits_uop_dst_rtype = _RANDOM[10'h2AD][18:17];	// lsu.scala:211:16
        stq_14_bits_uop_lrs1_rtype = _RANDOM[10'h2AD][20:19];	// lsu.scala:211:16
        stq_14_bits_uop_lrs2_rtype = _RANDOM[10'h2AD][22:21];	// lsu.scala:211:16
        stq_14_bits_uop_frs3_en = _RANDOM[10'h2AD][23];	// lsu.scala:211:16
        stq_14_bits_uop_fp_val = _RANDOM[10'h2AD][24];	// lsu.scala:211:16
        stq_14_bits_uop_fp_single = _RANDOM[10'h2AD][25];	// lsu.scala:211:16
        stq_14_bits_uop_xcpt_pf_if = _RANDOM[10'h2AD][26];	// lsu.scala:211:16
        stq_14_bits_uop_xcpt_ae_if = _RANDOM[10'h2AD][27];	// lsu.scala:211:16
        stq_14_bits_uop_xcpt_ma_if = _RANDOM[10'h2AD][28];	// lsu.scala:211:16
        stq_14_bits_uop_bp_debug_if = _RANDOM[10'h2AD][29];	// lsu.scala:211:16
        stq_14_bits_uop_bp_xcpt_if = _RANDOM[10'h2AD][30];	// lsu.scala:211:16
        stq_14_bits_uop_debug_fsrc = {_RANDOM[10'h2AD][31], _RANDOM[10'h2AE][0]};	// lsu.scala:211:16
        stq_14_bits_uop_debug_tsrc = _RANDOM[10'h2AE][2:1];	// lsu.scala:211:16
        stq_14_bits_addr_valid = _RANDOM[10'h2AE][3];	// lsu.scala:211:16
        stq_14_bits_addr_bits = {_RANDOM[10'h2AE][31:4], _RANDOM[10'h2AF][11:0]};	// lsu.scala:211:16
        stq_14_bits_addr_is_virtual = _RANDOM[10'h2AF][12];	// lsu.scala:211:16
        stq_14_bits_data_valid = _RANDOM[10'h2AF][13];	// lsu.scala:211:16
        stq_14_bits_data_bits =
          {_RANDOM[10'h2AF][31:14], _RANDOM[10'h2B0], _RANDOM[10'h2B1][13:0]};	// lsu.scala:211:16
        stq_14_bits_committed = _RANDOM[10'h2B1][14];	// lsu.scala:211:16
        stq_14_bits_succeeded = _RANDOM[10'h2B1][15];	// lsu.scala:211:16
        stq_15_valid = _RANDOM[10'h2B3][16];	// lsu.scala:211:16
        stq_15_bits_uop_uopc = _RANDOM[10'h2B3][23:17];	// lsu.scala:211:16
        stq_15_bits_uop_inst = {_RANDOM[10'h2B3][31:24], _RANDOM[10'h2B4][23:0]};	// lsu.scala:211:16
        stq_15_bits_uop_debug_inst = {_RANDOM[10'h2B4][31:24], _RANDOM[10'h2B5][23:0]};	// lsu.scala:211:16
        stq_15_bits_uop_is_rvc = _RANDOM[10'h2B5][24];	// lsu.scala:211:16
        stq_15_bits_uop_debug_pc =
          {_RANDOM[10'h2B5][31:25], _RANDOM[10'h2B6], _RANDOM[10'h2B7][0]};	// lsu.scala:211:16
        stq_15_bits_uop_iq_type = _RANDOM[10'h2B7][3:1];	// lsu.scala:211:16
        stq_15_bits_uop_fu_code = _RANDOM[10'h2B7][13:4];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_br_type = _RANDOM[10'h2B7][17:14];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op1_sel = _RANDOM[10'h2B7][19:18];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op2_sel = _RANDOM[10'h2B7][22:20];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_imm_sel = _RANDOM[10'h2B7][25:23];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op_fcn = _RANDOM[10'h2B7][29:26];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_fcn_dw = _RANDOM[10'h2B7][30];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h2B7][31], _RANDOM[10'h2B8][1:0]};	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_is_load = _RANDOM[10'h2B8][2];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_is_sta = _RANDOM[10'h2B8][3];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_is_std = _RANDOM[10'h2B8][4];	// lsu.scala:211:16
        stq_15_bits_uop_iw_state = _RANDOM[10'h2B8][6:5];	// lsu.scala:211:16
        stq_15_bits_uop_iw_p1_poisoned = _RANDOM[10'h2B8][7];	// lsu.scala:211:16
        stq_15_bits_uop_iw_p2_poisoned = _RANDOM[10'h2B8][8];	// lsu.scala:211:16
        stq_15_bits_uop_is_br = _RANDOM[10'h2B8][9];	// lsu.scala:211:16
        stq_15_bits_uop_is_jalr = _RANDOM[10'h2B8][10];	// lsu.scala:211:16
        stq_15_bits_uop_is_jal = _RANDOM[10'h2B8][11];	// lsu.scala:211:16
        stq_15_bits_uop_is_sfb = _RANDOM[10'h2B8][12];	// lsu.scala:211:16
        stq_15_bits_uop_br_mask = _RANDOM[10'h2B8][28:13];	// lsu.scala:211:16
        stq_15_bits_uop_br_tag = {_RANDOM[10'h2B8][31:29], _RANDOM[10'h2B9][0]};	// lsu.scala:211:16
        stq_15_bits_uop_ftq_idx = _RANDOM[10'h2B9][5:1];	// lsu.scala:211:16
        stq_15_bits_uop_edge_inst = _RANDOM[10'h2B9][6];	// lsu.scala:211:16
        stq_15_bits_uop_pc_lob = _RANDOM[10'h2B9][12:7];	// lsu.scala:211:16
        stq_15_bits_uop_taken = _RANDOM[10'h2B9][13];	// lsu.scala:211:16
        stq_15_bits_uop_imm_packed = {_RANDOM[10'h2B9][31:14], _RANDOM[10'h2BA][1:0]};	// lsu.scala:211:16
        stq_15_bits_uop_csr_addr = _RANDOM[10'h2BA][13:2];	// lsu.scala:211:16
        stq_15_bits_uop_rob_idx = _RANDOM[10'h2BA][20:14];	// lsu.scala:211:16
        stq_15_bits_uop_ldq_idx = _RANDOM[10'h2BA][25:21];	// lsu.scala:211:16
        stq_15_bits_uop_stq_idx = _RANDOM[10'h2BA][30:26];	// lsu.scala:211:16
        stq_15_bits_uop_rxq_idx = {_RANDOM[10'h2BA][31], _RANDOM[10'h2BB][0]};	// lsu.scala:211:16
        stq_15_bits_uop_pdst = _RANDOM[10'h2BB][7:1];	// lsu.scala:211:16
        stq_15_bits_uop_prs1 = _RANDOM[10'h2BB][14:8];	// lsu.scala:211:16
        stq_15_bits_uop_prs2 = _RANDOM[10'h2BB][21:15];	// lsu.scala:211:16
        stq_15_bits_uop_prs3 = _RANDOM[10'h2BB][28:22];	// lsu.scala:211:16
        stq_15_bits_uop_ppred = {_RANDOM[10'h2BB][31:29], _RANDOM[10'h2BC][1:0]};	// lsu.scala:211:16
        stq_15_bits_uop_prs1_busy = _RANDOM[10'h2BC][2];	// lsu.scala:211:16
        stq_15_bits_uop_prs2_busy = _RANDOM[10'h2BC][3];	// lsu.scala:211:16
        stq_15_bits_uop_prs3_busy = _RANDOM[10'h2BC][4];	// lsu.scala:211:16
        stq_15_bits_uop_ppred_busy = _RANDOM[10'h2BC][5];	// lsu.scala:211:16
        stq_15_bits_uop_stale_pdst = _RANDOM[10'h2BC][12:6];	// lsu.scala:211:16
        stq_15_bits_uop_exception = _RANDOM[10'h2BC][13];	// lsu.scala:211:16
        stq_15_bits_uop_exc_cause =
          {_RANDOM[10'h2BC][31:14], _RANDOM[10'h2BD], _RANDOM[10'h2BE][13:0]};	// lsu.scala:211:16
        stq_15_bits_uop_bypassable = _RANDOM[10'h2BE][14];	// lsu.scala:211:16
        stq_15_bits_uop_mem_cmd = _RANDOM[10'h2BE][19:15];	// lsu.scala:211:16
        stq_15_bits_uop_mem_size = _RANDOM[10'h2BE][21:20];	// lsu.scala:211:16
        stq_15_bits_uop_mem_signed = _RANDOM[10'h2BE][22];	// lsu.scala:211:16
        stq_15_bits_uop_is_fence = _RANDOM[10'h2BE][23];	// lsu.scala:211:16
        stq_15_bits_uop_is_fencei = _RANDOM[10'h2BE][24];	// lsu.scala:211:16
        stq_15_bits_uop_is_amo = _RANDOM[10'h2BE][25];	// lsu.scala:211:16
        stq_15_bits_uop_uses_ldq = _RANDOM[10'h2BE][26];	// lsu.scala:211:16
        stq_15_bits_uop_uses_stq = _RANDOM[10'h2BE][27];	// lsu.scala:211:16
        stq_15_bits_uop_is_sys_pc2epc = _RANDOM[10'h2BE][28];	// lsu.scala:211:16
        stq_15_bits_uop_is_unique = _RANDOM[10'h2BE][29];	// lsu.scala:211:16
        stq_15_bits_uop_flush_on_commit = _RANDOM[10'h2BE][30];	// lsu.scala:211:16
        stq_15_bits_uop_ldst_is_rs1 = _RANDOM[10'h2BE][31];	// lsu.scala:211:16
        stq_15_bits_uop_ldst = _RANDOM[10'h2BF][5:0];	// lsu.scala:211:16
        stq_15_bits_uop_lrs1 = _RANDOM[10'h2BF][11:6];	// lsu.scala:211:16
        stq_15_bits_uop_lrs2 = _RANDOM[10'h2BF][17:12];	// lsu.scala:211:16
        stq_15_bits_uop_lrs3 = _RANDOM[10'h2BF][23:18];	// lsu.scala:211:16
        stq_15_bits_uop_ldst_val = _RANDOM[10'h2BF][24];	// lsu.scala:211:16
        stq_15_bits_uop_dst_rtype = _RANDOM[10'h2BF][26:25];	// lsu.scala:211:16
        stq_15_bits_uop_lrs1_rtype = _RANDOM[10'h2BF][28:27];	// lsu.scala:211:16
        stq_15_bits_uop_lrs2_rtype = _RANDOM[10'h2BF][30:29];	// lsu.scala:211:16
        stq_15_bits_uop_frs3_en = _RANDOM[10'h2BF][31];	// lsu.scala:211:16
        stq_15_bits_uop_fp_val = _RANDOM[10'h2C0][0];	// lsu.scala:211:16
        stq_15_bits_uop_fp_single = _RANDOM[10'h2C0][1];	// lsu.scala:211:16
        stq_15_bits_uop_xcpt_pf_if = _RANDOM[10'h2C0][2];	// lsu.scala:211:16
        stq_15_bits_uop_xcpt_ae_if = _RANDOM[10'h2C0][3];	// lsu.scala:211:16
        stq_15_bits_uop_xcpt_ma_if = _RANDOM[10'h2C0][4];	// lsu.scala:211:16
        stq_15_bits_uop_bp_debug_if = _RANDOM[10'h2C0][5];	// lsu.scala:211:16
        stq_15_bits_uop_bp_xcpt_if = _RANDOM[10'h2C0][6];	// lsu.scala:211:16
        stq_15_bits_uop_debug_fsrc = _RANDOM[10'h2C0][8:7];	// lsu.scala:211:16
        stq_15_bits_uop_debug_tsrc = _RANDOM[10'h2C0][10:9];	// lsu.scala:211:16
        stq_15_bits_addr_valid = _RANDOM[10'h2C0][11];	// lsu.scala:211:16
        stq_15_bits_addr_bits = {_RANDOM[10'h2C0][31:12], _RANDOM[10'h2C1][19:0]};	// lsu.scala:211:16
        stq_15_bits_addr_is_virtual = _RANDOM[10'h2C1][20];	// lsu.scala:211:16
        stq_15_bits_data_valid = _RANDOM[10'h2C1][21];	// lsu.scala:211:16
        stq_15_bits_data_bits =
          {_RANDOM[10'h2C1][31:22], _RANDOM[10'h2C2], _RANDOM[10'h2C3][21:0]};	// lsu.scala:211:16
        stq_15_bits_committed = _RANDOM[10'h2C3][22];	// lsu.scala:211:16
        stq_15_bits_succeeded = _RANDOM[10'h2C3][23];	// lsu.scala:211:16
        stq_16_valid = _RANDOM[10'h2C5][24];	// lsu.scala:211:16
        stq_16_bits_uop_uopc = _RANDOM[10'h2C5][31:25];	// lsu.scala:211:16
        stq_16_bits_uop_inst = _RANDOM[10'h2C6];	// lsu.scala:211:16
        stq_16_bits_uop_debug_inst = _RANDOM[10'h2C7];	// lsu.scala:211:16
        stq_16_bits_uop_is_rvc = _RANDOM[10'h2C8][0];	// lsu.scala:211:16
        stq_16_bits_uop_debug_pc = {_RANDOM[10'h2C8][31:1], _RANDOM[10'h2C9][8:0]};	// lsu.scala:211:16
        stq_16_bits_uop_iq_type = _RANDOM[10'h2C9][11:9];	// lsu.scala:211:16
        stq_16_bits_uop_fu_code = _RANDOM[10'h2C9][21:12];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_br_type = _RANDOM[10'h2C9][25:22];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_op1_sel = _RANDOM[10'h2C9][27:26];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_op2_sel = _RANDOM[10'h2C9][30:28];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_imm_sel = {_RANDOM[10'h2C9][31], _RANDOM[10'h2CA][1:0]};	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_op_fcn = _RANDOM[10'h2CA][5:2];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_fcn_dw = _RANDOM[10'h2CA][6];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_csr_cmd = _RANDOM[10'h2CA][9:7];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_is_load = _RANDOM[10'h2CA][10];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_is_sta = _RANDOM[10'h2CA][11];	// lsu.scala:211:16
        stq_16_bits_uop_ctrl_is_std = _RANDOM[10'h2CA][12];	// lsu.scala:211:16
        stq_16_bits_uop_iw_state = _RANDOM[10'h2CA][14:13];	// lsu.scala:211:16
        stq_16_bits_uop_iw_p1_poisoned = _RANDOM[10'h2CA][15];	// lsu.scala:211:16
        stq_16_bits_uop_iw_p2_poisoned = _RANDOM[10'h2CA][16];	// lsu.scala:211:16
        stq_16_bits_uop_is_br = _RANDOM[10'h2CA][17];	// lsu.scala:211:16
        stq_16_bits_uop_is_jalr = _RANDOM[10'h2CA][18];	// lsu.scala:211:16
        stq_16_bits_uop_is_jal = _RANDOM[10'h2CA][19];	// lsu.scala:211:16
        stq_16_bits_uop_is_sfb = _RANDOM[10'h2CA][20];	// lsu.scala:211:16
        stq_16_bits_uop_br_mask = {_RANDOM[10'h2CA][31:21], _RANDOM[10'h2CB][4:0]};	// lsu.scala:211:16
        stq_16_bits_uop_br_tag = _RANDOM[10'h2CB][8:5];	// lsu.scala:211:16
        stq_16_bits_uop_ftq_idx = _RANDOM[10'h2CB][13:9];	// lsu.scala:211:16
        stq_16_bits_uop_edge_inst = _RANDOM[10'h2CB][14];	// lsu.scala:211:16
        stq_16_bits_uop_pc_lob = _RANDOM[10'h2CB][20:15];	// lsu.scala:211:16
        stq_16_bits_uop_taken = _RANDOM[10'h2CB][21];	// lsu.scala:211:16
        stq_16_bits_uop_imm_packed = {_RANDOM[10'h2CB][31:22], _RANDOM[10'h2CC][9:0]};	// lsu.scala:211:16
        stq_16_bits_uop_csr_addr = _RANDOM[10'h2CC][21:10];	// lsu.scala:211:16
        stq_16_bits_uop_rob_idx = _RANDOM[10'h2CC][28:22];	// lsu.scala:211:16
        stq_16_bits_uop_ldq_idx = {_RANDOM[10'h2CC][31:29], _RANDOM[10'h2CD][1:0]};	// lsu.scala:211:16
        stq_16_bits_uop_stq_idx = _RANDOM[10'h2CD][6:2];	// lsu.scala:211:16
        stq_16_bits_uop_rxq_idx = _RANDOM[10'h2CD][8:7];	// lsu.scala:211:16
        stq_16_bits_uop_pdst = _RANDOM[10'h2CD][15:9];	// lsu.scala:211:16
        stq_16_bits_uop_prs1 = _RANDOM[10'h2CD][22:16];	// lsu.scala:211:16
        stq_16_bits_uop_prs2 = _RANDOM[10'h2CD][29:23];	// lsu.scala:211:16
        stq_16_bits_uop_prs3 = {_RANDOM[10'h2CD][31:30], _RANDOM[10'h2CE][4:0]};	// lsu.scala:211:16
        stq_16_bits_uop_ppred = _RANDOM[10'h2CE][9:5];	// lsu.scala:211:16
        stq_16_bits_uop_prs1_busy = _RANDOM[10'h2CE][10];	// lsu.scala:211:16
        stq_16_bits_uop_prs2_busy = _RANDOM[10'h2CE][11];	// lsu.scala:211:16
        stq_16_bits_uop_prs3_busy = _RANDOM[10'h2CE][12];	// lsu.scala:211:16
        stq_16_bits_uop_ppred_busy = _RANDOM[10'h2CE][13];	// lsu.scala:211:16
        stq_16_bits_uop_stale_pdst = _RANDOM[10'h2CE][20:14];	// lsu.scala:211:16
        stq_16_bits_uop_exception = _RANDOM[10'h2CE][21];	// lsu.scala:211:16
        stq_16_bits_uop_exc_cause =
          {_RANDOM[10'h2CE][31:22], _RANDOM[10'h2CF], _RANDOM[10'h2D0][21:0]};	// lsu.scala:211:16
        stq_16_bits_uop_bypassable = _RANDOM[10'h2D0][22];	// lsu.scala:211:16
        stq_16_bits_uop_mem_cmd = _RANDOM[10'h2D0][27:23];	// lsu.scala:211:16
        stq_16_bits_uop_mem_size = _RANDOM[10'h2D0][29:28];	// lsu.scala:211:16
        stq_16_bits_uop_mem_signed = _RANDOM[10'h2D0][30];	// lsu.scala:211:16
        stq_16_bits_uop_is_fence = _RANDOM[10'h2D0][31];	// lsu.scala:211:16
        stq_16_bits_uop_is_fencei = _RANDOM[10'h2D1][0];	// lsu.scala:211:16
        stq_16_bits_uop_is_amo = _RANDOM[10'h2D1][1];	// lsu.scala:211:16
        stq_16_bits_uop_uses_ldq = _RANDOM[10'h2D1][2];	// lsu.scala:211:16
        stq_16_bits_uop_uses_stq = _RANDOM[10'h2D1][3];	// lsu.scala:211:16
        stq_16_bits_uop_is_sys_pc2epc = _RANDOM[10'h2D1][4];	// lsu.scala:211:16
        stq_16_bits_uop_is_unique = _RANDOM[10'h2D1][5];	// lsu.scala:211:16
        stq_16_bits_uop_flush_on_commit = _RANDOM[10'h2D1][6];	// lsu.scala:211:16
        stq_16_bits_uop_ldst_is_rs1 = _RANDOM[10'h2D1][7];	// lsu.scala:211:16
        stq_16_bits_uop_ldst = _RANDOM[10'h2D1][13:8];	// lsu.scala:211:16
        stq_16_bits_uop_lrs1 = _RANDOM[10'h2D1][19:14];	// lsu.scala:211:16
        stq_16_bits_uop_lrs2 = _RANDOM[10'h2D1][25:20];	// lsu.scala:211:16
        stq_16_bits_uop_lrs3 = _RANDOM[10'h2D1][31:26];	// lsu.scala:211:16
        stq_16_bits_uop_ldst_val = _RANDOM[10'h2D2][0];	// lsu.scala:211:16
        stq_16_bits_uop_dst_rtype = _RANDOM[10'h2D2][2:1];	// lsu.scala:211:16
        stq_16_bits_uop_lrs1_rtype = _RANDOM[10'h2D2][4:3];	// lsu.scala:211:16
        stq_16_bits_uop_lrs2_rtype = _RANDOM[10'h2D2][6:5];	// lsu.scala:211:16
        stq_16_bits_uop_frs3_en = _RANDOM[10'h2D2][7];	// lsu.scala:211:16
        stq_16_bits_uop_fp_val = _RANDOM[10'h2D2][8];	// lsu.scala:211:16
        stq_16_bits_uop_fp_single = _RANDOM[10'h2D2][9];	// lsu.scala:211:16
        stq_16_bits_uop_xcpt_pf_if = _RANDOM[10'h2D2][10];	// lsu.scala:211:16
        stq_16_bits_uop_xcpt_ae_if = _RANDOM[10'h2D2][11];	// lsu.scala:211:16
        stq_16_bits_uop_xcpt_ma_if = _RANDOM[10'h2D2][12];	// lsu.scala:211:16
        stq_16_bits_uop_bp_debug_if = _RANDOM[10'h2D2][13];	// lsu.scala:211:16
        stq_16_bits_uop_bp_xcpt_if = _RANDOM[10'h2D2][14];	// lsu.scala:211:16
        stq_16_bits_uop_debug_fsrc = _RANDOM[10'h2D2][16:15];	// lsu.scala:211:16
        stq_16_bits_uop_debug_tsrc = _RANDOM[10'h2D2][18:17];	// lsu.scala:211:16
        stq_16_bits_addr_valid = _RANDOM[10'h2D2][19];	// lsu.scala:211:16
        stq_16_bits_addr_bits = {_RANDOM[10'h2D2][31:20], _RANDOM[10'h2D3][27:0]};	// lsu.scala:211:16
        stq_16_bits_addr_is_virtual = _RANDOM[10'h2D3][28];	// lsu.scala:211:16
        stq_16_bits_data_valid = _RANDOM[10'h2D3][29];	// lsu.scala:211:16
        stq_16_bits_data_bits =
          {_RANDOM[10'h2D3][31:30], _RANDOM[10'h2D4], _RANDOM[10'h2D5][29:0]};	// lsu.scala:211:16
        stq_16_bits_committed = _RANDOM[10'h2D5][30];	// lsu.scala:211:16
        stq_16_bits_succeeded = _RANDOM[10'h2D5][31];	// lsu.scala:211:16
        stq_17_valid = _RANDOM[10'h2D8][0];	// lsu.scala:211:16
        stq_17_bits_uop_uopc = _RANDOM[10'h2D8][7:1];	// lsu.scala:211:16
        stq_17_bits_uop_inst = {_RANDOM[10'h2D8][31:8], _RANDOM[10'h2D9][7:0]};	// lsu.scala:211:16
        stq_17_bits_uop_debug_inst = {_RANDOM[10'h2D9][31:8], _RANDOM[10'h2DA][7:0]};	// lsu.scala:211:16
        stq_17_bits_uop_is_rvc = _RANDOM[10'h2DA][8];	// lsu.scala:211:16
        stq_17_bits_uop_debug_pc = {_RANDOM[10'h2DA][31:9], _RANDOM[10'h2DB][16:0]};	// lsu.scala:211:16
        stq_17_bits_uop_iq_type = _RANDOM[10'h2DB][19:17];	// lsu.scala:211:16
        stq_17_bits_uop_fu_code = _RANDOM[10'h2DB][29:20];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_br_type = {_RANDOM[10'h2DB][31:30], _RANDOM[10'h2DC][1:0]};	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_op1_sel = _RANDOM[10'h2DC][3:2];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_op2_sel = _RANDOM[10'h2DC][6:4];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_imm_sel = _RANDOM[10'h2DC][9:7];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_op_fcn = _RANDOM[10'h2DC][13:10];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_fcn_dw = _RANDOM[10'h2DC][14];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_csr_cmd = _RANDOM[10'h2DC][17:15];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_is_load = _RANDOM[10'h2DC][18];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_is_sta = _RANDOM[10'h2DC][19];	// lsu.scala:211:16
        stq_17_bits_uop_ctrl_is_std = _RANDOM[10'h2DC][20];	// lsu.scala:211:16
        stq_17_bits_uop_iw_state = _RANDOM[10'h2DC][22:21];	// lsu.scala:211:16
        stq_17_bits_uop_iw_p1_poisoned = _RANDOM[10'h2DC][23];	// lsu.scala:211:16
        stq_17_bits_uop_iw_p2_poisoned = _RANDOM[10'h2DC][24];	// lsu.scala:211:16
        stq_17_bits_uop_is_br = _RANDOM[10'h2DC][25];	// lsu.scala:211:16
        stq_17_bits_uop_is_jalr = _RANDOM[10'h2DC][26];	// lsu.scala:211:16
        stq_17_bits_uop_is_jal = _RANDOM[10'h2DC][27];	// lsu.scala:211:16
        stq_17_bits_uop_is_sfb = _RANDOM[10'h2DC][28];	// lsu.scala:211:16
        stq_17_bits_uop_br_mask = {_RANDOM[10'h2DC][31:29], _RANDOM[10'h2DD][12:0]};	// lsu.scala:211:16
        stq_17_bits_uop_br_tag = _RANDOM[10'h2DD][16:13];	// lsu.scala:211:16
        stq_17_bits_uop_ftq_idx = _RANDOM[10'h2DD][21:17];	// lsu.scala:211:16
        stq_17_bits_uop_edge_inst = _RANDOM[10'h2DD][22];	// lsu.scala:211:16
        stq_17_bits_uop_pc_lob = _RANDOM[10'h2DD][28:23];	// lsu.scala:211:16
        stq_17_bits_uop_taken = _RANDOM[10'h2DD][29];	// lsu.scala:211:16
        stq_17_bits_uop_imm_packed = {_RANDOM[10'h2DD][31:30], _RANDOM[10'h2DE][17:0]};	// lsu.scala:211:16
        stq_17_bits_uop_csr_addr = _RANDOM[10'h2DE][29:18];	// lsu.scala:211:16
        stq_17_bits_uop_rob_idx = {_RANDOM[10'h2DE][31:30], _RANDOM[10'h2DF][4:0]};	// lsu.scala:211:16
        stq_17_bits_uop_ldq_idx = _RANDOM[10'h2DF][9:5];	// lsu.scala:211:16
        stq_17_bits_uop_stq_idx = _RANDOM[10'h2DF][14:10];	// lsu.scala:211:16
        stq_17_bits_uop_rxq_idx = _RANDOM[10'h2DF][16:15];	// lsu.scala:211:16
        stq_17_bits_uop_pdst = _RANDOM[10'h2DF][23:17];	// lsu.scala:211:16
        stq_17_bits_uop_prs1 = _RANDOM[10'h2DF][30:24];	// lsu.scala:211:16
        stq_17_bits_uop_prs2 = {_RANDOM[10'h2DF][31], _RANDOM[10'h2E0][5:0]};	// lsu.scala:211:16
        stq_17_bits_uop_prs3 = _RANDOM[10'h2E0][12:6];	// lsu.scala:211:16
        stq_17_bits_uop_ppred = _RANDOM[10'h2E0][17:13];	// lsu.scala:211:16
        stq_17_bits_uop_prs1_busy = _RANDOM[10'h2E0][18];	// lsu.scala:211:16
        stq_17_bits_uop_prs2_busy = _RANDOM[10'h2E0][19];	// lsu.scala:211:16
        stq_17_bits_uop_prs3_busy = _RANDOM[10'h2E0][20];	// lsu.scala:211:16
        stq_17_bits_uop_ppred_busy = _RANDOM[10'h2E0][21];	// lsu.scala:211:16
        stq_17_bits_uop_stale_pdst = _RANDOM[10'h2E0][28:22];	// lsu.scala:211:16
        stq_17_bits_uop_exception = _RANDOM[10'h2E0][29];	// lsu.scala:211:16
        stq_17_bits_uop_exc_cause =
          {_RANDOM[10'h2E0][31:30], _RANDOM[10'h2E1], _RANDOM[10'h2E2][29:0]};	// lsu.scala:211:16
        stq_17_bits_uop_bypassable = _RANDOM[10'h2E2][30];	// lsu.scala:211:16
        stq_17_bits_uop_mem_cmd = {_RANDOM[10'h2E2][31], _RANDOM[10'h2E3][3:0]};	// lsu.scala:211:16
        stq_17_bits_uop_mem_size = _RANDOM[10'h2E3][5:4];	// lsu.scala:211:16
        stq_17_bits_uop_mem_signed = _RANDOM[10'h2E3][6];	// lsu.scala:211:16
        stq_17_bits_uop_is_fence = _RANDOM[10'h2E3][7];	// lsu.scala:211:16
        stq_17_bits_uop_is_fencei = _RANDOM[10'h2E3][8];	// lsu.scala:211:16
        stq_17_bits_uop_is_amo = _RANDOM[10'h2E3][9];	// lsu.scala:211:16
        stq_17_bits_uop_uses_ldq = _RANDOM[10'h2E3][10];	// lsu.scala:211:16
        stq_17_bits_uop_uses_stq = _RANDOM[10'h2E3][11];	// lsu.scala:211:16
        stq_17_bits_uop_is_sys_pc2epc = _RANDOM[10'h2E3][12];	// lsu.scala:211:16
        stq_17_bits_uop_is_unique = _RANDOM[10'h2E3][13];	// lsu.scala:211:16
        stq_17_bits_uop_flush_on_commit = _RANDOM[10'h2E3][14];	// lsu.scala:211:16
        stq_17_bits_uop_ldst_is_rs1 = _RANDOM[10'h2E3][15];	// lsu.scala:211:16
        stq_17_bits_uop_ldst = _RANDOM[10'h2E3][21:16];	// lsu.scala:211:16
        stq_17_bits_uop_lrs1 = _RANDOM[10'h2E3][27:22];	// lsu.scala:211:16
        stq_17_bits_uop_lrs2 = {_RANDOM[10'h2E3][31:28], _RANDOM[10'h2E4][1:0]};	// lsu.scala:211:16
        stq_17_bits_uop_lrs3 = _RANDOM[10'h2E4][7:2];	// lsu.scala:211:16
        stq_17_bits_uop_ldst_val = _RANDOM[10'h2E4][8];	// lsu.scala:211:16
        stq_17_bits_uop_dst_rtype = _RANDOM[10'h2E4][10:9];	// lsu.scala:211:16
        stq_17_bits_uop_lrs1_rtype = _RANDOM[10'h2E4][12:11];	// lsu.scala:211:16
        stq_17_bits_uop_lrs2_rtype = _RANDOM[10'h2E4][14:13];	// lsu.scala:211:16
        stq_17_bits_uop_frs3_en = _RANDOM[10'h2E4][15];	// lsu.scala:211:16
        stq_17_bits_uop_fp_val = _RANDOM[10'h2E4][16];	// lsu.scala:211:16
        stq_17_bits_uop_fp_single = _RANDOM[10'h2E4][17];	// lsu.scala:211:16
        stq_17_bits_uop_xcpt_pf_if = _RANDOM[10'h2E4][18];	// lsu.scala:211:16
        stq_17_bits_uop_xcpt_ae_if = _RANDOM[10'h2E4][19];	// lsu.scala:211:16
        stq_17_bits_uop_xcpt_ma_if = _RANDOM[10'h2E4][20];	// lsu.scala:211:16
        stq_17_bits_uop_bp_debug_if = _RANDOM[10'h2E4][21];	// lsu.scala:211:16
        stq_17_bits_uop_bp_xcpt_if = _RANDOM[10'h2E4][22];	// lsu.scala:211:16
        stq_17_bits_uop_debug_fsrc = _RANDOM[10'h2E4][24:23];	// lsu.scala:211:16
        stq_17_bits_uop_debug_tsrc = _RANDOM[10'h2E4][26:25];	// lsu.scala:211:16
        stq_17_bits_addr_valid = _RANDOM[10'h2E4][27];	// lsu.scala:211:16
        stq_17_bits_addr_bits =
          {_RANDOM[10'h2E4][31:28], _RANDOM[10'h2E5], _RANDOM[10'h2E6][3:0]};	// lsu.scala:211:16
        stq_17_bits_addr_is_virtual = _RANDOM[10'h2E6][4];	// lsu.scala:211:16
        stq_17_bits_data_valid = _RANDOM[10'h2E6][5];	// lsu.scala:211:16
        stq_17_bits_data_bits =
          {_RANDOM[10'h2E6][31:6], _RANDOM[10'h2E7], _RANDOM[10'h2E8][5:0]};	// lsu.scala:211:16
        stq_17_bits_committed = _RANDOM[10'h2E8][6];	// lsu.scala:211:16
        stq_17_bits_succeeded = _RANDOM[10'h2E8][7];	// lsu.scala:211:16
        stq_18_valid = _RANDOM[10'h2EA][8];	// lsu.scala:211:16
        stq_18_bits_uop_uopc = _RANDOM[10'h2EA][15:9];	// lsu.scala:211:16
        stq_18_bits_uop_inst = {_RANDOM[10'h2EA][31:16], _RANDOM[10'h2EB][15:0]};	// lsu.scala:211:16
        stq_18_bits_uop_debug_inst = {_RANDOM[10'h2EB][31:16], _RANDOM[10'h2EC][15:0]};	// lsu.scala:211:16
        stq_18_bits_uop_is_rvc = _RANDOM[10'h2EC][16];	// lsu.scala:211:16
        stq_18_bits_uop_debug_pc = {_RANDOM[10'h2EC][31:17], _RANDOM[10'h2ED][24:0]};	// lsu.scala:211:16
        stq_18_bits_uop_iq_type = _RANDOM[10'h2ED][27:25];	// lsu.scala:211:16
        stq_18_bits_uop_fu_code = {_RANDOM[10'h2ED][31:28], _RANDOM[10'h2EE][5:0]};	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_br_type = _RANDOM[10'h2EE][9:6];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_op1_sel = _RANDOM[10'h2EE][11:10];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_op2_sel = _RANDOM[10'h2EE][14:12];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_imm_sel = _RANDOM[10'h2EE][17:15];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_op_fcn = _RANDOM[10'h2EE][21:18];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_fcn_dw = _RANDOM[10'h2EE][22];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_csr_cmd = _RANDOM[10'h2EE][25:23];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_is_load = _RANDOM[10'h2EE][26];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_is_sta = _RANDOM[10'h2EE][27];	// lsu.scala:211:16
        stq_18_bits_uop_ctrl_is_std = _RANDOM[10'h2EE][28];	// lsu.scala:211:16
        stq_18_bits_uop_iw_state = _RANDOM[10'h2EE][30:29];	// lsu.scala:211:16
        stq_18_bits_uop_iw_p1_poisoned = _RANDOM[10'h2EE][31];	// lsu.scala:211:16
        stq_18_bits_uop_iw_p2_poisoned = _RANDOM[10'h2EF][0];	// lsu.scala:211:16
        stq_18_bits_uop_is_br = _RANDOM[10'h2EF][1];	// lsu.scala:211:16
        stq_18_bits_uop_is_jalr = _RANDOM[10'h2EF][2];	// lsu.scala:211:16
        stq_18_bits_uop_is_jal = _RANDOM[10'h2EF][3];	// lsu.scala:211:16
        stq_18_bits_uop_is_sfb = _RANDOM[10'h2EF][4];	// lsu.scala:211:16
        stq_18_bits_uop_br_mask = _RANDOM[10'h2EF][20:5];	// lsu.scala:211:16
        stq_18_bits_uop_br_tag = _RANDOM[10'h2EF][24:21];	// lsu.scala:211:16
        stq_18_bits_uop_ftq_idx = _RANDOM[10'h2EF][29:25];	// lsu.scala:211:16
        stq_18_bits_uop_edge_inst = _RANDOM[10'h2EF][30];	// lsu.scala:211:16
        stq_18_bits_uop_pc_lob = {_RANDOM[10'h2EF][31], _RANDOM[10'h2F0][4:0]};	// lsu.scala:211:16
        stq_18_bits_uop_taken = _RANDOM[10'h2F0][5];	// lsu.scala:211:16
        stq_18_bits_uop_imm_packed = _RANDOM[10'h2F0][25:6];	// lsu.scala:211:16
        stq_18_bits_uop_csr_addr = {_RANDOM[10'h2F0][31:26], _RANDOM[10'h2F1][5:0]};	// lsu.scala:211:16
        stq_18_bits_uop_rob_idx = _RANDOM[10'h2F1][12:6];	// lsu.scala:211:16
        stq_18_bits_uop_ldq_idx = _RANDOM[10'h2F1][17:13];	// lsu.scala:211:16
        stq_18_bits_uop_stq_idx = _RANDOM[10'h2F1][22:18];	// lsu.scala:211:16
        stq_18_bits_uop_rxq_idx = _RANDOM[10'h2F1][24:23];	// lsu.scala:211:16
        stq_18_bits_uop_pdst = _RANDOM[10'h2F1][31:25];	// lsu.scala:211:16
        stq_18_bits_uop_prs1 = _RANDOM[10'h2F2][6:0];	// lsu.scala:211:16
        stq_18_bits_uop_prs2 = _RANDOM[10'h2F2][13:7];	// lsu.scala:211:16
        stq_18_bits_uop_prs3 = _RANDOM[10'h2F2][20:14];	// lsu.scala:211:16
        stq_18_bits_uop_ppred = _RANDOM[10'h2F2][25:21];	// lsu.scala:211:16
        stq_18_bits_uop_prs1_busy = _RANDOM[10'h2F2][26];	// lsu.scala:211:16
        stq_18_bits_uop_prs2_busy = _RANDOM[10'h2F2][27];	// lsu.scala:211:16
        stq_18_bits_uop_prs3_busy = _RANDOM[10'h2F2][28];	// lsu.scala:211:16
        stq_18_bits_uop_ppred_busy = _RANDOM[10'h2F2][29];	// lsu.scala:211:16
        stq_18_bits_uop_stale_pdst = {_RANDOM[10'h2F2][31:30], _RANDOM[10'h2F3][4:0]};	// lsu.scala:211:16
        stq_18_bits_uop_exception = _RANDOM[10'h2F3][5];	// lsu.scala:211:16
        stq_18_bits_uop_exc_cause =
          {_RANDOM[10'h2F3][31:6], _RANDOM[10'h2F4], _RANDOM[10'h2F5][5:0]};	// lsu.scala:211:16
        stq_18_bits_uop_bypassable = _RANDOM[10'h2F5][6];	// lsu.scala:211:16
        stq_18_bits_uop_mem_cmd = _RANDOM[10'h2F5][11:7];	// lsu.scala:211:16
        stq_18_bits_uop_mem_size = _RANDOM[10'h2F5][13:12];	// lsu.scala:211:16
        stq_18_bits_uop_mem_signed = _RANDOM[10'h2F5][14];	// lsu.scala:211:16
        stq_18_bits_uop_is_fence = _RANDOM[10'h2F5][15];	// lsu.scala:211:16
        stq_18_bits_uop_is_fencei = _RANDOM[10'h2F5][16];	// lsu.scala:211:16
        stq_18_bits_uop_is_amo = _RANDOM[10'h2F5][17];	// lsu.scala:211:16
        stq_18_bits_uop_uses_ldq = _RANDOM[10'h2F5][18];	// lsu.scala:211:16
        stq_18_bits_uop_uses_stq = _RANDOM[10'h2F5][19];	// lsu.scala:211:16
        stq_18_bits_uop_is_sys_pc2epc = _RANDOM[10'h2F5][20];	// lsu.scala:211:16
        stq_18_bits_uop_is_unique = _RANDOM[10'h2F5][21];	// lsu.scala:211:16
        stq_18_bits_uop_flush_on_commit = _RANDOM[10'h2F5][22];	// lsu.scala:211:16
        stq_18_bits_uop_ldst_is_rs1 = _RANDOM[10'h2F5][23];	// lsu.scala:211:16
        stq_18_bits_uop_ldst = _RANDOM[10'h2F5][29:24];	// lsu.scala:211:16
        stq_18_bits_uop_lrs1 = {_RANDOM[10'h2F5][31:30], _RANDOM[10'h2F6][3:0]};	// lsu.scala:211:16
        stq_18_bits_uop_lrs2 = _RANDOM[10'h2F6][9:4];	// lsu.scala:211:16
        stq_18_bits_uop_lrs3 = _RANDOM[10'h2F6][15:10];	// lsu.scala:211:16
        stq_18_bits_uop_ldst_val = _RANDOM[10'h2F6][16];	// lsu.scala:211:16
        stq_18_bits_uop_dst_rtype = _RANDOM[10'h2F6][18:17];	// lsu.scala:211:16
        stq_18_bits_uop_lrs1_rtype = _RANDOM[10'h2F6][20:19];	// lsu.scala:211:16
        stq_18_bits_uop_lrs2_rtype = _RANDOM[10'h2F6][22:21];	// lsu.scala:211:16
        stq_18_bits_uop_frs3_en = _RANDOM[10'h2F6][23];	// lsu.scala:211:16
        stq_18_bits_uop_fp_val = _RANDOM[10'h2F6][24];	// lsu.scala:211:16
        stq_18_bits_uop_fp_single = _RANDOM[10'h2F6][25];	// lsu.scala:211:16
        stq_18_bits_uop_xcpt_pf_if = _RANDOM[10'h2F6][26];	// lsu.scala:211:16
        stq_18_bits_uop_xcpt_ae_if = _RANDOM[10'h2F6][27];	// lsu.scala:211:16
        stq_18_bits_uop_xcpt_ma_if = _RANDOM[10'h2F6][28];	// lsu.scala:211:16
        stq_18_bits_uop_bp_debug_if = _RANDOM[10'h2F6][29];	// lsu.scala:211:16
        stq_18_bits_uop_bp_xcpt_if = _RANDOM[10'h2F6][30];	// lsu.scala:211:16
        stq_18_bits_uop_debug_fsrc = {_RANDOM[10'h2F6][31], _RANDOM[10'h2F7][0]};	// lsu.scala:211:16
        stq_18_bits_uop_debug_tsrc = _RANDOM[10'h2F7][2:1];	// lsu.scala:211:16
        stq_18_bits_addr_valid = _RANDOM[10'h2F7][3];	// lsu.scala:211:16
        stq_18_bits_addr_bits = {_RANDOM[10'h2F7][31:4], _RANDOM[10'h2F8][11:0]};	// lsu.scala:211:16
        stq_18_bits_addr_is_virtual = _RANDOM[10'h2F8][12];	// lsu.scala:211:16
        stq_18_bits_data_valid = _RANDOM[10'h2F8][13];	// lsu.scala:211:16
        stq_18_bits_data_bits =
          {_RANDOM[10'h2F8][31:14], _RANDOM[10'h2F9], _RANDOM[10'h2FA][13:0]};	// lsu.scala:211:16
        stq_18_bits_committed = _RANDOM[10'h2FA][14];	// lsu.scala:211:16
        stq_18_bits_succeeded = _RANDOM[10'h2FA][15];	// lsu.scala:211:16
        stq_19_valid = _RANDOM[10'h2FC][16];	// lsu.scala:211:16
        stq_19_bits_uop_uopc = _RANDOM[10'h2FC][23:17];	// lsu.scala:211:16
        stq_19_bits_uop_inst = {_RANDOM[10'h2FC][31:24], _RANDOM[10'h2FD][23:0]};	// lsu.scala:211:16
        stq_19_bits_uop_debug_inst = {_RANDOM[10'h2FD][31:24], _RANDOM[10'h2FE][23:0]};	// lsu.scala:211:16
        stq_19_bits_uop_is_rvc = _RANDOM[10'h2FE][24];	// lsu.scala:211:16
        stq_19_bits_uop_debug_pc =
          {_RANDOM[10'h2FE][31:25], _RANDOM[10'h2FF], _RANDOM[10'h300][0]};	// lsu.scala:211:16
        stq_19_bits_uop_iq_type = _RANDOM[10'h300][3:1];	// lsu.scala:211:16
        stq_19_bits_uop_fu_code = _RANDOM[10'h300][13:4];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_br_type = _RANDOM[10'h300][17:14];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_op1_sel = _RANDOM[10'h300][19:18];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_op2_sel = _RANDOM[10'h300][22:20];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_imm_sel = _RANDOM[10'h300][25:23];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_op_fcn = _RANDOM[10'h300][29:26];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_fcn_dw = _RANDOM[10'h300][30];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h300][31], _RANDOM[10'h301][1:0]};	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_is_load = _RANDOM[10'h301][2];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_is_sta = _RANDOM[10'h301][3];	// lsu.scala:211:16
        stq_19_bits_uop_ctrl_is_std = _RANDOM[10'h301][4];	// lsu.scala:211:16
        stq_19_bits_uop_iw_state = _RANDOM[10'h301][6:5];	// lsu.scala:211:16
        stq_19_bits_uop_iw_p1_poisoned = _RANDOM[10'h301][7];	// lsu.scala:211:16
        stq_19_bits_uop_iw_p2_poisoned = _RANDOM[10'h301][8];	// lsu.scala:211:16
        stq_19_bits_uop_is_br = _RANDOM[10'h301][9];	// lsu.scala:211:16
        stq_19_bits_uop_is_jalr = _RANDOM[10'h301][10];	// lsu.scala:211:16
        stq_19_bits_uop_is_jal = _RANDOM[10'h301][11];	// lsu.scala:211:16
        stq_19_bits_uop_is_sfb = _RANDOM[10'h301][12];	// lsu.scala:211:16
        stq_19_bits_uop_br_mask = _RANDOM[10'h301][28:13];	// lsu.scala:211:16
        stq_19_bits_uop_br_tag = {_RANDOM[10'h301][31:29], _RANDOM[10'h302][0]};	// lsu.scala:211:16
        stq_19_bits_uop_ftq_idx = _RANDOM[10'h302][5:1];	// lsu.scala:211:16
        stq_19_bits_uop_edge_inst = _RANDOM[10'h302][6];	// lsu.scala:211:16
        stq_19_bits_uop_pc_lob = _RANDOM[10'h302][12:7];	// lsu.scala:211:16
        stq_19_bits_uop_taken = _RANDOM[10'h302][13];	// lsu.scala:211:16
        stq_19_bits_uop_imm_packed = {_RANDOM[10'h302][31:14], _RANDOM[10'h303][1:0]};	// lsu.scala:211:16
        stq_19_bits_uop_csr_addr = _RANDOM[10'h303][13:2];	// lsu.scala:211:16
        stq_19_bits_uop_rob_idx = _RANDOM[10'h303][20:14];	// lsu.scala:211:16
        stq_19_bits_uop_ldq_idx = _RANDOM[10'h303][25:21];	// lsu.scala:211:16
        stq_19_bits_uop_stq_idx = _RANDOM[10'h303][30:26];	// lsu.scala:211:16
        stq_19_bits_uop_rxq_idx = {_RANDOM[10'h303][31], _RANDOM[10'h304][0]};	// lsu.scala:211:16
        stq_19_bits_uop_pdst = _RANDOM[10'h304][7:1];	// lsu.scala:211:16
        stq_19_bits_uop_prs1 = _RANDOM[10'h304][14:8];	// lsu.scala:211:16
        stq_19_bits_uop_prs2 = _RANDOM[10'h304][21:15];	// lsu.scala:211:16
        stq_19_bits_uop_prs3 = _RANDOM[10'h304][28:22];	// lsu.scala:211:16
        stq_19_bits_uop_ppred = {_RANDOM[10'h304][31:29], _RANDOM[10'h305][1:0]};	// lsu.scala:211:16
        stq_19_bits_uop_prs1_busy = _RANDOM[10'h305][2];	// lsu.scala:211:16
        stq_19_bits_uop_prs2_busy = _RANDOM[10'h305][3];	// lsu.scala:211:16
        stq_19_bits_uop_prs3_busy = _RANDOM[10'h305][4];	// lsu.scala:211:16
        stq_19_bits_uop_ppred_busy = _RANDOM[10'h305][5];	// lsu.scala:211:16
        stq_19_bits_uop_stale_pdst = _RANDOM[10'h305][12:6];	// lsu.scala:211:16
        stq_19_bits_uop_exception = _RANDOM[10'h305][13];	// lsu.scala:211:16
        stq_19_bits_uop_exc_cause =
          {_RANDOM[10'h305][31:14], _RANDOM[10'h306], _RANDOM[10'h307][13:0]};	// lsu.scala:211:16
        stq_19_bits_uop_bypassable = _RANDOM[10'h307][14];	// lsu.scala:211:16
        stq_19_bits_uop_mem_cmd = _RANDOM[10'h307][19:15];	// lsu.scala:211:16
        stq_19_bits_uop_mem_size = _RANDOM[10'h307][21:20];	// lsu.scala:211:16
        stq_19_bits_uop_mem_signed = _RANDOM[10'h307][22];	// lsu.scala:211:16
        stq_19_bits_uop_is_fence = _RANDOM[10'h307][23];	// lsu.scala:211:16
        stq_19_bits_uop_is_fencei = _RANDOM[10'h307][24];	// lsu.scala:211:16
        stq_19_bits_uop_is_amo = _RANDOM[10'h307][25];	// lsu.scala:211:16
        stq_19_bits_uop_uses_ldq = _RANDOM[10'h307][26];	// lsu.scala:211:16
        stq_19_bits_uop_uses_stq = _RANDOM[10'h307][27];	// lsu.scala:211:16
        stq_19_bits_uop_is_sys_pc2epc = _RANDOM[10'h307][28];	// lsu.scala:211:16
        stq_19_bits_uop_is_unique = _RANDOM[10'h307][29];	// lsu.scala:211:16
        stq_19_bits_uop_flush_on_commit = _RANDOM[10'h307][30];	// lsu.scala:211:16
        stq_19_bits_uop_ldst_is_rs1 = _RANDOM[10'h307][31];	// lsu.scala:211:16
        stq_19_bits_uop_ldst = _RANDOM[10'h308][5:0];	// lsu.scala:211:16
        stq_19_bits_uop_lrs1 = _RANDOM[10'h308][11:6];	// lsu.scala:211:16
        stq_19_bits_uop_lrs2 = _RANDOM[10'h308][17:12];	// lsu.scala:211:16
        stq_19_bits_uop_lrs3 = _RANDOM[10'h308][23:18];	// lsu.scala:211:16
        stq_19_bits_uop_ldst_val = _RANDOM[10'h308][24];	// lsu.scala:211:16
        stq_19_bits_uop_dst_rtype = _RANDOM[10'h308][26:25];	// lsu.scala:211:16
        stq_19_bits_uop_lrs1_rtype = _RANDOM[10'h308][28:27];	// lsu.scala:211:16
        stq_19_bits_uop_lrs2_rtype = _RANDOM[10'h308][30:29];	// lsu.scala:211:16
        stq_19_bits_uop_frs3_en = _RANDOM[10'h308][31];	// lsu.scala:211:16
        stq_19_bits_uop_fp_val = _RANDOM[10'h309][0];	// lsu.scala:211:16
        stq_19_bits_uop_fp_single = _RANDOM[10'h309][1];	// lsu.scala:211:16
        stq_19_bits_uop_xcpt_pf_if = _RANDOM[10'h309][2];	// lsu.scala:211:16
        stq_19_bits_uop_xcpt_ae_if = _RANDOM[10'h309][3];	// lsu.scala:211:16
        stq_19_bits_uop_xcpt_ma_if = _RANDOM[10'h309][4];	// lsu.scala:211:16
        stq_19_bits_uop_bp_debug_if = _RANDOM[10'h309][5];	// lsu.scala:211:16
        stq_19_bits_uop_bp_xcpt_if = _RANDOM[10'h309][6];	// lsu.scala:211:16
        stq_19_bits_uop_debug_fsrc = _RANDOM[10'h309][8:7];	// lsu.scala:211:16
        stq_19_bits_uop_debug_tsrc = _RANDOM[10'h309][10:9];	// lsu.scala:211:16
        stq_19_bits_addr_valid = _RANDOM[10'h309][11];	// lsu.scala:211:16
        stq_19_bits_addr_bits = {_RANDOM[10'h309][31:12], _RANDOM[10'h30A][19:0]};	// lsu.scala:211:16
        stq_19_bits_addr_is_virtual = _RANDOM[10'h30A][20];	// lsu.scala:211:16
        stq_19_bits_data_valid = _RANDOM[10'h30A][21];	// lsu.scala:211:16
        stq_19_bits_data_bits =
          {_RANDOM[10'h30A][31:22], _RANDOM[10'h30B], _RANDOM[10'h30C][21:0]};	// lsu.scala:211:16
        stq_19_bits_committed = _RANDOM[10'h30C][22];	// lsu.scala:211:16
        stq_19_bits_succeeded = _RANDOM[10'h30C][23];	// lsu.scala:211:16
        stq_20_valid = _RANDOM[10'h30E][24];	// lsu.scala:211:16
        stq_20_bits_uop_uopc = _RANDOM[10'h30E][31:25];	// lsu.scala:211:16
        stq_20_bits_uop_inst = _RANDOM[10'h30F];	// lsu.scala:211:16
        stq_20_bits_uop_debug_inst = _RANDOM[10'h310];	// lsu.scala:211:16
        stq_20_bits_uop_is_rvc = _RANDOM[10'h311][0];	// lsu.scala:211:16
        stq_20_bits_uop_debug_pc = {_RANDOM[10'h311][31:1], _RANDOM[10'h312][8:0]};	// lsu.scala:211:16
        stq_20_bits_uop_iq_type = _RANDOM[10'h312][11:9];	// lsu.scala:211:16
        stq_20_bits_uop_fu_code = _RANDOM[10'h312][21:12];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_br_type = _RANDOM[10'h312][25:22];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_op1_sel = _RANDOM[10'h312][27:26];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_op2_sel = _RANDOM[10'h312][30:28];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_imm_sel = {_RANDOM[10'h312][31], _RANDOM[10'h313][1:0]};	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_op_fcn = _RANDOM[10'h313][5:2];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_fcn_dw = _RANDOM[10'h313][6];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_csr_cmd = _RANDOM[10'h313][9:7];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_is_load = _RANDOM[10'h313][10];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_is_sta = _RANDOM[10'h313][11];	// lsu.scala:211:16
        stq_20_bits_uop_ctrl_is_std = _RANDOM[10'h313][12];	// lsu.scala:211:16
        stq_20_bits_uop_iw_state = _RANDOM[10'h313][14:13];	// lsu.scala:211:16
        stq_20_bits_uop_iw_p1_poisoned = _RANDOM[10'h313][15];	// lsu.scala:211:16
        stq_20_bits_uop_iw_p2_poisoned = _RANDOM[10'h313][16];	// lsu.scala:211:16
        stq_20_bits_uop_is_br = _RANDOM[10'h313][17];	// lsu.scala:211:16
        stq_20_bits_uop_is_jalr = _RANDOM[10'h313][18];	// lsu.scala:211:16
        stq_20_bits_uop_is_jal = _RANDOM[10'h313][19];	// lsu.scala:211:16
        stq_20_bits_uop_is_sfb = _RANDOM[10'h313][20];	// lsu.scala:211:16
        stq_20_bits_uop_br_mask = {_RANDOM[10'h313][31:21], _RANDOM[10'h314][4:0]};	// lsu.scala:211:16
        stq_20_bits_uop_br_tag = _RANDOM[10'h314][8:5];	// lsu.scala:211:16
        stq_20_bits_uop_ftq_idx = _RANDOM[10'h314][13:9];	// lsu.scala:211:16
        stq_20_bits_uop_edge_inst = _RANDOM[10'h314][14];	// lsu.scala:211:16
        stq_20_bits_uop_pc_lob = _RANDOM[10'h314][20:15];	// lsu.scala:211:16
        stq_20_bits_uop_taken = _RANDOM[10'h314][21];	// lsu.scala:211:16
        stq_20_bits_uop_imm_packed = {_RANDOM[10'h314][31:22], _RANDOM[10'h315][9:0]};	// lsu.scala:211:16
        stq_20_bits_uop_csr_addr = _RANDOM[10'h315][21:10];	// lsu.scala:211:16
        stq_20_bits_uop_rob_idx = _RANDOM[10'h315][28:22];	// lsu.scala:211:16
        stq_20_bits_uop_ldq_idx = {_RANDOM[10'h315][31:29], _RANDOM[10'h316][1:0]};	// lsu.scala:211:16
        stq_20_bits_uop_stq_idx = _RANDOM[10'h316][6:2];	// lsu.scala:211:16
        stq_20_bits_uop_rxq_idx = _RANDOM[10'h316][8:7];	// lsu.scala:211:16
        stq_20_bits_uop_pdst = _RANDOM[10'h316][15:9];	// lsu.scala:211:16
        stq_20_bits_uop_prs1 = _RANDOM[10'h316][22:16];	// lsu.scala:211:16
        stq_20_bits_uop_prs2 = _RANDOM[10'h316][29:23];	// lsu.scala:211:16
        stq_20_bits_uop_prs3 = {_RANDOM[10'h316][31:30], _RANDOM[10'h317][4:0]};	// lsu.scala:211:16
        stq_20_bits_uop_ppred = _RANDOM[10'h317][9:5];	// lsu.scala:211:16
        stq_20_bits_uop_prs1_busy = _RANDOM[10'h317][10];	// lsu.scala:211:16
        stq_20_bits_uop_prs2_busy = _RANDOM[10'h317][11];	// lsu.scala:211:16
        stq_20_bits_uop_prs3_busy = _RANDOM[10'h317][12];	// lsu.scala:211:16
        stq_20_bits_uop_ppred_busy = _RANDOM[10'h317][13];	// lsu.scala:211:16
        stq_20_bits_uop_stale_pdst = _RANDOM[10'h317][20:14];	// lsu.scala:211:16
        stq_20_bits_uop_exception = _RANDOM[10'h317][21];	// lsu.scala:211:16
        stq_20_bits_uop_exc_cause =
          {_RANDOM[10'h317][31:22], _RANDOM[10'h318], _RANDOM[10'h319][21:0]};	// lsu.scala:211:16
        stq_20_bits_uop_bypassable = _RANDOM[10'h319][22];	// lsu.scala:211:16
        stq_20_bits_uop_mem_cmd = _RANDOM[10'h319][27:23];	// lsu.scala:211:16
        stq_20_bits_uop_mem_size = _RANDOM[10'h319][29:28];	// lsu.scala:211:16
        stq_20_bits_uop_mem_signed = _RANDOM[10'h319][30];	// lsu.scala:211:16
        stq_20_bits_uop_is_fence = _RANDOM[10'h319][31];	// lsu.scala:211:16
        stq_20_bits_uop_is_fencei = _RANDOM[10'h31A][0];	// lsu.scala:211:16
        stq_20_bits_uop_is_amo = _RANDOM[10'h31A][1];	// lsu.scala:211:16
        stq_20_bits_uop_uses_ldq = _RANDOM[10'h31A][2];	// lsu.scala:211:16
        stq_20_bits_uop_uses_stq = _RANDOM[10'h31A][3];	// lsu.scala:211:16
        stq_20_bits_uop_is_sys_pc2epc = _RANDOM[10'h31A][4];	// lsu.scala:211:16
        stq_20_bits_uop_is_unique = _RANDOM[10'h31A][5];	// lsu.scala:211:16
        stq_20_bits_uop_flush_on_commit = _RANDOM[10'h31A][6];	// lsu.scala:211:16
        stq_20_bits_uop_ldst_is_rs1 = _RANDOM[10'h31A][7];	// lsu.scala:211:16
        stq_20_bits_uop_ldst = _RANDOM[10'h31A][13:8];	// lsu.scala:211:16
        stq_20_bits_uop_lrs1 = _RANDOM[10'h31A][19:14];	// lsu.scala:211:16
        stq_20_bits_uop_lrs2 = _RANDOM[10'h31A][25:20];	// lsu.scala:211:16
        stq_20_bits_uop_lrs3 = _RANDOM[10'h31A][31:26];	// lsu.scala:211:16
        stq_20_bits_uop_ldst_val = _RANDOM[10'h31B][0];	// lsu.scala:211:16
        stq_20_bits_uop_dst_rtype = _RANDOM[10'h31B][2:1];	// lsu.scala:211:16
        stq_20_bits_uop_lrs1_rtype = _RANDOM[10'h31B][4:3];	// lsu.scala:211:16
        stq_20_bits_uop_lrs2_rtype = _RANDOM[10'h31B][6:5];	// lsu.scala:211:16
        stq_20_bits_uop_frs3_en = _RANDOM[10'h31B][7];	// lsu.scala:211:16
        stq_20_bits_uop_fp_val = _RANDOM[10'h31B][8];	// lsu.scala:211:16
        stq_20_bits_uop_fp_single = _RANDOM[10'h31B][9];	// lsu.scala:211:16
        stq_20_bits_uop_xcpt_pf_if = _RANDOM[10'h31B][10];	// lsu.scala:211:16
        stq_20_bits_uop_xcpt_ae_if = _RANDOM[10'h31B][11];	// lsu.scala:211:16
        stq_20_bits_uop_xcpt_ma_if = _RANDOM[10'h31B][12];	// lsu.scala:211:16
        stq_20_bits_uop_bp_debug_if = _RANDOM[10'h31B][13];	// lsu.scala:211:16
        stq_20_bits_uop_bp_xcpt_if = _RANDOM[10'h31B][14];	// lsu.scala:211:16
        stq_20_bits_uop_debug_fsrc = _RANDOM[10'h31B][16:15];	// lsu.scala:211:16
        stq_20_bits_uop_debug_tsrc = _RANDOM[10'h31B][18:17];	// lsu.scala:211:16
        stq_20_bits_addr_valid = _RANDOM[10'h31B][19];	// lsu.scala:211:16
        stq_20_bits_addr_bits = {_RANDOM[10'h31B][31:20], _RANDOM[10'h31C][27:0]};	// lsu.scala:211:16
        stq_20_bits_addr_is_virtual = _RANDOM[10'h31C][28];	// lsu.scala:211:16
        stq_20_bits_data_valid = _RANDOM[10'h31C][29];	// lsu.scala:211:16
        stq_20_bits_data_bits =
          {_RANDOM[10'h31C][31:30], _RANDOM[10'h31D], _RANDOM[10'h31E][29:0]};	// lsu.scala:211:16
        stq_20_bits_committed = _RANDOM[10'h31E][30];	// lsu.scala:211:16
        stq_20_bits_succeeded = _RANDOM[10'h31E][31];	// lsu.scala:211:16
        stq_21_valid = _RANDOM[10'h321][0];	// lsu.scala:211:16
        stq_21_bits_uop_uopc = _RANDOM[10'h321][7:1];	// lsu.scala:211:16
        stq_21_bits_uop_inst = {_RANDOM[10'h321][31:8], _RANDOM[10'h322][7:0]};	// lsu.scala:211:16
        stq_21_bits_uop_debug_inst = {_RANDOM[10'h322][31:8], _RANDOM[10'h323][7:0]};	// lsu.scala:211:16
        stq_21_bits_uop_is_rvc = _RANDOM[10'h323][8];	// lsu.scala:211:16
        stq_21_bits_uop_debug_pc = {_RANDOM[10'h323][31:9], _RANDOM[10'h324][16:0]};	// lsu.scala:211:16
        stq_21_bits_uop_iq_type = _RANDOM[10'h324][19:17];	// lsu.scala:211:16
        stq_21_bits_uop_fu_code = _RANDOM[10'h324][29:20];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_br_type = {_RANDOM[10'h324][31:30], _RANDOM[10'h325][1:0]};	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_op1_sel = _RANDOM[10'h325][3:2];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_op2_sel = _RANDOM[10'h325][6:4];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_imm_sel = _RANDOM[10'h325][9:7];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_op_fcn = _RANDOM[10'h325][13:10];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_fcn_dw = _RANDOM[10'h325][14];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_csr_cmd = _RANDOM[10'h325][17:15];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_is_load = _RANDOM[10'h325][18];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_is_sta = _RANDOM[10'h325][19];	// lsu.scala:211:16
        stq_21_bits_uop_ctrl_is_std = _RANDOM[10'h325][20];	// lsu.scala:211:16
        stq_21_bits_uop_iw_state = _RANDOM[10'h325][22:21];	// lsu.scala:211:16
        stq_21_bits_uop_iw_p1_poisoned = _RANDOM[10'h325][23];	// lsu.scala:211:16
        stq_21_bits_uop_iw_p2_poisoned = _RANDOM[10'h325][24];	// lsu.scala:211:16
        stq_21_bits_uop_is_br = _RANDOM[10'h325][25];	// lsu.scala:211:16
        stq_21_bits_uop_is_jalr = _RANDOM[10'h325][26];	// lsu.scala:211:16
        stq_21_bits_uop_is_jal = _RANDOM[10'h325][27];	// lsu.scala:211:16
        stq_21_bits_uop_is_sfb = _RANDOM[10'h325][28];	// lsu.scala:211:16
        stq_21_bits_uop_br_mask = {_RANDOM[10'h325][31:29], _RANDOM[10'h326][12:0]};	// lsu.scala:211:16
        stq_21_bits_uop_br_tag = _RANDOM[10'h326][16:13];	// lsu.scala:211:16
        stq_21_bits_uop_ftq_idx = _RANDOM[10'h326][21:17];	// lsu.scala:211:16
        stq_21_bits_uop_edge_inst = _RANDOM[10'h326][22];	// lsu.scala:211:16
        stq_21_bits_uop_pc_lob = _RANDOM[10'h326][28:23];	// lsu.scala:211:16
        stq_21_bits_uop_taken = _RANDOM[10'h326][29];	// lsu.scala:211:16
        stq_21_bits_uop_imm_packed = {_RANDOM[10'h326][31:30], _RANDOM[10'h327][17:0]};	// lsu.scala:211:16
        stq_21_bits_uop_csr_addr = _RANDOM[10'h327][29:18];	// lsu.scala:211:16
        stq_21_bits_uop_rob_idx = {_RANDOM[10'h327][31:30], _RANDOM[10'h328][4:0]};	// lsu.scala:211:16
        stq_21_bits_uop_ldq_idx = _RANDOM[10'h328][9:5];	// lsu.scala:211:16
        stq_21_bits_uop_stq_idx = _RANDOM[10'h328][14:10];	// lsu.scala:211:16
        stq_21_bits_uop_rxq_idx = _RANDOM[10'h328][16:15];	// lsu.scala:211:16
        stq_21_bits_uop_pdst = _RANDOM[10'h328][23:17];	// lsu.scala:211:16
        stq_21_bits_uop_prs1 = _RANDOM[10'h328][30:24];	// lsu.scala:211:16
        stq_21_bits_uop_prs2 = {_RANDOM[10'h328][31], _RANDOM[10'h329][5:0]};	// lsu.scala:211:16
        stq_21_bits_uop_prs3 = _RANDOM[10'h329][12:6];	// lsu.scala:211:16
        stq_21_bits_uop_ppred = _RANDOM[10'h329][17:13];	// lsu.scala:211:16
        stq_21_bits_uop_prs1_busy = _RANDOM[10'h329][18];	// lsu.scala:211:16
        stq_21_bits_uop_prs2_busy = _RANDOM[10'h329][19];	// lsu.scala:211:16
        stq_21_bits_uop_prs3_busy = _RANDOM[10'h329][20];	// lsu.scala:211:16
        stq_21_bits_uop_ppred_busy = _RANDOM[10'h329][21];	// lsu.scala:211:16
        stq_21_bits_uop_stale_pdst = _RANDOM[10'h329][28:22];	// lsu.scala:211:16
        stq_21_bits_uop_exception = _RANDOM[10'h329][29];	// lsu.scala:211:16
        stq_21_bits_uop_exc_cause =
          {_RANDOM[10'h329][31:30], _RANDOM[10'h32A], _RANDOM[10'h32B][29:0]};	// lsu.scala:211:16
        stq_21_bits_uop_bypassable = _RANDOM[10'h32B][30];	// lsu.scala:211:16
        stq_21_bits_uop_mem_cmd = {_RANDOM[10'h32B][31], _RANDOM[10'h32C][3:0]};	// lsu.scala:211:16
        stq_21_bits_uop_mem_size = _RANDOM[10'h32C][5:4];	// lsu.scala:211:16
        stq_21_bits_uop_mem_signed = _RANDOM[10'h32C][6];	// lsu.scala:211:16
        stq_21_bits_uop_is_fence = _RANDOM[10'h32C][7];	// lsu.scala:211:16
        stq_21_bits_uop_is_fencei = _RANDOM[10'h32C][8];	// lsu.scala:211:16
        stq_21_bits_uop_is_amo = _RANDOM[10'h32C][9];	// lsu.scala:211:16
        stq_21_bits_uop_uses_ldq = _RANDOM[10'h32C][10];	// lsu.scala:211:16
        stq_21_bits_uop_uses_stq = _RANDOM[10'h32C][11];	// lsu.scala:211:16
        stq_21_bits_uop_is_sys_pc2epc = _RANDOM[10'h32C][12];	// lsu.scala:211:16
        stq_21_bits_uop_is_unique = _RANDOM[10'h32C][13];	// lsu.scala:211:16
        stq_21_bits_uop_flush_on_commit = _RANDOM[10'h32C][14];	// lsu.scala:211:16
        stq_21_bits_uop_ldst_is_rs1 = _RANDOM[10'h32C][15];	// lsu.scala:211:16
        stq_21_bits_uop_ldst = _RANDOM[10'h32C][21:16];	// lsu.scala:211:16
        stq_21_bits_uop_lrs1 = _RANDOM[10'h32C][27:22];	// lsu.scala:211:16
        stq_21_bits_uop_lrs2 = {_RANDOM[10'h32C][31:28], _RANDOM[10'h32D][1:0]};	// lsu.scala:211:16
        stq_21_bits_uop_lrs3 = _RANDOM[10'h32D][7:2];	// lsu.scala:211:16
        stq_21_bits_uop_ldst_val = _RANDOM[10'h32D][8];	// lsu.scala:211:16
        stq_21_bits_uop_dst_rtype = _RANDOM[10'h32D][10:9];	// lsu.scala:211:16
        stq_21_bits_uop_lrs1_rtype = _RANDOM[10'h32D][12:11];	// lsu.scala:211:16
        stq_21_bits_uop_lrs2_rtype = _RANDOM[10'h32D][14:13];	// lsu.scala:211:16
        stq_21_bits_uop_frs3_en = _RANDOM[10'h32D][15];	// lsu.scala:211:16
        stq_21_bits_uop_fp_val = _RANDOM[10'h32D][16];	// lsu.scala:211:16
        stq_21_bits_uop_fp_single = _RANDOM[10'h32D][17];	// lsu.scala:211:16
        stq_21_bits_uop_xcpt_pf_if = _RANDOM[10'h32D][18];	// lsu.scala:211:16
        stq_21_bits_uop_xcpt_ae_if = _RANDOM[10'h32D][19];	// lsu.scala:211:16
        stq_21_bits_uop_xcpt_ma_if = _RANDOM[10'h32D][20];	// lsu.scala:211:16
        stq_21_bits_uop_bp_debug_if = _RANDOM[10'h32D][21];	// lsu.scala:211:16
        stq_21_bits_uop_bp_xcpt_if = _RANDOM[10'h32D][22];	// lsu.scala:211:16
        stq_21_bits_uop_debug_fsrc = _RANDOM[10'h32D][24:23];	// lsu.scala:211:16
        stq_21_bits_uop_debug_tsrc = _RANDOM[10'h32D][26:25];	// lsu.scala:211:16
        stq_21_bits_addr_valid = _RANDOM[10'h32D][27];	// lsu.scala:211:16
        stq_21_bits_addr_bits =
          {_RANDOM[10'h32D][31:28], _RANDOM[10'h32E], _RANDOM[10'h32F][3:0]};	// lsu.scala:211:16
        stq_21_bits_addr_is_virtual = _RANDOM[10'h32F][4];	// lsu.scala:211:16
        stq_21_bits_data_valid = _RANDOM[10'h32F][5];	// lsu.scala:211:16
        stq_21_bits_data_bits =
          {_RANDOM[10'h32F][31:6], _RANDOM[10'h330], _RANDOM[10'h331][5:0]};	// lsu.scala:211:16
        stq_21_bits_committed = _RANDOM[10'h331][6];	// lsu.scala:211:16
        stq_21_bits_succeeded = _RANDOM[10'h331][7];	// lsu.scala:211:16
        stq_22_valid = _RANDOM[10'h333][8];	// lsu.scala:211:16
        stq_22_bits_uop_uopc = _RANDOM[10'h333][15:9];	// lsu.scala:211:16
        stq_22_bits_uop_inst = {_RANDOM[10'h333][31:16], _RANDOM[10'h334][15:0]};	// lsu.scala:211:16
        stq_22_bits_uop_debug_inst = {_RANDOM[10'h334][31:16], _RANDOM[10'h335][15:0]};	// lsu.scala:211:16
        stq_22_bits_uop_is_rvc = _RANDOM[10'h335][16];	// lsu.scala:211:16
        stq_22_bits_uop_debug_pc = {_RANDOM[10'h335][31:17], _RANDOM[10'h336][24:0]};	// lsu.scala:211:16
        stq_22_bits_uop_iq_type = _RANDOM[10'h336][27:25];	// lsu.scala:211:16
        stq_22_bits_uop_fu_code = {_RANDOM[10'h336][31:28], _RANDOM[10'h337][5:0]};	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_br_type = _RANDOM[10'h337][9:6];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_op1_sel = _RANDOM[10'h337][11:10];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_op2_sel = _RANDOM[10'h337][14:12];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_imm_sel = _RANDOM[10'h337][17:15];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_op_fcn = _RANDOM[10'h337][21:18];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_fcn_dw = _RANDOM[10'h337][22];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_csr_cmd = _RANDOM[10'h337][25:23];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_is_load = _RANDOM[10'h337][26];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_is_sta = _RANDOM[10'h337][27];	// lsu.scala:211:16
        stq_22_bits_uop_ctrl_is_std = _RANDOM[10'h337][28];	// lsu.scala:211:16
        stq_22_bits_uop_iw_state = _RANDOM[10'h337][30:29];	// lsu.scala:211:16
        stq_22_bits_uop_iw_p1_poisoned = _RANDOM[10'h337][31];	// lsu.scala:211:16
        stq_22_bits_uop_iw_p2_poisoned = _RANDOM[10'h338][0];	// lsu.scala:211:16
        stq_22_bits_uop_is_br = _RANDOM[10'h338][1];	// lsu.scala:211:16
        stq_22_bits_uop_is_jalr = _RANDOM[10'h338][2];	// lsu.scala:211:16
        stq_22_bits_uop_is_jal = _RANDOM[10'h338][3];	// lsu.scala:211:16
        stq_22_bits_uop_is_sfb = _RANDOM[10'h338][4];	// lsu.scala:211:16
        stq_22_bits_uop_br_mask = _RANDOM[10'h338][20:5];	// lsu.scala:211:16
        stq_22_bits_uop_br_tag = _RANDOM[10'h338][24:21];	// lsu.scala:211:16
        stq_22_bits_uop_ftq_idx = _RANDOM[10'h338][29:25];	// lsu.scala:211:16
        stq_22_bits_uop_edge_inst = _RANDOM[10'h338][30];	// lsu.scala:211:16
        stq_22_bits_uop_pc_lob = {_RANDOM[10'h338][31], _RANDOM[10'h339][4:0]};	// lsu.scala:211:16
        stq_22_bits_uop_taken = _RANDOM[10'h339][5];	// lsu.scala:211:16
        stq_22_bits_uop_imm_packed = _RANDOM[10'h339][25:6];	// lsu.scala:211:16
        stq_22_bits_uop_csr_addr = {_RANDOM[10'h339][31:26], _RANDOM[10'h33A][5:0]};	// lsu.scala:211:16
        stq_22_bits_uop_rob_idx = _RANDOM[10'h33A][12:6];	// lsu.scala:211:16
        stq_22_bits_uop_ldq_idx = _RANDOM[10'h33A][17:13];	// lsu.scala:211:16
        stq_22_bits_uop_stq_idx = _RANDOM[10'h33A][22:18];	// lsu.scala:211:16
        stq_22_bits_uop_rxq_idx = _RANDOM[10'h33A][24:23];	// lsu.scala:211:16
        stq_22_bits_uop_pdst = _RANDOM[10'h33A][31:25];	// lsu.scala:211:16
        stq_22_bits_uop_prs1 = _RANDOM[10'h33B][6:0];	// lsu.scala:211:16
        stq_22_bits_uop_prs2 = _RANDOM[10'h33B][13:7];	// lsu.scala:211:16
        stq_22_bits_uop_prs3 = _RANDOM[10'h33B][20:14];	// lsu.scala:211:16
        stq_22_bits_uop_ppred = _RANDOM[10'h33B][25:21];	// lsu.scala:211:16
        stq_22_bits_uop_prs1_busy = _RANDOM[10'h33B][26];	// lsu.scala:211:16
        stq_22_bits_uop_prs2_busy = _RANDOM[10'h33B][27];	// lsu.scala:211:16
        stq_22_bits_uop_prs3_busy = _RANDOM[10'h33B][28];	// lsu.scala:211:16
        stq_22_bits_uop_ppred_busy = _RANDOM[10'h33B][29];	// lsu.scala:211:16
        stq_22_bits_uop_stale_pdst = {_RANDOM[10'h33B][31:30], _RANDOM[10'h33C][4:0]};	// lsu.scala:211:16
        stq_22_bits_uop_exception = _RANDOM[10'h33C][5];	// lsu.scala:211:16
        stq_22_bits_uop_exc_cause =
          {_RANDOM[10'h33C][31:6], _RANDOM[10'h33D], _RANDOM[10'h33E][5:0]};	// lsu.scala:211:16
        stq_22_bits_uop_bypassable = _RANDOM[10'h33E][6];	// lsu.scala:211:16
        stq_22_bits_uop_mem_cmd = _RANDOM[10'h33E][11:7];	// lsu.scala:211:16
        stq_22_bits_uop_mem_size = _RANDOM[10'h33E][13:12];	// lsu.scala:211:16
        stq_22_bits_uop_mem_signed = _RANDOM[10'h33E][14];	// lsu.scala:211:16
        stq_22_bits_uop_is_fence = _RANDOM[10'h33E][15];	// lsu.scala:211:16
        stq_22_bits_uop_is_fencei = _RANDOM[10'h33E][16];	// lsu.scala:211:16
        stq_22_bits_uop_is_amo = _RANDOM[10'h33E][17];	// lsu.scala:211:16
        stq_22_bits_uop_uses_ldq = _RANDOM[10'h33E][18];	// lsu.scala:211:16
        stq_22_bits_uop_uses_stq = _RANDOM[10'h33E][19];	// lsu.scala:211:16
        stq_22_bits_uop_is_sys_pc2epc = _RANDOM[10'h33E][20];	// lsu.scala:211:16
        stq_22_bits_uop_is_unique = _RANDOM[10'h33E][21];	// lsu.scala:211:16
        stq_22_bits_uop_flush_on_commit = _RANDOM[10'h33E][22];	// lsu.scala:211:16
        stq_22_bits_uop_ldst_is_rs1 = _RANDOM[10'h33E][23];	// lsu.scala:211:16
        stq_22_bits_uop_ldst = _RANDOM[10'h33E][29:24];	// lsu.scala:211:16
        stq_22_bits_uop_lrs1 = {_RANDOM[10'h33E][31:30], _RANDOM[10'h33F][3:0]};	// lsu.scala:211:16
        stq_22_bits_uop_lrs2 = _RANDOM[10'h33F][9:4];	// lsu.scala:211:16
        stq_22_bits_uop_lrs3 = _RANDOM[10'h33F][15:10];	// lsu.scala:211:16
        stq_22_bits_uop_ldst_val = _RANDOM[10'h33F][16];	// lsu.scala:211:16
        stq_22_bits_uop_dst_rtype = _RANDOM[10'h33F][18:17];	// lsu.scala:211:16
        stq_22_bits_uop_lrs1_rtype = _RANDOM[10'h33F][20:19];	// lsu.scala:211:16
        stq_22_bits_uop_lrs2_rtype = _RANDOM[10'h33F][22:21];	// lsu.scala:211:16
        stq_22_bits_uop_frs3_en = _RANDOM[10'h33F][23];	// lsu.scala:211:16
        stq_22_bits_uop_fp_val = _RANDOM[10'h33F][24];	// lsu.scala:211:16
        stq_22_bits_uop_fp_single = _RANDOM[10'h33F][25];	// lsu.scala:211:16
        stq_22_bits_uop_xcpt_pf_if = _RANDOM[10'h33F][26];	// lsu.scala:211:16
        stq_22_bits_uop_xcpt_ae_if = _RANDOM[10'h33F][27];	// lsu.scala:211:16
        stq_22_bits_uop_xcpt_ma_if = _RANDOM[10'h33F][28];	// lsu.scala:211:16
        stq_22_bits_uop_bp_debug_if = _RANDOM[10'h33F][29];	// lsu.scala:211:16
        stq_22_bits_uop_bp_xcpt_if = _RANDOM[10'h33F][30];	// lsu.scala:211:16
        stq_22_bits_uop_debug_fsrc = {_RANDOM[10'h33F][31], _RANDOM[10'h340][0]};	// lsu.scala:211:16
        stq_22_bits_uop_debug_tsrc = _RANDOM[10'h340][2:1];	// lsu.scala:211:16
        stq_22_bits_addr_valid = _RANDOM[10'h340][3];	// lsu.scala:211:16
        stq_22_bits_addr_bits = {_RANDOM[10'h340][31:4], _RANDOM[10'h341][11:0]};	// lsu.scala:211:16
        stq_22_bits_addr_is_virtual = _RANDOM[10'h341][12];	// lsu.scala:211:16
        stq_22_bits_data_valid = _RANDOM[10'h341][13];	// lsu.scala:211:16
        stq_22_bits_data_bits =
          {_RANDOM[10'h341][31:14], _RANDOM[10'h342], _RANDOM[10'h343][13:0]};	// lsu.scala:211:16
        stq_22_bits_committed = _RANDOM[10'h343][14];	// lsu.scala:211:16
        stq_22_bits_succeeded = _RANDOM[10'h343][15];	// lsu.scala:211:16
        stq_23_valid = _RANDOM[10'h345][16];	// lsu.scala:211:16
        stq_23_bits_uop_uopc = _RANDOM[10'h345][23:17];	// lsu.scala:211:16
        stq_23_bits_uop_inst = {_RANDOM[10'h345][31:24], _RANDOM[10'h346][23:0]};	// lsu.scala:211:16
        stq_23_bits_uop_debug_inst = {_RANDOM[10'h346][31:24], _RANDOM[10'h347][23:0]};	// lsu.scala:211:16
        stq_23_bits_uop_is_rvc = _RANDOM[10'h347][24];	// lsu.scala:211:16
        stq_23_bits_uop_debug_pc =
          {_RANDOM[10'h347][31:25], _RANDOM[10'h348], _RANDOM[10'h349][0]};	// lsu.scala:211:16
        stq_23_bits_uop_iq_type = _RANDOM[10'h349][3:1];	// lsu.scala:211:16
        stq_23_bits_uop_fu_code = _RANDOM[10'h349][13:4];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_br_type = _RANDOM[10'h349][17:14];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_op1_sel = _RANDOM[10'h349][19:18];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_op2_sel = _RANDOM[10'h349][22:20];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_imm_sel = _RANDOM[10'h349][25:23];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_op_fcn = _RANDOM[10'h349][29:26];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_fcn_dw = _RANDOM[10'h349][30];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h349][31], _RANDOM[10'h34A][1:0]};	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_is_load = _RANDOM[10'h34A][2];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_is_sta = _RANDOM[10'h34A][3];	// lsu.scala:211:16
        stq_23_bits_uop_ctrl_is_std = _RANDOM[10'h34A][4];	// lsu.scala:211:16
        stq_23_bits_uop_iw_state = _RANDOM[10'h34A][6:5];	// lsu.scala:211:16
        stq_23_bits_uop_iw_p1_poisoned = _RANDOM[10'h34A][7];	// lsu.scala:211:16
        stq_23_bits_uop_iw_p2_poisoned = _RANDOM[10'h34A][8];	// lsu.scala:211:16
        stq_23_bits_uop_is_br = _RANDOM[10'h34A][9];	// lsu.scala:211:16
        stq_23_bits_uop_is_jalr = _RANDOM[10'h34A][10];	// lsu.scala:211:16
        stq_23_bits_uop_is_jal = _RANDOM[10'h34A][11];	// lsu.scala:211:16
        stq_23_bits_uop_is_sfb = _RANDOM[10'h34A][12];	// lsu.scala:211:16
        stq_23_bits_uop_br_mask = _RANDOM[10'h34A][28:13];	// lsu.scala:211:16
        stq_23_bits_uop_br_tag = {_RANDOM[10'h34A][31:29], _RANDOM[10'h34B][0]};	// lsu.scala:211:16
        stq_23_bits_uop_ftq_idx = _RANDOM[10'h34B][5:1];	// lsu.scala:211:16
        stq_23_bits_uop_edge_inst = _RANDOM[10'h34B][6];	// lsu.scala:211:16
        stq_23_bits_uop_pc_lob = _RANDOM[10'h34B][12:7];	// lsu.scala:211:16
        stq_23_bits_uop_taken = _RANDOM[10'h34B][13];	// lsu.scala:211:16
        stq_23_bits_uop_imm_packed = {_RANDOM[10'h34B][31:14], _RANDOM[10'h34C][1:0]};	// lsu.scala:211:16
        stq_23_bits_uop_csr_addr = _RANDOM[10'h34C][13:2];	// lsu.scala:211:16
        stq_23_bits_uop_rob_idx = _RANDOM[10'h34C][20:14];	// lsu.scala:211:16
        stq_23_bits_uop_ldq_idx = _RANDOM[10'h34C][25:21];	// lsu.scala:211:16
        stq_23_bits_uop_stq_idx = _RANDOM[10'h34C][30:26];	// lsu.scala:211:16
        stq_23_bits_uop_rxq_idx = {_RANDOM[10'h34C][31], _RANDOM[10'h34D][0]};	// lsu.scala:211:16
        stq_23_bits_uop_pdst = _RANDOM[10'h34D][7:1];	// lsu.scala:211:16
        stq_23_bits_uop_prs1 = _RANDOM[10'h34D][14:8];	// lsu.scala:211:16
        stq_23_bits_uop_prs2 = _RANDOM[10'h34D][21:15];	// lsu.scala:211:16
        stq_23_bits_uop_prs3 = _RANDOM[10'h34D][28:22];	// lsu.scala:211:16
        stq_23_bits_uop_ppred = {_RANDOM[10'h34D][31:29], _RANDOM[10'h34E][1:0]};	// lsu.scala:211:16
        stq_23_bits_uop_prs1_busy = _RANDOM[10'h34E][2];	// lsu.scala:211:16
        stq_23_bits_uop_prs2_busy = _RANDOM[10'h34E][3];	// lsu.scala:211:16
        stq_23_bits_uop_prs3_busy = _RANDOM[10'h34E][4];	// lsu.scala:211:16
        stq_23_bits_uop_ppred_busy = _RANDOM[10'h34E][5];	// lsu.scala:211:16
        stq_23_bits_uop_stale_pdst = _RANDOM[10'h34E][12:6];	// lsu.scala:211:16
        stq_23_bits_uop_exception = _RANDOM[10'h34E][13];	// lsu.scala:211:16
        stq_23_bits_uop_exc_cause =
          {_RANDOM[10'h34E][31:14], _RANDOM[10'h34F], _RANDOM[10'h350][13:0]};	// lsu.scala:211:16
        stq_23_bits_uop_bypassable = _RANDOM[10'h350][14];	// lsu.scala:211:16
        stq_23_bits_uop_mem_cmd = _RANDOM[10'h350][19:15];	// lsu.scala:211:16
        stq_23_bits_uop_mem_size = _RANDOM[10'h350][21:20];	// lsu.scala:211:16
        stq_23_bits_uop_mem_signed = _RANDOM[10'h350][22];	// lsu.scala:211:16
        stq_23_bits_uop_is_fence = _RANDOM[10'h350][23];	// lsu.scala:211:16
        stq_23_bits_uop_is_fencei = _RANDOM[10'h350][24];	// lsu.scala:211:16
        stq_23_bits_uop_is_amo = _RANDOM[10'h350][25];	// lsu.scala:211:16
        stq_23_bits_uop_uses_ldq = _RANDOM[10'h350][26];	// lsu.scala:211:16
        stq_23_bits_uop_uses_stq = _RANDOM[10'h350][27];	// lsu.scala:211:16
        stq_23_bits_uop_is_sys_pc2epc = _RANDOM[10'h350][28];	// lsu.scala:211:16
        stq_23_bits_uop_is_unique = _RANDOM[10'h350][29];	// lsu.scala:211:16
        stq_23_bits_uop_flush_on_commit = _RANDOM[10'h350][30];	// lsu.scala:211:16
        stq_23_bits_uop_ldst_is_rs1 = _RANDOM[10'h350][31];	// lsu.scala:211:16
        stq_23_bits_uop_ldst = _RANDOM[10'h351][5:0];	// lsu.scala:211:16
        stq_23_bits_uop_lrs1 = _RANDOM[10'h351][11:6];	// lsu.scala:211:16
        stq_23_bits_uop_lrs2 = _RANDOM[10'h351][17:12];	// lsu.scala:211:16
        stq_23_bits_uop_lrs3 = _RANDOM[10'h351][23:18];	// lsu.scala:211:16
        stq_23_bits_uop_ldst_val = _RANDOM[10'h351][24];	// lsu.scala:211:16
        stq_23_bits_uop_dst_rtype = _RANDOM[10'h351][26:25];	// lsu.scala:211:16
        stq_23_bits_uop_lrs1_rtype = _RANDOM[10'h351][28:27];	// lsu.scala:211:16
        stq_23_bits_uop_lrs2_rtype = _RANDOM[10'h351][30:29];	// lsu.scala:211:16
        stq_23_bits_uop_frs3_en = _RANDOM[10'h351][31];	// lsu.scala:211:16
        stq_23_bits_uop_fp_val = _RANDOM[10'h352][0];	// lsu.scala:211:16
        stq_23_bits_uop_fp_single = _RANDOM[10'h352][1];	// lsu.scala:211:16
        stq_23_bits_uop_xcpt_pf_if = _RANDOM[10'h352][2];	// lsu.scala:211:16
        stq_23_bits_uop_xcpt_ae_if = _RANDOM[10'h352][3];	// lsu.scala:211:16
        stq_23_bits_uop_xcpt_ma_if = _RANDOM[10'h352][4];	// lsu.scala:211:16
        stq_23_bits_uop_bp_debug_if = _RANDOM[10'h352][5];	// lsu.scala:211:16
        stq_23_bits_uop_bp_xcpt_if = _RANDOM[10'h352][6];	// lsu.scala:211:16
        stq_23_bits_uop_debug_fsrc = _RANDOM[10'h352][8:7];	// lsu.scala:211:16
        stq_23_bits_uop_debug_tsrc = _RANDOM[10'h352][10:9];	// lsu.scala:211:16
        stq_23_bits_addr_valid = _RANDOM[10'h352][11];	// lsu.scala:211:16
        stq_23_bits_addr_bits = {_RANDOM[10'h352][31:12], _RANDOM[10'h353][19:0]};	// lsu.scala:211:16
        stq_23_bits_addr_is_virtual = _RANDOM[10'h353][20];	// lsu.scala:211:16
        stq_23_bits_data_valid = _RANDOM[10'h353][21];	// lsu.scala:211:16
        stq_23_bits_data_bits =
          {_RANDOM[10'h353][31:22], _RANDOM[10'h354], _RANDOM[10'h355][21:0]};	// lsu.scala:211:16
        stq_23_bits_committed = _RANDOM[10'h355][22];	// lsu.scala:211:16
        stq_23_bits_succeeded = _RANDOM[10'h355][23];	// lsu.scala:211:16
        ldq_head = _RANDOM[10'h357][28:24];	// lsu.scala:215:29
        ldq_tail = {_RANDOM[10'h357][31:29], _RANDOM[10'h358][1:0]};	// lsu.scala:215:29, :216:29
        stq_head = _RANDOM[10'h358][6:2];	// lsu.scala:216:29, :217:29
        stq_tail = _RANDOM[10'h358][11:7];	// lsu.scala:216:29, :218:29
        stq_commit_head = _RANDOM[10'h358][16:12];	// lsu.scala:216:29, :219:29
        stq_execute_head = _RANDOM[10'h358][21:17];	// lsu.scala:216:29, :220:29
        hella_state = _RANDOM[10'h358][24:22];	// lsu.scala:216:29, :242:38
        hella_req_addr = {_RANDOM[10'h358][31:25], _RANDOM[10'h359], _RANDOM[10'h35A][0]};	// lsu.scala:216:29, :243:34
        hella_req_cmd = _RANDOM[10'h35A][12:8];	// lsu.scala:243:34
        hella_req_size = _RANDOM[10'h35A][14:13];	// lsu.scala:243:34
        hella_req_signed = _RANDOM[10'h35A][15];	// lsu.scala:243:34
        hella_req_phys = _RANDOM[10'h35A][18];	// lsu.scala:243:34
        hella_data_data =
          {_RANDOM[10'h35C][31:29], _RANDOM[10'h35D], _RANDOM[10'h35E][28:0]};	// lsu.scala:244:34
        hella_paddr = {_RANDOM[10'h35F][31:5], _RANDOM[10'h360][4:0]};	// lsu.scala:245:34
        hella_xcpt_ma_ld = _RANDOM[10'h360][5];	// lsu.scala:245:34, :246:34
        hella_xcpt_ma_st = _RANDOM[10'h360][6];	// lsu.scala:245:34, :246:34
        hella_xcpt_pf_ld = _RANDOM[10'h360][7];	// lsu.scala:245:34, :246:34
        hella_xcpt_pf_st = _RANDOM[10'h360][8];	// lsu.scala:245:34, :246:34
        hella_xcpt_ae_ld = _RANDOM[10'h360][9];	// lsu.scala:245:34, :246:34
        hella_xcpt_ae_st = _RANDOM[10'h360][10];	// lsu.scala:245:34, :246:34
        live_store_mask = {_RANDOM[10'h360][31:11], _RANDOM[10'h361][2:0]};	// lsu.scala:245:34, :259:32
        p1_block_load_mask_0 = _RANDOM[10'h361][3];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_1 = _RANDOM[10'h361][4];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_2 = _RANDOM[10'h361][5];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_3 = _RANDOM[10'h361][6];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_4 = _RANDOM[10'h361][7];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_5 = _RANDOM[10'h361][8];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_6 = _RANDOM[10'h361][9];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_7 = _RANDOM[10'h361][10];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_8 = _RANDOM[10'h361][11];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_9 = _RANDOM[10'h361][12];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_10 = _RANDOM[10'h361][13];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_11 = _RANDOM[10'h361][14];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_12 = _RANDOM[10'h361][15];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_13 = _RANDOM[10'h361][16];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_14 = _RANDOM[10'h361][17];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_15 = _RANDOM[10'h361][18];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_16 = _RANDOM[10'h361][19];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_17 = _RANDOM[10'h361][20];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_18 = _RANDOM[10'h361][21];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_19 = _RANDOM[10'h361][22];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_20 = _RANDOM[10'h361][23];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_21 = _RANDOM[10'h361][24];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_22 = _RANDOM[10'h361][25];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_23 = _RANDOM[10'h361][26];	// lsu.scala:259:32, :398:35
        p2_block_load_mask_0 = _RANDOM[10'h361][27];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_1 = _RANDOM[10'h361][28];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_2 = _RANDOM[10'h361][29];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_3 = _RANDOM[10'h361][30];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_4 = _RANDOM[10'h361][31];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_5 = _RANDOM[10'h362][0];	// lsu.scala:399:35
        p2_block_load_mask_6 = _RANDOM[10'h362][1];	// lsu.scala:399:35
        p2_block_load_mask_7 = _RANDOM[10'h362][2];	// lsu.scala:399:35
        p2_block_load_mask_8 = _RANDOM[10'h362][3];	// lsu.scala:399:35
        p2_block_load_mask_9 = _RANDOM[10'h362][4];	// lsu.scala:399:35
        p2_block_load_mask_10 = _RANDOM[10'h362][5];	// lsu.scala:399:35
        p2_block_load_mask_11 = _RANDOM[10'h362][6];	// lsu.scala:399:35
        p2_block_load_mask_12 = _RANDOM[10'h362][7];	// lsu.scala:399:35
        p2_block_load_mask_13 = _RANDOM[10'h362][8];	// lsu.scala:399:35
        p2_block_load_mask_14 = _RANDOM[10'h362][9];	// lsu.scala:399:35
        p2_block_load_mask_15 = _RANDOM[10'h362][10];	// lsu.scala:399:35
        p2_block_load_mask_16 = _RANDOM[10'h362][11];	// lsu.scala:399:35
        p2_block_load_mask_17 = _RANDOM[10'h362][12];	// lsu.scala:399:35
        p2_block_load_mask_18 = _RANDOM[10'h362][13];	// lsu.scala:399:35
        p2_block_load_mask_19 = _RANDOM[10'h362][14];	// lsu.scala:399:35
        p2_block_load_mask_20 = _RANDOM[10'h362][15];	// lsu.scala:399:35
        p2_block_load_mask_21 = _RANDOM[10'h362][16];	// lsu.scala:399:35
        p2_block_load_mask_22 = _RANDOM[10'h362][17];	// lsu.scala:399:35
        p2_block_load_mask_23 = _RANDOM[10'h362][18];	// lsu.scala:399:35
        ldq_retry_idx = _RANDOM[10'h362][24:20];	// lsu.scala:399:35, :415:30
        stq_retry_idx = _RANDOM[10'h362][29:25];	// lsu.scala:399:35, :422:30
        ldq_wakeup_idx = {_RANDOM[10'h362][31:30], _RANDOM[10'h363][2:0]};	// lsu.scala:399:35, :430:31
        can_fire_load_retry_REG = _RANDOM[10'h363][3];	// lsu.scala:430:31, :470:40
        can_fire_sta_retry_REG = _RANDOM[10'h363][4];	// lsu.scala:430:31, :482:41
        mem_xcpt_valids_0 = _RANDOM[10'h363][5];	// lsu.scala:430:31, :667:32
        mem_xcpt_uops_0_br_mask = _RANDOM[10'h368][17:2];	// lsu.scala:671:32
        mem_xcpt_uops_0_rob_idx = _RANDOM[10'h36A][9:3];	// lsu.scala:671:32
        mem_xcpt_uops_0_ldq_idx = _RANDOM[10'h36A][14:10];	// lsu.scala:671:32
        mem_xcpt_uops_0_stq_idx = _RANDOM[10'h36A][19:15];	// lsu.scala:671:32
        mem_xcpt_uops_0_uses_ldq = _RANDOM[10'h36E][15];	// lsu.scala:671:32
        mem_xcpt_uops_0_uses_stq = _RANDOM[10'h36E][16];	// lsu.scala:671:32
        mem_xcpt_causes_0 = _RANDOM[10'h370][3:0];	// lsu.scala:672:32
        mem_xcpt_vaddrs_0 = {_RANDOM[10'h370][31:4], _RANDOM[10'h371][11:0]};	// lsu.scala:672:32, :679:32
        REG = _RANDOM[10'h371][12];	// lsu.scala:679:32, :718:21
        fired_load_incoming_REG = _RANDOM[10'h371][13];	// lsu.scala:679:32, :894:51
        fired_stad_incoming_REG = _RANDOM[10'h371][14];	// lsu.scala:679:32, :895:51
        fired_sta_incoming_REG = _RANDOM[10'h371][15];	// lsu.scala:679:32, :896:51
        fired_std_incoming_REG = _RANDOM[10'h371][16];	// lsu.scala:679:32, :897:51
        fired_stdf_incoming = _RANDOM[10'h371][17];	// lsu.scala:679:32, :898:37
        fired_sfence_0 = _RANDOM[10'h371][18];	// lsu.scala:679:32, :899:37
        fired_release_0 = _RANDOM[10'h371][19];	// lsu.scala:679:32, :900:37
        fired_load_retry_REG = _RANDOM[10'h371][20];	// lsu.scala:679:32, :901:51
        fired_sta_retry_REG = _RANDOM[10'h371][21];	// lsu.scala:679:32, :902:51
        fired_load_wakeup_REG = _RANDOM[10'h371][23];	// lsu.scala:679:32, :904:51
        mem_incoming_uop_0_br_mask = {_RANDOM[10'h376][31:22], _RANDOM[10'h377][5:0]};	// lsu.scala:908:37
        mem_incoming_uop_0_rob_idx = _RANDOM[10'h378][29:23];	// lsu.scala:908:37
        mem_incoming_uop_0_ldq_idx = {_RANDOM[10'h378][31:30], _RANDOM[10'h379][2:0]};	// lsu.scala:908:37
        mem_incoming_uop_0_stq_idx = _RANDOM[10'h379][7:3];	// lsu.scala:908:37
        mem_incoming_uop_0_pdst = _RANDOM[10'h379][16:10];	// lsu.scala:908:37
        mem_incoming_uop_0_fp_val = _RANDOM[10'h37E][9];	// lsu.scala:908:37
        mem_ldq_incoming_e_0_bits_uop_br_mask =
          {_RANDOM[10'h383][31:17], _RANDOM[10'h384][0]};	// lsu.scala:909:37
        mem_ldq_incoming_e_0_bits_uop_stq_idx =
          {_RANDOM[10'h385][31:30], _RANDOM[10'h386][2:0]};	// lsu.scala:909:37
        mem_ldq_incoming_e_0_bits_uop_mem_size = _RANDOM[10'h389][25:24];	// lsu.scala:909:37
        mem_ldq_incoming_e_0_bits_st_dep_mask =
          {_RANDOM[10'h38C][31:30], _RANDOM[10'h38D][21:0]};	// lsu.scala:909:37
        mem_stq_incoming_e_0_valid = _RANDOM[10'h390][1];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_br_mask =
          {_RANDOM[10'h394][31:30], _RANDOM[10'h395][13:0]};	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_rob_idx =
          {_RANDOM[10'h396][31], _RANDOM[10'h397][5:0]};	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_stq_idx = _RANDOM[10'h397][15:11];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_mem_size = _RANDOM[10'h39B][6:5];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_is_amo = _RANDOM[10'h39B][10];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_addr_valid = _RANDOM[10'h39C][28];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_addr_is_virtual = _RANDOM[10'h39E][5];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_data_valid = _RANDOM[10'h39E][6];	// lsu.scala:910:37
        mem_ldq_wakeup_e_bits_uop_br_mask = _RANDOM[10'h3A7][21:6];	// lsu.scala:911:37
        mem_ldq_wakeup_e_bits_uop_stq_idx = _RANDOM[10'h3A9][23:19];	// lsu.scala:911:37
        mem_ldq_wakeup_e_bits_uop_mem_size = _RANDOM[10'h3AD][14:13];	// lsu.scala:911:37
        mem_ldq_wakeup_e_bits_st_dep_mask =
          {_RANDOM[10'h3B0][31:19], _RANDOM[10'h3B1][10:0]};	// lsu.scala:911:37
        mem_ldq_retry_e_bits_uop_br_mask =
          {_RANDOM[10'h3B8][31:19], _RANDOM[10'h3B9][2:0]};	// lsu.scala:912:37
        mem_ldq_retry_e_bits_uop_stq_idx = _RANDOM[10'h3BB][4:0];	// lsu.scala:912:37
        mem_ldq_retry_e_bits_uop_mem_size = _RANDOM[10'h3BE][27:26];	// lsu.scala:912:37
        mem_ldq_retry_e_bits_st_dep_mask = _RANDOM[10'h3C2][23:0];	// lsu.scala:912:37
        mem_stq_retry_e_valid = _RANDOM[10'h3C5][3];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_br_mask = _RANDOM[10'h3CA][15:0];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_rob_idx = _RANDOM[10'h3CC][7:1];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_stq_idx = _RANDOM[10'h3CC][17:13];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_mem_size = _RANDOM[10'h3D0][8:7];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_is_amo = _RANDOM[10'h3D0][12];	// lsu.scala:913:37
        mem_stq_retry_e_bits_data_valid = _RANDOM[10'h3D3][8];	// lsu.scala:913:37
        mem_stdf_uop_br_mask = _RANDOM[10'h3DC][22:7];	// lsu.scala:922:37
        mem_stdf_uop_rob_idx = _RANDOM[10'h3DE][14:8];	// lsu.scala:922:37
        mem_stdf_uop_stq_idx = _RANDOM[10'h3DE][24:20];	// lsu.scala:922:37
        mem_tlb_miss_0 = _RANDOM[10'h3E4][5];	// lsu.scala:925:41
        mem_tlb_uncacheable_0 = _RANDOM[10'h3E4][6];	// lsu.scala:925:41, :926:41
        mem_paddr_0 = {_RANDOM[10'h3E4][31:7], _RANDOM[10'h3E5][14:0]};	// lsu.scala:925:41, :927:41
        clr_bsy_valid_0 = _RANDOM[10'h3E5][15];	// lsu.scala:927:41, :930:32
        clr_bsy_rob_idx_0 = _RANDOM[10'h3E5][22:16];	// lsu.scala:927:41, :931:28
        clr_bsy_brmask_0 = {_RANDOM[10'h3E5][31:23], _RANDOM[10'h3E6][6:0]};	// lsu.scala:927:41, :932:28
        io_core_clr_bsy_0_valid_REG = _RANDOM[10'h3E6][7];	// lsu.scala:932:28, :979:62
        io_core_clr_bsy_0_valid_REG_1 = _RANDOM[10'h3E6][8];	// lsu.scala:932:28, :979:101
        io_core_clr_bsy_0_valid_REG_2 = _RANDOM[10'h3E6][9];	// lsu.scala:932:28, :979:93
        stdf_clr_bsy_valid = _RANDOM[10'h3E6][10];	// lsu.scala:932:28, :983:37
        stdf_clr_bsy_rob_idx = _RANDOM[10'h3E6][17:11];	// lsu.scala:932:28, :984:33
        stdf_clr_bsy_brmask = {_RANDOM[10'h3E6][31:18], _RANDOM[10'h3E7][1:0]};	// lsu.scala:932:28, :985:33
        io_core_clr_bsy_1_valid_REG = _RANDOM[10'h3E7][2];	// lsu.scala:985:33, :1004:67
        io_core_clr_bsy_1_valid_REG_1 = _RANDOM[10'h3E7][3];	// lsu.scala:985:33, :1004:106
        io_core_clr_bsy_1_valid_REG_2 = _RANDOM[10'h3E7][4];	// lsu.scala:985:33, :1004:98
        lcam_addr_REG = {_RANDOM[10'h3E7][31:5], _RANDOM[10'h3E8][4:0]};	// lsu.scala:985:33, :1026:45
        lcam_addr_REG_1 = {_RANDOM[10'h3E8][31:5], _RANDOM[10'h3E9][4:0]};	// lsu.scala:1026:45, :1027:67
        lcam_ldq_idx_REG = _RANDOM[10'h3E9][9:5];	// lsu.scala:1027:67, :1037:58
        lcam_ldq_idx_REG_1 = _RANDOM[10'h3E9][14:10];	// lsu.scala:1027:67, :1038:58
        lcam_stq_idx_REG = _RANDOM[10'h3E9][19:15];	// lsu.scala:1027:67, :1042:58
        s1_executing_loads_0 = _RANDOM[10'h3E9][20];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_1 = _RANDOM[10'h3E9][21];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_2 = _RANDOM[10'h3E9][22];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_3 = _RANDOM[10'h3E9][23];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_4 = _RANDOM[10'h3E9][24];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_5 = _RANDOM[10'h3E9][25];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_6 = _RANDOM[10'h3E9][26];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_7 = _RANDOM[10'h3E9][27];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_8 = _RANDOM[10'h3E9][28];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_9 = _RANDOM[10'h3E9][29];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_10 = _RANDOM[10'h3E9][30];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_11 = _RANDOM[10'h3E9][31];	// lsu.scala:1027:67, :1056:35
        s1_executing_loads_12 = _RANDOM[10'h3EA][0];	// lsu.scala:1056:35
        s1_executing_loads_13 = _RANDOM[10'h3EA][1];	// lsu.scala:1056:35
        s1_executing_loads_14 = _RANDOM[10'h3EA][2];	// lsu.scala:1056:35
        s1_executing_loads_15 = _RANDOM[10'h3EA][3];	// lsu.scala:1056:35
        s1_executing_loads_16 = _RANDOM[10'h3EA][4];	// lsu.scala:1056:35
        s1_executing_loads_17 = _RANDOM[10'h3EA][5];	// lsu.scala:1056:35
        s1_executing_loads_18 = _RANDOM[10'h3EA][6];	// lsu.scala:1056:35
        s1_executing_loads_19 = _RANDOM[10'h3EA][7];	// lsu.scala:1056:35
        s1_executing_loads_20 = _RANDOM[10'h3EA][8];	// lsu.scala:1056:35
        s1_executing_loads_21 = _RANDOM[10'h3EA][9];	// lsu.scala:1056:35
        s1_executing_loads_22 = _RANDOM[10'h3EA][10];	// lsu.scala:1056:35
        s1_executing_loads_23 = _RANDOM[10'h3EA][11];	// lsu.scala:1056:35
        wb_forward_valid_0 = _RANDOM[10'h3EA][12];	// lsu.scala:1056:35, :1064:36
        wb_forward_ldq_idx_0 = _RANDOM[10'h3EA][17:13];	// lsu.scala:1056:35, :1065:36
        wb_forward_ld_addr_0 = {_RANDOM[10'h3EA][31:18], _RANDOM[10'h3EB][25:0]};	// lsu.scala:1056:35, :1066:36
        wb_forward_stq_idx_0 = _RANDOM[10'h3EB][30:26];	// lsu.scala:1066:36, :1067:36
        older_nacked_REG = _RANDOM[10'h3EB][31];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG = _RANDOM[10'h3EC][0];	// lsu.scala:1131:58
        older_nacked_REG_1 = _RANDOM[10'h3EC][1];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_1 = _RANDOM[10'h3EC][2];	// lsu.scala:1131:58
        older_nacked_REG_2 = _RANDOM[10'h3EC][3];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_2 = _RANDOM[10'h3EC][4];	// lsu.scala:1131:58
        older_nacked_REG_3 = _RANDOM[10'h3EC][5];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_3 = _RANDOM[10'h3EC][6];	// lsu.scala:1131:58
        older_nacked_REG_4 = _RANDOM[10'h3EC][7];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_4 = _RANDOM[10'h3EC][8];	// lsu.scala:1131:58
        older_nacked_REG_5 = _RANDOM[10'h3EC][9];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_5 = _RANDOM[10'h3EC][10];	// lsu.scala:1131:58
        older_nacked_REG_6 = _RANDOM[10'h3EC][11];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_6 = _RANDOM[10'h3EC][12];	// lsu.scala:1131:58
        older_nacked_REG_7 = _RANDOM[10'h3EC][13];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_7 = _RANDOM[10'h3EC][14];	// lsu.scala:1131:58
        older_nacked_REG_8 = _RANDOM[10'h3EC][15];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_8 = _RANDOM[10'h3EC][16];	// lsu.scala:1131:58
        older_nacked_REG_9 = _RANDOM[10'h3EC][17];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_9 = _RANDOM[10'h3EC][18];	// lsu.scala:1131:58
        older_nacked_REG_10 = _RANDOM[10'h3EC][19];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_10 = _RANDOM[10'h3EC][20];	// lsu.scala:1131:58
        older_nacked_REG_11 = _RANDOM[10'h3EC][21];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_11 = _RANDOM[10'h3EC][22];	// lsu.scala:1131:58
        older_nacked_REG_12 = _RANDOM[10'h3EC][23];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_12 = _RANDOM[10'h3EC][24];	// lsu.scala:1131:58
        older_nacked_REG_13 = _RANDOM[10'h3EC][25];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_13 = _RANDOM[10'h3EC][26];	// lsu.scala:1131:58
        older_nacked_REG_14 = _RANDOM[10'h3EC][27];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_14 = _RANDOM[10'h3EC][28];	// lsu.scala:1131:58
        older_nacked_REG_15 = _RANDOM[10'h3EC][29];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_15 = _RANDOM[10'h3EC][30];	// lsu.scala:1131:58
        older_nacked_REG_16 = _RANDOM[10'h3EC][31];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_16 = _RANDOM[10'h3ED][0];	// lsu.scala:1131:58
        older_nacked_REG_17 = _RANDOM[10'h3ED][1];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_17 = _RANDOM[10'h3ED][2];	// lsu.scala:1131:58
        older_nacked_REG_18 = _RANDOM[10'h3ED][3];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_18 = _RANDOM[10'h3ED][4];	// lsu.scala:1131:58
        older_nacked_REG_19 = _RANDOM[10'h3ED][5];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_19 = _RANDOM[10'h3ED][6];	// lsu.scala:1131:58
        older_nacked_REG_20 = _RANDOM[10'h3ED][7];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_20 = _RANDOM[10'h3ED][8];	// lsu.scala:1131:58
        older_nacked_REG_21 = _RANDOM[10'h3ED][9];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_21 = _RANDOM[10'h3ED][10];	// lsu.scala:1131:58
        older_nacked_REG_22 = _RANDOM[10'h3ED][11];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_22 = _RANDOM[10'h3ED][12];	// lsu.scala:1131:58
        older_nacked_REG_23 = _RANDOM[10'h3ED][13];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_23 = _RANDOM[10'h3ED][14];	// lsu.scala:1131:58
        io_dmem_s1_kill_0_REG_24 = _RANDOM[10'h3ED][15];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_25 = _RANDOM[10'h3ED][16];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_26 = _RANDOM[10'h3ED][17];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_27 = _RANDOM[10'h3ED][18];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_28 = _RANDOM[10'h3ED][19];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_29 = _RANDOM[10'h3ED][20];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_30 = _RANDOM[10'h3ED][21];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_31 = _RANDOM[10'h3ED][22];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_32 = _RANDOM[10'h3ED][23];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_33 = _RANDOM[10'h3ED][24];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_34 = _RANDOM[10'h3ED][25];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_35 = _RANDOM[10'h3ED][26];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_36 = _RANDOM[10'h3ED][27];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_37 = _RANDOM[10'h3ED][28];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_38 = _RANDOM[10'h3ED][29];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_39 = _RANDOM[10'h3ED][30];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_40 = _RANDOM[10'h3ED][31];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_41 = _RANDOM[10'h3EE][0];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_42 = _RANDOM[10'h3EE][1];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_43 = _RANDOM[10'h3EE][2];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_44 = _RANDOM[10'h3EE][3];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_45 = _RANDOM[10'h3EE][4];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_46 = _RANDOM[10'h3EE][5];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_47 = _RANDOM[10'h3EE][6];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_48 = _RANDOM[10'h3EE][7];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_49 = _RANDOM[10'h3EE][8];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_50 = _RANDOM[10'h3EE][9];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_51 = _RANDOM[10'h3EE][10];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_52 = _RANDOM[10'h3EE][11];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_53 = _RANDOM[10'h3EE][12];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_54 = _RANDOM[10'h3EE][13];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_55 = _RANDOM[10'h3EE][14];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_56 = _RANDOM[10'h3EE][15];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_57 = _RANDOM[10'h3EE][16];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_58 = _RANDOM[10'h3EE][17];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_59 = _RANDOM[10'h3EE][18];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_60 = _RANDOM[10'h3EE][19];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_61 = _RANDOM[10'h3EE][20];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_62 = _RANDOM[10'h3EE][21];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_63 = _RANDOM[10'h3EE][22];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_64 = _RANDOM[10'h3EE][23];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_65 = _RANDOM[10'h3EE][24];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_66 = _RANDOM[10'h3EE][25];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_67 = _RANDOM[10'h3EE][26];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_68 = _RANDOM[10'h3EE][27];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_69 = _RANDOM[10'h3EE][28];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_70 = _RANDOM[10'h3EE][29];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_71 = _RANDOM[10'h3EE][30];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_72 = _RANDOM[10'h3EE][31];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_73 = _RANDOM[10'h3EF][0];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_74 = _RANDOM[10'h3EF][1];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_75 = _RANDOM[10'h3EF][2];	// lsu.scala:1153:56, :1159:56
        io_dmem_s1_kill_0_REG_76 = _RANDOM[10'h3EF][3];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_77 = _RANDOM[10'h3EF][4];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_78 = _RANDOM[10'h3EF][5];	// lsu.scala:1153:56, :1159:56
        io_dmem_s1_kill_0_REG_79 = _RANDOM[10'h3EF][6];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_80 = _RANDOM[10'h3EF][7];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_81 = _RANDOM[10'h3EF][8];	// lsu.scala:1153:56, :1159:56
        io_dmem_s1_kill_0_REG_82 = _RANDOM[10'h3EF][9];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_83 = _RANDOM[10'h3EF][10];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_84 = _RANDOM[10'h3EF][11];	// lsu.scala:1153:56, :1159:56
        io_dmem_s1_kill_0_REG_85 = _RANDOM[10'h3EF][12];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_86 = _RANDOM[10'h3EF][13];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_87 = _RANDOM[10'h3EF][14];	// lsu.scala:1153:56, :1159:56
        io_dmem_s1_kill_0_REG_88 = _RANDOM[10'h3EF][15];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_89 = _RANDOM[10'h3EF][16];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_90 = _RANDOM[10'h3EF][17];	// lsu.scala:1153:56, :1159:56
        io_dmem_s1_kill_0_REG_91 = _RANDOM[10'h3EF][18];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_92 = _RANDOM[10'h3EF][19];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_93 = _RANDOM[10'h3EF][20];	// lsu.scala:1153:56, :1159:56
        io_dmem_s1_kill_0_REG_94 = _RANDOM[10'h3EF][21];	// lsu.scala:1159:56
        io_dmem_s1_kill_0_REG_95 = _RANDOM[10'h3EF][22];	// lsu.scala:1159:56, :1165:56
        REG_1 = _RANDOM[10'h3EF][23];	// lsu.scala:1159:56, :1189:64
        REG_2 = _RANDOM[10'h3EF][24];	// lsu.scala:1159:56, :1199:18
        store_blocked_counter = _RANDOM[10'h3EF][28:25];	// lsu.scala:1159:56, :1204:36
        r_xcpt_valid = _RANDOM[10'h3F0][5];	// lsu.scala:1235:29
        r_xcpt_uop_br_mask = _RANDOM[10'h3F5][17:2];	// lsu.scala:1236:25
        r_xcpt_uop_rob_idx = _RANDOM[10'h3F7][9:3];	// lsu.scala:1236:25
        r_xcpt_cause = _RANDOM[10'h3FD][4:0];	// lsu.scala:1236:25
        r_xcpt_badvaddr = {_RANDOM[10'h3FD][31:5], _RANDOM[10'h3FE][12:0]};	// lsu.scala:1236:25
        io_core_ld_miss_REG = _RANDOM[10'h3FE][13];	// lsu.scala:1236:25, :1380:37
        spec_ld_succeed_REG = _RANDOM[10'h3FE][14];	// lsu.scala:1236:25, :1382:13
        spec_ld_succeed_REG_1 = _RANDOM[10'h3FE][19:15];	// lsu.scala:1236:25, :1384:56
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  NBDTLB_1 dtlb (	// lsu.scala:249:20
    .clock                        (clock),
    .reset                        (reset),
    .io_req_0_valid               (~_will_fire_store_commit_0_T_2),	// lsu.scala:538:31, :576:25
    .io_req_0_bits_vaddr          (exe_tlb_vaddr_0),	// lsu.scala:607:24
    .io_req_0_bits_passthrough    (will_fire_hella_incoming_0 & hella_req_phys),	// lsu.scala:243:34, :535:65, :643:23
    .io_req_0_bits_size
      (_exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0 | will_fire_load_retry_0
       | will_fire_sta_retry_0
         ? exe_tlb_uop_0_mem_size
         : will_fire_hella_incoming_0 ? hella_req_size : 2'h0),	// lsu.scala:243:34, :535:65, :536:61, :567:63, :597:24, :624:23, :628:52, :630:23
    .io_req_0_bits_cmd
      (_exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0 | will_fire_load_retry_0
       | will_fire_sta_retry_0
         ? exe_tlb_uop_0_mem_cmd
         : will_fire_hella_incoming_0 ? hella_req_cmd : 5'h0),	// lsu.scala:243:34, :535:65, :536:61, :567:63, :597:24, :633:23, :637:52, :639:23
    .io_sfence_valid
      (will_fire_sfence_0 & io_core_exe_0_req_bits_sfence_valid),	// lsu.scala:536:61, :618:32, :619:18
    .io_sfence_bits_rs1
      (will_fire_sfence_0 & io_core_exe_0_req_bits_sfence_bits_rs1),	// lsu.scala:536:61, :618:32, :619:18
    .io_sfence_bits_rs2
      (will_fire_sfence_0 & io_core_exe_0_req_bits_sfence_bits_rs2),	// lsu.scala:536:61, :618:32, :619:18
    .io_sfence_bits_addr
      (will_fire_sfence_0 ? io_core_exe_0_req_bits_sfence_bits_addr : 39'h0),	// lsu.scala:536:61, :616:43, :618:32, :619:18
    .io_ptw_req_ready             (io_ptw_req_ready),
    .io_ptw_resp_valid            (io_ptw_resp_valid),
    .io_ptw_resp_bits_ae          (io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn     (io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d       (io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a       (io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g       (io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u       (io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x       (io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w       (io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r       (io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v       (io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level       (io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous (io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode             (io_ptw_ptbr_mode),
    .io_ptw_status_dprv           (io_ptw_status_dprv),
    .io_ptw_status_mxr            (io_ptw_status_mxr),
    .io_ptw_status_sum            (io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l           (io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a           (io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x           (io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w           (io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r           (io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr            (io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask            (io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l           (io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a           (io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x           (io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w           (io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r           (io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr            (io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask            (io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l           (io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a           (io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x           (io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w           (io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r           (io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr            (io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask            (io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l           (io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a           (io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x           (io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w           (io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r           (io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr            (io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask            (io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l           (io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a           (io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x           (io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w           (io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r           (io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr            (io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask            (io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l           (io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a           (io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x           (io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w           (io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r           (io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr            (io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask            (io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l           (io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a           (io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x           (io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w           (io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r           (io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr            (io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask            (io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l           (io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a           (io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x           (io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w           (io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r           (io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr            (io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask            (io_ptw_pmp_7_mask),
    .io_kill                      (will_fire_hella_incoming_0 & io_hellacache_s1_kill),	// lsu.scala:535:65, :646:23
    .io_miss_rdy                  (_dtlb_io_miss_rdy),
    .io_resp_0_miss               (_dtlb_io_resp_0_miss),
    .io_resp_0_paddr              (_dtlb_io_resp_0_paddr),
    .io_resp_0_pf_ld              (_dtlb_io_resp_0_pf_ld),
    .io_resp_0_pf_st              (_dtlb_io_resp_0_pf_st),
    .io_resp_0_ae_ld              (_dtlb_io_resp_0_ae_ld),
    .io_resp_0_ae_st              (_dtlb_io_resp_0_ae_st),
    .io_resp_0_ma_ld              (_dtlb_io_resp_0_ma_ld),
    .io_resp_0_ma_st              (_dtlb_io_resp_0_ma_st),
    .io_resp_0_cacheable          (_dtlb_io_resp_0_cacheable),
    .io_ptw_req_valid             (io_ptw_req_valid),
    .io_ptw_req_bits_valid        (io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr    (io_ptw_req_bits_bits_addr)
  );
  ForwardingAgeLogic_2 forwarding_age_logic_0 (	// lsu.scala:1178:57
    .io_addr_matches
      ({ldst_addr_matches_0_23,
        ldst_addr_matches_0_22,
        ldst_addr_matches_0_21,
        ldst_addr_matches_0_20,
        ldst_addr_matches_0_19,
        ldst_addr_matches_0_18,
        ldst_addr_matches_0_17,
        ldst_addr_matches_0_16,
        ldst_addr_matches_0_15,
        ldst_addr_matches_0_14,
        ldst_addr_matches_0_13,
        ldst_addr_matches_0_12,
        ldst_addr_matches_0_11,
        ldst_addr_matches_0_10,
        ldst_addr_matches_0_9,
        ldst_addr_matches_0_8,
        ldst_addr_matches_0_7,
        ldst_addr_matches_0_6,
        ldst_addr_matches_0_5,
        ldst_addr_matches_0_4,
        ldst_addr_matches_0_3,
        ldst_addr_matches_0_2,
        ldst_addr_matches_0_1,
        ldst_addr_matches_0_0}),	// lsu.scala:1148:72, :1150:9, :1180:72
    .io_youngest_st_idx
      (do_st_search_0
         ? (_lcam_stq_idx_T
              ? mem_stq_incoming_e_0_bits_uop_stq_idx
              : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_stq_idx : 5'h0)
         : do_ld_search_0
             ? (fired_load_incoming_REG
                  ? mem_ldq_incoming_e_0_bits_uop_stq_idx
                  : fired_load_retry_REG
                      ? mem_ldq_retry_e_bits_uop_stq_idx
                      : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_uop_stq_idx : 5'h0)
             : 5'h0),	// lsu.scala:894:51, :901:51, :902:51, :904:51, :909:37, :910:37, :911:37, :912:37, :913:37, :915:33, :916:33, :917:33, :919:{33,57}, :921:33, :1014:108, :1016:106, :1029:37, :1030:37
    .io_forwarding_idx  (_forwarding_age_logic_0_io_forwarding_idx)
  );
  assign io_core_exe_0_iresp_valid = _io_core_exe_0_iresp_valid_output;	// lsu.scala:1306:5, :1344:5, :1348:5
  assign io_core_exe_0_iresp_bits_uop_rob_idx =
    _GEN_801
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_148[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_36[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_790;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_pdst =
    _GEN_801
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_153[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_40[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_791;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_is_amo =
    _GEN_801
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_171[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_61[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_794;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_uses_stq =
    _GEN_801
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_174[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_64[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_795;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_dst_rtype =
    _GEN_801
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_185[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_74[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_796;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_data =
    _GEN_801
      ? io_dmem_resp_0_bits_data
      : {_ldq_bits_debug_wb_data_T_17
           ? {56{_GEN_793 & io_core_exe_0_iresp_bits_data_lo_2[7]}}
           : {_ldq_bits_debug_wb_data_T_9
                ? {48{_GEN_793 & io_core_exe_0_iresp_bits_data_lo_1[15]}}
                : {_ldq_bits_debug_wb_data_T_1
                     ? {32{_GEN_793 & io_core_exe_0_iresp_bits_data_lo[31]}}
                     : _GEN_800[63:32],
                   io_core_exe_0_iresp_bits_data_lo[31:16]},
              io_core_exe_0_iresp_bits_data_lo_1[15:8]},
         io_core_exe_0_iresp_bits_data_lo_2};	// AMOALU.scala:26:13, :39:{24,37}, :42:{20,26,76,85,98}, Bitwise.scala:72:12, Cat.scala:30:58, lsu.scala:1306:5, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_valid = _io_core_exe_0_fresp_valid_output;	// lsu.scala:1306:5, :1344:5, :1348:5
  assign io_core_exe_0_fresp_bits_uop_uopc =
    _GEN_801 ? _GEN_116[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_116[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_br_mask =
    _GEN_801 ? _GEN_110[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_789;	// lsu.scala:264:49, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_rob_idx =
    _GEN_801 ? _GEN_148[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_790;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_stq_idx =
    _GEN_801 ? _GEN_111[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_111[wb_forward_ldq_idx_0];	// lsu.scala:264:49, :1065:36, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_pdst =
    _GEN_801 ? _GEN_153[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_791;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_mem_size =
    _GEN_801 ? _GEN_112[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_792;	// lsu.scala:264:49, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_is_amo =
    _GEN_801 ? _GEN_171[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_794;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_uses_stq =
    _GEN_801 ? _GEN_174[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_795;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_dst_rtype =
    _GEN_801 ? _GEN_185[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_796;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_fp_val =
    _GEN_801 ? _GEN_189[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_189[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_data =
    {1'h0,
     _GEN_801
       ? io_dmem_resp_0_bits_data
       : {_ldq_bits_debug_wb_data_T_17
            ? {56{_GEN_793 & io_core_exe_0_fresp_bits_data_lo_2[7]}}
            : {_ldq_bits_debug_wb_data_T_9
                 ? {48{_GEN_793 & io_core_exe_0_fresp_bits_data_lo_1[15]}}
                 : {_ldq_bits_debug_wb_data_T_1
                      ? {32{_GEN_793 & io_core_exe_0_fresp_bits_data_lo[31]}}
                      : _GEN_800[63:32],
                    io_core_exe_0_fresp_bits_data_lo[31:16]},
               io_core_exe_0_fresp_bits_data_lo_1[15:8]},
          io_core_exe_0_fresp_bits_data_lo_2}};	// AMOALU.scala:26:13, :39:{24,37}, :42:{20,26,76,85,98}, Bitwise.scala:72:12, lsu.scala:249:20, :708:86, :1306:5, :1344:5, :1348:5, :1367:38, util.scala:118:51
  assign io_core_dis_ldq_idx_0 = ldq_tail;	// lsu.scala:216:29
  assign io_core_dis_ldq_idx_1 = _GEN_100;	// lsu.scala:333:21
  assign io_core_dis_ldq_idx_2 = _GEN_106;	// lsu.scala:333:21
  assign io_core_dis_stq_idx_0 = stq_tail;	// lsu.scala:218:29
  assign io_core_dis_stq_idx_1 = _GEN_101;	// lsu.scala:338:21
  assign io_core_dis_stq_idx_2 = _GEN_107;	// lsu.scala:338:21
  assign io_core_ldq_full_0 = _GEN_96 == ldq_head;	// lsu.scala:215:29, :293:51, util.scala:206:10
  assign io_core_ldq_full_1 = _GEN_103 == ldq_head;	// lsu.scala:215:29, :293:51, util.scala:206:10
  assign io_core_ldq_full_2 = (wrap_8 ? 5'h0 : _GEN_108) == ldq_head;	// lsu.scala:215:29, :293:51, util.scala:205:25, :206:{10,28}
  assign io_core_stq_full_0 = _GEN_98 == stq_head;	// lsu.scala:217:29, :297:51, util.scala:206:10
  assign io_core_stq_full_1 = _GEN_105 == stq_head;	// lsu.scala:217:29, :297:51, util.scala:206:10
  assign io_core_stq_full_2 = (wrap_9 ? 5'h0 : _GEN_109) == stq_head;	// lsu.scala:217:29, :297:51, util.scala:205:25, :206:{10,28}
  assign io_core_fp_stdata_ready = _io_core_fp_stdata_ready_output;	// lsu.scala:866:61
  assign io_core_clr_bsy_0_valid =
    clr_bsy_valid_0 & (io_core_brupdate_b1_mispredict_mask & clr_bsy_brmask_0) == 16'h0
    & ~io_core_exception & ~io_core_clr_bsy_0_valid_REG & ~io_core_clr_bsy_0_valid_REG_2;	// lsu.scala:669:22, :930:32, :932:28, :979:{54,62,82,85,93}, util.scala:118:{51,59}
  assign io_core_clr_bsy_0_bits = clr_bsy_rob_idx_0;	// lsu.scala:931:28
  assign io_core_clr_bsy_1_valid =
    stdf_clr_bsy_valid
    & (io_core_brupdate_b1_mispredict_mask & stdf_clr_bsy_brmask) == 16'h0
    & ~io_core_exception & ~io_core_clr_bsy_1_valid_REG & ~io_core_clr_bsy_1_valid_REG_2;	// lsu.scala:669:22, :983:37, :985:33, :1004:{59,67,87,90,98}, util.scala:118:{51,59}
  assign io_core_clr_bsy_1_bits = stdf_clr_bsy_rob_idx;	// lsu.scala:984:33
  assign io_core_spec_ld_wakeup_0_valid = _io_core_spec_ld_wakeup_0_valid_output;	// lsu.scala:1260:69
  assign io_core_spec_ld_wakeup_0_bits = mem_incoming_uop_0_pdst;	// lsu.scala:908:37
  assign io_core_ld_miss =
    ~(~spec_ld_succeed_REG | _io_core_exe_0_iresp_valid_output
      & (_GEN_801
           ? (io_dmem_resp_0_bits_uop_uses_ldq
                ? _GEN_150[io_dmem_resp_0_bits_uop_ldq_idx]
                : _GEN_37[io_dmem_resp_0_bits_uop_stq_idx])
           : _GEN_150[wb_forward_ldq_idx_0]) == spec_ld_succeed_REG_1)
    & io_core_ld_miss_REG;	// lsu.scala:224:42, :465:79, :1065:36, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, :1380:{27,37}, :1382:{5,13,47}, :1383:33, :1384:{45,56}, :1387:26, :1388:21, util.scala:118:51
  assign io_core_fencei_rdy =
    ~(stq_0_valid | stq_1_valid | stq_2_valid | stq_3_valid | stq_4_valid | stq_5_valid
      | stq_6_valid | stq_7_valid | stq_8_valid | stq_9_valid | stq_10_valid
      | stq_11_valid | stq_12_valid | stq_13_valid | stq_14_valid | stq_15_valid
      | stq_16_valid | stq_17_valid | stq_18_valid | stq_19_valid | stq_20_valid
      | stq_21_valid | stq_22_valid | stq_23_valid) & io_dmem_ordered;	// lsu.scala:211:16, :286:79, :348:{28,42}
  assign io_core_lxcpt_valid =
    r_xcpt_valid & ~io_core_exception
    & (io_core_brupdate_b1_mispredict_mask & r_xcpt_uop_br_mask) == 16'h0;	// lsu.scala:669:22, :1235:29, :1236:25, :1253:61, util.scala:118:{51,59}
  assign io_core_lxcpt_bits_uop_br_mask = r_xcpt_uop_br_mask;	// lsu.scala:1236:25
  assign io_core_lxcpt_bits_uop_rob_idx = r_xcpt_uop_rob_idx;	// lsu.scala:1236:25
  assign io_core_lxcpt_bits_cause = r_xcpt_cause;	// lsu.scala:1236:25
  assign io_core_lxcpt_bits_badvaddr = r_xcpt_badvaddr;	// lsu.scala:1236:25
  assign io_dmem_req_valid = dmem_req_0_valid;	// lsu.scala:766:39, :767:30, :773:43
  assign io_dmem_req_bits_0_valid = dmem_req_0_valid;	// lsu.scala:766:39, :767:30, :773:43
  assign io_dmem_req_bits_0_bits_uop_uopc =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_uopc
           : will_fire_load_retry_0
               ? _GEN_116[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_4[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_4[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_116[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_inst =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_inst
           : will_fire_load_retry_0
               ? _GEN_117[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_5[stq_retry_idx] : 32'h0)
      : will_fire_store_commit_0
          ? _GEN_5[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_117[ldq_wakeup_idx] : 32'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_inst =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_inst
           : will_fire_load_retry_0
               ? _GEN_118[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_6[stq_retry_idx] : 32'h0)
      : will_fire_store_commit_0
          ? _GEN_6[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_118[ldq_wakeup_idx] : 32'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_rvc =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_rvc
           : will_fire_load_retry_0
               ? _GEN_119[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_7[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_7[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_119[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_pc =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_pc
           : will_fire_load_retry_0
               ? _GEN_120[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_8[stq_retry_idx] : 40'h0)
      : will_fire_store_commit_0
          ? _GEN_8[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_120[ldq_wakeup_idx] : 40'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iq_type =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iq_type
           : will_fire_load_retry_0
               ? _GEN_121[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_9[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_9[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_121[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_fu_code =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_fu_code
           : will_fire_load_retry_0
               ? _GEN_122[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_10[stq_retry_idx] : 10'h0)
      : will_fire_store_commit_0
          ? _GEN_10[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_122[ldq_wakeup_idx] : 10'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_br_type =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_br_type
           : will_fire_load_retry_0
               ? _GEN_123[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_11[stq_retry_idx] : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_11[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_123[ldq_wakeup_idx] : 4'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_op1_sel =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_op1_sel
           : will_fire_load_retry_0
               ? _GEN_124[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_12[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_12[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_124[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_op2_sel =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_op2_sel
           : will_fire_load_retry_0
               ? _GEN_125[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_13[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_13[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_125[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_imm_sel =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_imm_sel
           : will_fire_load_retry_0
               ? _GEN_126[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_14[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_14[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_126[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_op_fcn =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_op_fcn
           : will_fire_load_retry_0
               ? _GEN_127[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_15[stq_retry_idx] : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_15[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_127[ldq_wakeup_idx] : 4'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_fcn_dw
           : will_fire_load_retry_0
               ? _GEN_128[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_16[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_16[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_128[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_csr_cmd
           : will_fire_load_retry_0
               ? _GEN_129[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_17[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_17[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_129[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_load =
    _GEN_315
      ? exe_tlb_uop_0_ctrl_is_load
      : will_fire_store_commit_0
          ? _GEN_18[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_130[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_sta =
    _GEN_315
      ? exe_tlb_uop_0_ctrl_is_sta
      : will_fire_store_commit_0
          ? _GEN_19[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_131[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_std =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_is_std
           : will_fire_load_retry_0
               ? _GEN_132[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_20[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_20[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_132[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iw_state =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iw_state
           : will_fire_load_retry_0
               ? _GEN_133[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_21[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_21[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_133[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iw_p1_poisoned =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iw_p1_poisoned
           : will_fire_load_retry_0
               ? _GEN_134[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_22[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_22[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_134[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iw_p2_poisoned =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iw_p2_poisoned
           : will_fire_load_retry_0
               ? _GEN_135[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_23[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_23[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_135[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_br =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_br
           : will_fire_load_retry_0
               ? _GEN_136[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_24[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_24[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_136[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_jalr =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_jalr
           : will_fire_load_retry_0
               ? _GEN_137[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_25[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_25[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_137[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_jal =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_jal
           : will_fire_load_retry_0
               ? _GEN_138[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_26[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_26[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_138[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_sfb =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_sfb
           : will_fire_load_retry_0
               ? _GEN_139[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_27[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_27[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_139[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_br_mask =
    _GEN_315
      ? exe_tlb_uop_0_br_mask
      : will_fire_store_commit_0
          ? _GEN_28[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_209 : 16'h0;	// lsu.scala:220:29, :224:42, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_br_tag =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_br_tag
           : will_fire_load_retry_0
               ? _GEN_141[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_29[stq_retry_idx] : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_29[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_141[ldq_wakeup_idx] : 4'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ftq_idx =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ftq_idx
           : will_fire_load_retry_0
               ? _GEN_142[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_30[stq_retry_idx] : 5'h0)
      : will_fire_store_commit_0
          ? _GEN_30[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_142[ldq_wakeup_idx] : 5'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_edge_inst =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_edge_inst
           : will_fire_load_retry_0
               ? _GEN_143[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_31[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_31[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_143[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_pc_lob =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_pc_lob
           : will_fire_load_retry_0
               ? _GEN_144[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_32[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_32[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_144[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_taken =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_taken
           : will_fire_load_retry_0
               ? _GEN_145[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_33[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_33[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_145[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_imm_packed =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_imm_packed
           : will_fire_load_retry_0
               ? _GEN_146[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_34[stq_retry_idx] : 20'h0)
      : will_fire_store_commit_0
          ? _GEN_34[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_146[ldq_wakeup_idx] : 20'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_csr_addr =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_csr_addr
           : will_fire_load_retry_0
               ? _GEN_147[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_35[stq_retry_idx] : 12'h0)
      : will_fire_store_commit_0
          ? _GEN_35[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_147[ldq_wakeup_idx] : 12'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_rob_idx =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_rob_idx
           : will_fire_load_retry_0
               ? _GEN_149
               : will_fire_sta_retry_0 ? mem_stq_retry_e_out_bits_uop_rob_idx : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_36[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_148[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldq_idx =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldq_idx
           : will_fire_load_retry_0 ? _GEN_151 : will_fire_sta_retry_0 ? _GEN_206 : 5'h0)
      : will_fire_store_commit_0
          ? _GEN_37[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_150[ldq_wakeup_idx] : 5'h0;	// lsu.scala:220:29, :224:42, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_stq_idx =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_stq_idx
           : will_fire_load_retry_0
               ? mem_ldq_retry_e_out_bits_uop_stq_idx
               : will_fire_sta_retry_0 ? mem_stq_retry_e_out_bits_uop_stq_idx : 5'h0)
      : will_fire_store_commit_0
          ? _GEN_38[stq_execute_head]
          : will_fire_load_wakeup_0 ? mem_ldq_wakeup_e_out_bits_uop_stq_idx : 5'h0;	// lsu.scala:220:29, :224:42, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_rxq_idx =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_rxq_idx
           : will_fire_load_retry_0
               ? _GEN_152[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_39[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_39[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_152[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_pdst =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_pdst
           : will_fire_load_retry_0 ? _GEN_154 : will_fire_sta_retry_0 ? _GEN_207 : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_40[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_153[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs1 =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs1
           : will_fire_load_retry_0
               ? _GEN_155[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_41[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_41[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_155[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs2 =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs2
           : will_fire_load_retry_0
               ? _GEN_156[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_42[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_42[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_156[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs3 =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs3
           : will_fire_load_retry_0
               ? _GEN_157[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_43[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_43[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_157[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ppred =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ppred
           : will_fire_load_retry_0
               ? _GEN_158[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_44[stq_retry_idx] : 5'h0)
      : will_fire_store_commit_0
          ? _GEN_44[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_158[ldq_wakeup_idx] : 5'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs1_busy =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs1_busy
           : will_fire_load_retry_0
               ? _GEN_159[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_45[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_45[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_159[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs2_busy =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs2_busy
           : will_fire_load_retry_0
               ? _GEN_160[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_46[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_46[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_160[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs3_busy =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs3_busy
           : will_fire_load_retry_0
               ? _GEN_161[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_47[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_47[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_161[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ppred_busy =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ppred_busy
           : will_fire_load_retry_0
               ? _GEN_162[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_48[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_48[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_162[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_stale_pdst =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_stale_pdst
           : will_fire_load_retry_0
               ? _GEN_163[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_49[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_49[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_163[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_exception =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_exception
           : will_fire_load_retry_0
               ? _GEN_164[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_50[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_51
          : will_fire_load_wakeup_0 & _GEN_164[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_exc_cause =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_exc_cause
           : will_fire_load_retry_0
               ? _GEN_165[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_52[stq_retry_idx] : 64'h0)
      : will_fire_store_commit_0
          ? _GEN_52[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_165[ldq_wakeup_idx] : 64'h0;	// AMOALU.scala:26:13, lsu.scala:220:29, :224:42, :249:20, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_bypassable =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_bypassable
           : will_fire_load_retry_0
               ? _GEN_166[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_53[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_53[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_166[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_mem_cmd =
    _GEN_315
      ? exe_tlb_uop_0_mem_cmd
      : will_fire_store_commit_0
          ? _GEN_54[stq_execute_head]
          : will_fire_load_wakeup_0
              ? _GEN_167[ldq_wakeup_idx]
              : _GEN_320 ? hella_req_cmd : 5'h0;	// lsu.scala:220:29, :224:42, :243:34, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, :802:47, :811:39, :819:5, :827:39
  assign io_dmem_req_bits_0_bits_uop_mem_size =
    _GEN_315
      ? exe_tlb_uop_0_mem_size
      : will_fire_store_commit_0
          ? _GEN_56
          : will_fire_load_wakeup_0
              ? mem_ldq_wakeup_e_out_bits_uop_mem_size
              : _GEN_320 ? hella_req_size : 2'h0;	// lsu.scala:220:29, :224:42, :243:34, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, :802:47, :811:39, :812:39, :819:5, :827:39, :828:39
  assign io_dmem_req_bits_0_bits_uop_mem_signed =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_mem_signed
           : will_fire_load_retry_0
               ? _GEN_168[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_57[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_57[stq_execute_head]
          : will_fire_load_wakeup_0
              ? _GEN_168[ldq_wakeup_idx]
              : _GEN_320 & hella_req_signed;	// lsu.scala:220:29, :224:42, :243:34, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, :802:47, :811:39, :813:39, :819:5, :827:39, :829:39
  assign io_dmem_req_bits_0_bits_uop_is_fence =
    _GEN_315
      ? exe_tlb_uop_0_is_fence
      : will_fire_store_commit_0
          ? _GEN_59
          : will_fire_load_wakeup_0 & _GEN_169[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_fencei =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_fencei
           : will_fire_load_retry_0
               ? _GEN_170[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_60[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_60[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_170[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_amo =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_amo
           : will_fire_load_retry_0
               ? _GEN_171[ldq_retry_idx]
               : will_fire_sta_retry_0 & mem_stq_retry_e_out_bits_uop_is_amo)
      : will_fire_store_commit_0
          ? _GEN_62
          : will_fire_load_wakeup_0 & _GEN_171[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_uses_ldq =
    _GEN_315
      ? _mem_xcpt_uops_WIRE_0_uses_ldq
      : will_fire_store_commit_0
          ? _GEN_63[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_172[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_uses_stq =
    _GEN_315
      ? _mem_xcpt_uops_WIRE_0_uses_stq
      : will_fire_store_commit_0
          ? _GEN_64[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_174[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_sys_pc2epc =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_sys_pc2epc
           : will_fire_load_retry_0
               ? _GEN_176[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_65[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_65[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_176[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_unique =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_unique
           : will_fire_load_retry_0
               ? _GEN_177[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_66[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_66[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_177[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_flush_on_commit =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_flush_on_commit
           : will_fire_load_retry_0
               ? _GEN_178[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_67[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_67[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_178[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldst_is_rs1 =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldst_is_rs1
           : will_fire_load_retry_0
               ? _GEN_179[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_68[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_68[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_179[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldst =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldst
           : will_fire_load_retry_0
               ? _GEN_180[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_69[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_69[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_180[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs1 =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs1
           : will_fire_load_retry_0
               ? _GEN_181[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_70[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_70[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_181[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs2 =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs2
           : will_fire_load_retry_0
               ? _GEN_182[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_71[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_71[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_182[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs3 =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs3
           : will_fire_load_retry_0
               ? _GEN_183[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_72[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_72[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_183[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldst_val =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldst_val
           : will_fire_load_retry_0
               ? _GEN_184[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_73[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_73[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_184[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_dst_rtype =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_dst_rtype
           : will_fire_load_retry_0
               ? _GEN_185[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_74[stq_retry_idx] : 2'h2)
      : will_fire_store_commit_0
          ? _GEN_74[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_185[ldq_wakeup_idx] : 2'h2;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, util.scala:351:72
  assign io_dmem_req_bits_0_bits_uop_lrs1_rtype =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs1_rtype
           : will_fire_load_retry_0
               ? _GEN_186[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_75[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_75[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_186[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs2_rtype =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs2_rtype
           : will_fire_load_retry_0
               ? _GEN_187[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_76[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_76[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_187[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_frs3_en =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_frs3_en
           : will_fire_load_retry_0
               ? _GEN_188[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_77[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_77[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_188[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_fp_val =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_fp_val
           : will_fire_load_retry_0
               ? _GEN_189[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_78[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_78[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_189[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_fp_single =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_fp_single
           : will_fire_load_retry_0
               ? _GEN_190[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_79[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_79[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_190[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_xcpt_pf_if =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_xcpt_pf_if
           : will_fire_load_retry_0
               ? _GEN_191[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_80[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_80[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_191[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_xcpt_ae_if =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_xcpt_ae_if
           : will_fire_load_retry_0
               ? _GEN_192[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_81[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_81[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_192[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_xcpt_ma_if =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_xcpt_ma_if
           : will_fire_load_retry_0
               ? _GEN_193[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_82[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_82[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_193[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_bp_debug_if =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_bp_debug_if
           : will_fire_load_retry_0
               ? _GEN_194[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_83[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_83[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_194[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_bp_xcpt_if =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_bp_xcpt_if
           : will_fire_load_retry_0
               ? _GEN_195[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_84[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_84[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_195[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_fsrc =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_fsrc
           : will_fire_load_retry_0
               ? _GEN_196[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_85[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_85[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_196[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_tsrc =
    _GEN_315
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_tsrc
           : will_fire_load_retry_0
               ? _GEN_197[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_86[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_86[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_197[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_addr =
    _GEN_318
      ? _GEN_313
      : will_fire_store_commit_0
          ? _GEN_89
          : will_fire_load_wakeup_0
              ? _GEN_210
              : will_fire_hella_incoming_0
                  ? _GEN_313
                  : will_fire_hella_wakeup_0 ? _GEN_317 : 40'h0;	// lsu.scala:224:42, :502:88, :535:65, :760:28, :766:39, :768:30, :773:43, :780:45, :782:33, :794:44, :796:30, :802:47, :806:39, :819:5, :822:39
  assign io_dmem_req_bits_0_bits_data =
    _GEN_315
      ? 64'h0
      : will_fire_store_commit_0
          ? _GEN_314[_GEN_56]
          : will_fire_load_wakeup_0 | will_fire_hella_incoming_0
            | ~will_fire_hella_wakeup_0
              ? 64'h0
              : _GEN_319[hella_req_size];	// AMOALU.scala:26:{13,19}, lsu.scala:220:29, :224:42, :243:34, :249:20, :535:65, :761:28, :766:39, :773:43, :780:45, :783:33, :794:44, :802:47, :807:39, :819:5
  assign io_dmem_req_bits_0_bits_is_hella =
    ~(_GEN_315 | will_fire_store_commit_0 | will_fire_load_wakeup_0)
    & (will_fire_hella_incoming_0 | will_fire_hella_wakeup_0);	// lsu.scala:220:29, :535:65, :762:31, :766:39, :773:43, :780:45, :794:44, :802:47, :814:39, :819:5
  assign io_dmem_s1_kill_0 =
    _GEN_753
      ? (_GEN_755
           ? io_dmem_s1_kill_0_REG_93
           : _GEN_756
               ? io_dmem_s1_kill_0_REG_94
               : _GEN_757 ? io_dmem_s1_kill_0_REG_95 : _GEN_751)
      : _GEN_751;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  assign io_dmem_brupdate_b1_resolve_mask = io_core_brupdate_b1_resolve_mask;
  assign io_dmem_brupdate_b1_mispredict_mask = io_core_brupdate_b1_mispredict_mask;
  assign io_dmem_exception = io_core_exception;
  assign io_dmem_release_ready = will_fire_release_0;	// lsu.scala:534:63
  assign io_dmem_force_order = _GEN_847 & _GEN_848 | io_core_fence_dmem;	// lsu.scala:347:25, :1494:29, :1495:3, :1496:{43,64}, :1497:27
  assign io_hellacache_req_ready = ~(|hella_state);	// lsu.scala:242:38, :593:24, :1527:21
  assign io_hellacache_s2_nack = ~_GEN_850 & _GEN_849;	// lsu.scala:1524:27, :1527:34, :1533:38, :1550:{28,43}
  assign io_hellacache_resp_valid =
    ~(_GEN_850 | _GEN_849 | _GEN_851) & _GEN_759 & _GEN_852;	// lsu.scala:1288:28, :1524:27, :1526:28, :1527:34, :1533:38, :1550:{28,43}, :1553:{28,38}, :1560:40, :1562:35
  assign io_hellacache_resp_bits_data = io_dmem_resp_0_bits_data;
  assign io_hellacache_s2_xcpt_ae_ld =
    ~(~(|hella_state) | _GEN_1 | _GEN_849) & _GEN_851 & hella_xcpt_ae_ld;	// lsu.scala:242:38, :246:34, :593:24, :803:26, :1525:27, :1527:{21,34}, :1533:38, :1550:{28,43}, :1553:{28,38}
endmodule

