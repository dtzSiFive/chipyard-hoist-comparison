// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module MemoryBus(
  input         auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready,
                auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid,
  input  [2:0]  auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode,
  input  [1:0]  auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param,
  input  [2:0]  auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size,
  input  [3:0]  auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source,
  input         auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink,
                auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied,
  input  [63:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data,
  input         auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt,
                auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready,
                auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready,
                auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid,
  input  [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id,
  input  [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp,
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready,
                auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid,
  input  [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id,
  input  [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data,
  input  [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp,
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last,
                auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock,
                auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset,
                auto_bus_xing_in_a_valid,
  input  [2:0]  auto_bus_xing_in_a_bits_opcode,
                auto_bus_xing_in_a_bits_param,
                auto_bus_xing_in_a_bits_size,
  input  [3:0]  auto_bus_xing_in_a_bits_source,
  input  [31:0] auto_bus_xing_in_a_bits_address,
  input  [7:0]  auto_bus_xing_in_a_bits_mask,
  input  [63:0] auto_bus_xing_in_a_bits_data,
  input         auto_bus_xing_in_a_bits_corrupt,
                auto_bus_xing_in_d_ready,
  output        auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid,
  output [28:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address,
  output        auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready,
                auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id,
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr,
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size,
  output [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid,
  output [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data,
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last,
                auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready,
                auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id,
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr,
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size,
  output [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready,
                auto_bus_xing_in_a_ready,
                auto_bus_xing_in_d_valid,
  output [2:0]  auto_bus_xing_in_d_bits_opcode,
  output [1:0]  auto_bus_xing_in_d_bits_param,
  output [2:0]  auto_bus_xing_in_d_bits_size,
  output [3:0]  auto_bus_xing_in_d_bits_source,
  output        auto_bus_xing_in_d_bits_sink,
                auto_bus_xing_in_d_bits_denied,
  output [63:0] auto_bus_xing_in_d_bits_data,
  output        auto_bus_xing_in_d_bits_corrupt
);

  wire        _coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready;	// LazyModule.scala:432:27
  wire        _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid;	// LazyModule.scala:432:27
  wire [2:0]  _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode;	// LazyModule.scala:432:27
  wire [2:0]  _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size;	// LazyModule.scala:432:27
  wire [3:0]  _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source;	// LazyModule.scala:432:27
  wire        _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied;	// LazyModule.scala:432:27
  wire        _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt;	// LazyModule.scala:432:27
  wire        _subsystem_mbus_xbar_auto_in_a_ready;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_in_d_valid;	// MemoryBus.scala:42:32
  wire [2:0]  _subsystem_mbus_xbar_auto_in_d_bits_opcode;	// MemoryBus.scala:42:32
  wire [1:0]  _subsystem_mbus_xbar_auto_in_d_bits_param;	// MemoryBus.scala:42:32
  wire [2:0]  _subsystem_mbus_xbar_auto_in_d_bits_size;	// MemoryBus.scala:42:32
  wire [3:0]  _subsystem_mbus_xbar_auto_in_d_bits_source;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_in_d_bits_sink;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_in_d_bits_denied;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_in_d_bits_corrupt;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_out_1_a_valid;	// MemoryBus.scala:42:32
  wire [28:0] _subsystem_mbus_xbar_auto_out_1_a_bits_address;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_out_1_d_ready;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_out_0_a_valid;	// MemoryBus.scala:42:32
  wire        _subsystem_mbus_xbar_auto_out_0_d_ready;	// MemoryBus.scala:42:32
  TLXbar_6 subsystem_mbus_xbar (	// MemoryBus.scala:42:32
    .clock
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),
    .reset
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),
    .auto_in_a_valid           (auto_bus_xing_in_a_valid),
    .auto_in_a_bits_opcode     (auto_bus_xing_in_a_bits_opcode),
    .auto_in_a_bits_param      (auto_bus_xing_in_a_bits_param),
    .auto_in_a_bits_size       (auto_bus_xing_in_a_bits_size),
    .auto_in_a_bits_source     (auto_bus_xing_in_a_bits_source),
    .auto_in_a_bits_address    (auto_bus_xing_in_a_bits_address),
    .auto_in_a_bits_mask       (auto_bus_xing_in_a_bits_mask),
    .auto_in_a_bits_corrupt    (auto_bus_xing_in_a_bits_corrupt),
    .auto_in_d_ready           (auto_bus_xing_in_d_ready),
    .auto_out_1_a_ready
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready),
    .auto_out_1_d_valid
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid),
    .auto_out_1_d_bits_opcode
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode),
    .auto_out_1_d_bits_param
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param),
    .auto_out_1_d_bits_size
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size),
    .auto_out_1_d_bits_source
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source),
    .auto_out_1_d_bits_sink
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink),
    .auto_out_1_d_bits_denied
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied),
    .auto_out_1_d_bits_data
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data),
    .auto_out_1_d_bits_corrupt
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt),
    .auto_out_0_a_ready
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready),	// LazyModule.scala:432:27
    .auto_out_0_d_valid
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_opcode
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_param   (2'h0),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_size
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_source
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_sink    (1'h0),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_denied
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_data
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data),
    .auto_out_0_d_bits_corrupt
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt),	// LazyModule.scala:432:27
    .auto_in_a_ready           (_subsystem_mbus_xbar_auto_in_a_ready),
    .auto_in_d_valid           (_subsystem_mbus_xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode     (_subsystem_mbus_xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param      (_subsystem_mbus_xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size       (_subsystem_mbus_xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source     (_subsystem_mbus_xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink       (_subsystem_mbus_xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied     (_subsystem_mbus_xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data       (auto_bus_xing_in_d_bits_data),
    .auto_in_d_bits_corrupt    (_subsystem_mbus_xbar_auto_in_d_bits_corrupt),
    .auto_out_1_a_valid        (_subsystem_mbus_xbar_auto_out_1_a_valid),
    .auto_out_1_a_bits_address (_subsystem_mbus_xbar_auto_out_1_a_bits_address),
    .auto_out_1_d_ready        (_subsystem_mbus_xbar_auto_out_1_d_ready),
    .auto_out_0_a_valid        (_subsystem_mbus_xbar_auto_out_0_a_valid),
    .auto_out_0_d_ready        (_subsystem_mbus_xbar_auto_out_0_d_ready)
  );
  TLFIFOFixer_3 fixer (	// FIFOFixer.scala:144:27
    .clock
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),
    .reset
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),
    .auto_in_a_valid         (auto_bus_xing_in_a_valid),
    .auto_in_a_bits_opcode   (auto_bus_xing_in_a_bits_opcode),
    .auto_in_a_bits_param    (auto_bus_xing_in_a_bits_param),
    .auto_in_a_bits_size     (auto_bus_xing_in_a_bits_size),
    .auto_in_a_bits_source   (auto_bus_xing_in_a_bits_source),
    .auto_in_a_bits_address  (auto_bus_xing_in_a_bits_address),
    .auto_in_a_bits_mask     (auto_bus_xing_in_a_bits_mask),
    .auto_in_a_bits_corrupt  (auto_bus_xing_in_a_bits_corrupt),
    .auto_in_d_ready         (auto_bus_xing_in_d_ready),
    .auto_out_a_ready        (_subsystem_mbus_xbar_auto_in_a_ready),	// MemoryBus.scala:42:32
    .auto_out_d_valid        (_subsystem_mbus_xbar_auto_in_d_valid),	// MemoryBus.scala:42:32
    .auto_out_d_bits_opcode  (_subsystem_mbus_xbar_auto_in_d_bits_opcode),	// MemoryBus.scala:42:32
    .auto_out_d_bits_param   (_subsystem_mbus_xbar_auto_in_d_bits_param),	// MemoryBus.scala:42:32
    .auto_out_d_bits_size    (_subsystem_mbus_xbar_auto_in_d_bits_size),	// MemoryBus.scala:42:32
    .auto_out_d_bits_source  (_subsystem_mbus_xbar_auto_in_d_bits_source),	// MemoryBus.scala:42:32
    .auto_out_d_bits_sink    (_subsystem_mbus_xbar_auto_in_d_bits_sink),	// MemoryBus.scala:42:32
    .auto_out_d_bits_denied  (_subsystem_mbus_xbar_auto_in_d_bits_denied),	// MemoryBus.scala:42:32
    .auto_out_d_bits_corrupt (_subsystem_mbus_xbar_auto_in_d_bits_corrupt)	// MemoryBus.scala:42:32
  );
  ProbePicker picker (	// ProbePicker.scala:65:28
    .clock
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),
    .reset
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),
    .auto_in_1_a_valid         (_subsystem_mbus_xbar_auto_out_1_a_valid),	// MemoryBus.scala:42:32
    .auto_in_1_a_bits_opcode   (auto_bus_xing_in_a_bits_opcode),
    .auto_in_1_a_bits_param    (auto_bus_xing_in_a_bits_param),
    .auto_in_1_a_bits_size     (auto_bus_xing_in_a_bits_size),
    .auto_in_1_a_bits_source   (auto_bus_xing_in_a_bits_source),
    .auto_in_1_a_bits_address  (_subsystem_mbus_xbar_auto_out_1_a_bits_address),	// MemoryBus.scala:42:32
    .auto_in_1_a_bits_mask     (auto_bus_xing_in_a_bits_mask),
    .auto_in_1_a_bits_corrupt  (auto_bus_xing_in_a_bits_corrupt),
    .auto_in_1_d_ready         (_subsystem_mbus_xbar_auto_out_1_d_ready),	// MemoryBus.scala:42:32
    .auto_in_0_a_valid         (_subsystem_mbus_xbar_auto_out_0_a_valid),	// MemoryBus.scala:42:32
    .auto_in_0_a_bits_opcode   (auto_bus_xing_in_a_bits_opcode),
    .auto_in_0_a_bits_param    (auto_bus_xing_in_a_bits_param),
    .auto_in_0_a_bits_size     (auto_bus_xing_in_a_bits_size),
    .auto_in_0_a_bits_source   (auto_bus_xing_in_a_bits_source),
    .auto_in_0_a_bits_address  (auto_bus_xing_in_a_bits_address),
    .auto_in_0_a_bits_mask     (auto_bus_xing_in_a_bits_mask),
    .auto_in_0_a_bits_corrupt  (auto_bus_xing_in_a_bits_corrupt),
    .auto_in_0_d_ready         (_subsystem_mbus_xbar_auto_out_0_d_ready),	// MemoryBus.scala:42:32
    .auto_out_1_a_ready
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready),
    .auto_out_1_d_valid
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid),
    .auto_out_1_d_bits_opcode
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode),
    .auto_out_1_d_bits_param
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param),
    .auto_out_1_d_bits_size
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size),
    .auto_out_1_d_bits_source
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source),
    .auto_out_1_d_bits_sink
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink),
    .auto_out_1_d_bits_denied
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied),
    .auto_out_1_d_bits_corrupt
      (auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt),
    .auto_out_0_a_ready
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready),	// LazyModule.scala:432:27
    .auto_out_0_d_valid
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_opcode
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_param   (2'h0),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_size
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_source
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_sink    (1'h0),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_denied
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied),	// LazyModule.scala:432:27
    .auto_out_0_d_bits_corrupt
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt)	// LazyModule.scala:432:27
  );
  TLInterconnectCoupler_27 coupler_to_memory_controller_port_named_axi4 (	// LazyModule.scala:432:27
    .clock
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),
    .reset
      (auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),
    .auto_axi4yank_out_aw_ready
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready),
    .auto_axi4yank_out_w_ready
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready),
    .auto_axi4yank_out_b_valid
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid),
    .auto_axi4yank_out_b_bits_id
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id),
    .auto_axi4yank_out_b_bits_resp
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp),
    .auto_axi4yank_out_ar_ready
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready),
    .auto_axi4yank_out_r_valid
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid),
    .auto_axi4yank_out_r_bits_id
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id),
    .auto_axi4yank_out_r_bits_resp
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp),
    .auto_axi4yank_out_r_bits_last
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last),
    .auto_tl_in_a_valid              (_subsystem_mbus_xbar_auto_out_0_a_valid),	// MemoryBus.scala:42:32
    .auto_tl_in_a_bits_opcode        (auto_bus_xing_in_a_bits_opcode),
    .auto_tl_in_a_bits_param         (auto_bus_xing_in_a_bits_param),
    .auto_tl_in_a_bits_size          (auto_bus_xing_in_a_bits_size),
    .auto_tl_in_a_bits_source        (auto_bus_xing_in_a_bits_source),
    .auto_tl_in_a_bits_address       (auto_bus_xing_in_a_bits_address),
    .auto_tl_in_a_bits_mask          (auto_bus_xing_in_a_bits_mask),
    .auto_tl_in_a_bits_data          (auto_bus_xing_in_a_bits_data),
    .auto_tl_in_a_bits_corrupt       (auto_bus_xing_in_a_bits_corrupt),
    .auto_tl_in_d_ready              (_subsystem_mbus_xbar_auto_out_0_d_ready),	// MemoryBus.scala:42:32
    .auto_axi4yank_out_aw_valid
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid),
    .auto_axi4yank_out_aw_bits_id
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id),
    .auto_axi4yank_out_aw_bits_addr
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr),
    .auto_axi4yank_out_aw_bits_len
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len),
    .auto_axi4yank_out_aw_bits_size
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size),
    .auto_axi4yank_out_aw_bits_burst
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst),
    .auto_axi4yank_out_aw_bits_lock
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock),
    .auto_axi4yank_out_aw_bits_cache
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache),
    .auto_axi4yank_out_aw_bits_prot
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot),
    .auto_axi4yank_out_aw_bits_qos
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos),
    .auto_axi4yank_out_w_valid
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid),
    .auto_axi4yank_out_w_bits_data
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data),
    .auto_axi4yank_out_w_bits_strb
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb),
    .auto_axi4yank_out_w_bits_last
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last),
    .auto_axi4yank_out_b_ready
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready),
    .auto_axi4yank_out_ar_valid
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid),
    .auto_axi4yank_out_ar_bits_id
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id),
    .auto_axi4yank_out_ar_bits_addr
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr),
    .auto_axi4yank_out_ar_bits_len
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len),
    .auto_axi4yank_out_ar_bits_size
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size),
    .auto_axi4yank_out_ar_bits_burst
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst),
    .auto_axi4yank_out_ar_bits_lock
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock),
    .auto_axi4yank_out_ar_bits_cache
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache),
    .auto_axi4yank_out_ar_bits_prot
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot),
    .auto_axi4yank_out_ar_bits_qos
      (auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos),
    .auto_tl_in_a_ready
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready),
    .auto_tl_in_d_valid
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_opcode
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode),
    .auto_tl_in_d_bits_size
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_denied
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied),
    .auto_tl_in_d_bits_corrupt
      (_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt)
  );
  assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid =
    _subsystem_mbus_xbar_auto_out_1_a_valid;	// MemoryBus.scala:42:32
  assign
    auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address
    = _subsystem_mbus_xbar_auto_out_1_a_bits_address;	// MemoryBus.scala:42:32
  assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready =
    _subsystem_mbus_xbar_auto_out_1_d_ready;	// MemoryBus.scala:42:32
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready =
    _subsystem_mbus_xbar_auto_out_0_d_ready;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_a_ready = _subsystem_mbus_xbar_auto_in_a_ready;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_valid = _subsystem_mbus_xbar_auto_in_d_valid;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_bits_opcode = _subsystem_mbus_xbar_auto_in_d_bits_opcode;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_bits_param = _subsystem_mbus_xbar_auto_in_d_bits_param;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_bits_size = _subsystem_mbus_xbar_auto_in_d_bits_size;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_bits_source = _subsystem_mbus_xbar_auto_in_d_bits_source;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_bits_sink = _subsystem_mbus_xbar_auto_in_d_bits_sink;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_bits_denied = _subsystem_mbus_xbar_auto_in_d_bits_denied;	// MemoryBus.scala:42:32
  assign auto_bus_xing_in_d_bits_corrupt = _subsystem_mbus_xbar_auto_in_d_bits_corrupt;	// MemoryBus.scala:42:32
endmodule

