// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module LSU_2(
  input         clock,
                reset,
                io_ptw_req_ready,
                io_ptw_resp_valid,
                io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
                io_ptw_resp_bits_pte_a,
                io_ptw_resp_bits_pte_g,
                io_ptw_resp_bits_pte_u,
                io_ptw_resp_bits_pte_x,
                io_ptw_resp_bits_pte_w,
                io_ptw_resp_bits_pte_r,
                io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
                io_ptw_status_sum,
                io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
                io_ptw_pmp_0_cfg_w,
                io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
                io_ptw_pmp_1_cfg_w,
                io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
                io_ptw_pmp_2_cfg_w,
                io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
                io_ptw_pmp_3_cfg_w,
                io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
                io_ptw_pmp_4_cfg_w,
                io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
                io_ptw_pmp_5_cfg_w,
                io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
                io_ptw_pmp_6_cfg_w,
                io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
                io_ptw_pmp_7_cfg_w,
                io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_core_exe_0_req_valid,
  input  [6:0]  io_core_exe_0_req_bits_uop_uopc,
  input  [31:0] io_core_exe_0_req_bits_uop_inst,
                io_core_exe_0_req_bits_uop_debug_inst,
  input         io_core_exe_0_req_bits_uop_is_rvc,
  input  [39:0] io_core_exe_0_req_bits_uop_debug_pc,
  input  [2:0]  io_core_exe_0_req_bits_uop_iq_type,
  input  [9:0]  io_core_exe_0_req_bits_uop_fu_code,
  input  [3:0]  io_core_exe_0_req_bits_uop_ctrl_br_type,
  input  [1:0]  io_core_exe_0_req_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_core_exe_0_req_bits_uop_ctrl_op2_sel,
                io_core_exe_0_req_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_core_exe_0_req_bits_uop_ctrl_op_fcn,
  input         io_core_exe_0_req_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_core_exe_0_req_bits_uop_ctrl_csr_cmd,
  input         io_core_exe_0_req_bits_uop_ctrl_is_load,
                io_core_exe_0_req_bits_uop_ctrl_is_sta,
                io_core_exe_0_req_bits_uop_ctrl_is_std,
  input  [1:0]  io_core_exe_0_req_bits_uop_iw_state,
  input         io_core_exe_0_req_bits_uop_iw_p1_poisoned,
                io_core_exe_0_req_bits_uop_iw_p2_poisoned,
                io_core_exe_0_req_bits_uop_is_br,
                io_core_exe_0_req_bits_uop_is_jalr,
                io_core_exe_0_req_bits_uop_is_jal,
                io_core_exe_0_req_bits_uop_is_sfb,
  input  [11:0] io_core_exe_0_req_bits_uop_br_mask,
  input  [3:0]  io_core_exe_0_req_bits_uop_br_tag,
  input  [4:0]  io_core_exe_0_req_bits_uop_ftq_idx,
  input         io_core_exe_0_req_bits_uop_edge_inst,
  input  [5:0]  io_core_exe_0_req_bits_uop_pc_lob,
  input         io_core_exe_0_req_bits_uop_taken,
  input  [19:0] io_core_exe_0_req_bits_uop_imm_packed,
  input  [11:0] io_core_exe_0_req_bits_uop_csr_addr,
  input  [5:0]  io_core_exe_0_req_bits_uop_rob_idx,
  input  [3:0]  io_core_exe_0_req_bits_uop_ldq_idx,
                io_core_exe_0_req_bits_uop_stq_idx,
  input  [1:0]  io_core_exe_0_req_bits_uop_rxq_idx,
  input  [6:0]  io_core_exe_0_req_bits_uop_pdst,
                io_core_exe_0_req_bits_uop_prs1,
                io_core_exe_0_req_bits_uop_prs2,
                io_core_exe_0_req_bits_uop_prs3,
  input  [4:0]  io_core_exe_0_req_bits_uop_ppred,
  input         io_core_exe_0_req_bits_uop_prs1_busy,
                io_core_exe_0_req_bits_uop_prs2_busy,
                io_core_exe_0_req_bits_uop_prs3_busy,
                io_core_exe_0_req_bits_uop_ppred_busy,
  input  [6:0]  io_core_exe_0_req_bits_uop_stale_pdst,
  input         io_core_exe_0_req_bits_uop_exception,
  input  [63:0] io_core_exe_0_req_bits_uop_exc_cause,
  input         io_core_exe_0_req_bits_uop_bypassable,
  input  [4:0]  io_core_exe_0_req_bits_uop_mem_cmd,
  input  [1:0]  io_core_exe_0_req_bits_uop_mem_size,
  input         io_core_exe_0_req_bits_uop_mem_signed,
                io_core_exe_0_req_bits_uop_is_fence,
                io_core_exe_0_req_bits_uop_is_fencei,
                io_core_exe_0_req_bits_uop_is_amo,
                io_core_exe_0_req_bits_uop_uses_ldq,
                io_core_exe_0_req_bits_uop_uses_stq,
                io_core_exe_0_req_bits_uop_is_sys_pc2epc,
                io_core_exe_0_req_bits_uop_is_unique,
                io_core_exe_0_req_bits_uop_flush_on_commit,
                io_core_exe_0_req_bits_uop_ldst_is_rs1,
  input  [5:0]  io_core_exe_0_req_bits_uop_ldst,
                io_core_exe_0_req_bits_uop_lrs1,
                io_core_exe_0_req_bits_uop_lrs2,
                io_core_exe_0_req_bits_uop_lrs3,
  input         io_core_exe_0_req_bits_uop_ldst_val,
  input  [1:0]  io_core_exe_0_req_bits_uop_dst_rtype,
                io_core_exe_0_req_bits_uop_lrs1_rtype,
                io_core_exe_0_req_bits_uop_lrs2_rtype,
  input         io_core_exe_0_req_bits_uop_frs3_en,
                io_core_exe_0_req_bits_uop_fp_val,
                io_core_exe_0_req_bits_uop_fp_single,
                io_core_exe_0_req_bits_uop_xcpt_pf_if,
                io_core_exe_0_req_bits_uop_xcpt_ae_if,
                io_core_exe_0_req_bits_uop_xcpt_ma_if,
                io_core_exe_0_req_bits_uop_bp_debug_if,
                io_core_exe_0_req_bits_uop_bp_xcpt_if,
  input  [1:0]  io_core_exe_0_req_bits_uop_debug_fsrc,
                io_core_exe_0_req_bits_uop_debug_tsrc,
  input  [63:0] io_core_exe_0_req_bits_data,
  input  [39:0] io_core_exe_0_req_bits_addr,
  input         io_core_exe_0_req_bits_mxcpt_valid,
                io_core_exe_0_req_bits_sfence_valid,
                io_core_exe_0_req_bits_sfence_bits_rs1,
                io_core_exe_0_req_bits_sfence_bits_rs2,
  input  [38:0] io_core_exe_0_req_bits_sfence_bits_addr,
  input         io_core_dis_uops_0_valid,
  input  [6:0]  io_core_dis_uops_0_bits_uopc,
  input  [31:0] io_core_dis_uops_0_bits_inst,
                io_core_dis_uops_0_bits_debug_inst,
  input         io_core_dis_uops_0_bits_is_rvc,
  input  [39:0] io_core_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_0_bits_iq_type,
  input  [9:0]  io_core_dis_uops_0_bits_fu_code,
  input  [3:0]  io_core_dis_uops_0_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_0_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_0_bits_ctrl_op2_sel,
                io_core_dis_uops_0_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_0_bits_ctrl_op_fcn,
  input         io_core_dis_uops_0_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_0_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_0_bits_ctrl_is_load,
                io_core_dis_uops_0_bits_ctrl_is_sta,
                io_core_dis_uops_0_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_0_bits_iw_state,
  input         io_core_dis_uops_0_bits_iw_p1_poisoned,
                io_core_dis_uops_0_bits_iw_p2_poisoned,
                io_core_dis_uops_0_bits_is_br,
                io_core_dis_uops_0_bits_is_jalr,
                io_core_dis_uops_0_bits_is_jal,
                io_core_dis_uops_0_bits_is_sfb,
  input  [11:0] io_core_dis_uops_0_bits_br_mask,
  input  [3:0]  io_core_dis_uops_0_bits_br_tag,
  input  [4:0]  io_core_dis_uops_0_bits_ftq_idx,
  input         io_core_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_0_bits_pc_lob,
  input         io_core_dis_uops_0_bits_taken,
  input  [19:0] io_core_dis_uops_0_bits_imm_packed,
  input  [11:0] io_core_dis_uops_0_bits_csr_addr,
  input  [5:0]  io_core_dis_uops_0_bits_rob_idx,
  input  [3:0]  io_core_dis_uops_0_bits_ldq_idx,
                io_core_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_0_bits_pdst,
                io_core_dis_uops_0_bits_prs1,
                io_core_dis_uops_0_bits_prs2,
                io_core_dis_uops_0_bits_prs3,
  input         io_core_dis_uops_0_bits_prs1_busy,
                io_core_dis_uops_0_bits_prs2_busy,
                io_core_dis_uops_0_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_0_bits_stale_pdst,
  input         io_core_dis_uops_0_bits_exception,
  input  [63:0] io_core_dis_uops_0_bits_exc_cause,
  input         io_core_dis_uops_0_bits_bypassable,
  input  [4:0]  io_core_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_0_bits_mem_size,
  input         io_core_dis_uops_0_bits_mem_signed,
                io_core_dis_uops_0_bits_is_fence,
                io_core_dis_uops_0_bits_is_fencei,
                io_core_dis_uops_0_bits_is_amo,
                io_core_dis_uops_0_bits_uses_ldq,
                io_core_dis_uops_0_bits_uses_stq,
                io_core_dis_uops_0_bits_is_sys_pc2epc,
                io_core_dis_uops_0_bits_is_unique,
                io_core_dis_uops_0_bits_flush_on_commit,
                io_core_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_0_bits_ldst,
                io_core_dis_uops_0_bits_lrs1,
                io_core_dis_uops_0_bits_lrs2,
                io_core_dis_uops_0_bits_lrs3,
  input         io_core_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_0_bits_dst_rtype,
                io_core_dis_uops_0_bits_lrs1_rtype,
                io_core_dis_uops_0_bits_lrs2_rtype,
  input         io_core_dis_uops_0_bits_frs3_en,
                io_core_dis_uops_0_bits_fp_val,
                io_core_dis_uops_0_bits_fp_single,
                io_core_dis_uops_0_bits_xcpt_pf_if,
                io_core_dis_uops_0_bits_xcpt_ae_if,
                io_core_dis_uops_0_bits_xcpt_ma_if,
                io_core_dis_uops_0_bits_bp_debug_if,
                io_core_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_0_bits_debug_fsrc,
                io_core_dis_uops_0_bits_debug_tsrc,
  input         io_core_dis_uops_1_valid,
  input  [6:0]  io_core_dis_uops_1_bits_uopc,
  input  [31:0] io_core_dis_uops_1_bits_inst,
                io_core_dis_uops_1_bits_debug_inst,
  input         io_core_dis_uops_1_bits_is_rvc,
  input  [39:0] io_core_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_1_bits_iq_type,
  input  [9:0]  io_core_dis_uops_1_bits_fu_code,
  input  [3:0]  io_core_dis_uops_1_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_1_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_1_bits_ctrl_op2_sel,
                io_core_dis_uops_1_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_1_bits_ctrl_op_fcn,
  input         io_core_dis_uops_1_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_1_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_1_bits_ctrl_is_load,
                io_core_dis_uops_1_bits_ctrl_is_sta,
                io_core_dis_uops_1_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_1_bits_iw_state,
  input         io_core_dis_uops_1_bits_iw_p1_poisoned,
                io_core_dis_uops_1_bits_iw_p2_poisoned,
                io_core_dis_uops_1_bits_is_br,
                io_core_dis_uops_1_bits_is_jalr,
                io_core_dis_uops_1_bits_is_jal,
                io_core_dis_uops_1_bits_is_sfb,
  input  [11:0] io_core_dis_uops_1_bits_br_mask,
  input  [3:0]  io_core_dis_uops_1_bits_br_tag,
  input  [4:0]  io_core_dis_uops_1_bits_ftq_idx,
  input         io_core_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_1_bits_pc_lob,
  input         io_core_dis_uops_1_bits_taken,
  input  [19:0] io_core_dis_uops_1_bits_imm_packed,
  input  [11:0] io_core_dis_uops_1_bits_csr_addr,
  input  [5:0]  io_core_dis_uops_1_bits_rob_idx,
  input  [3:0]  io_core_dis_uops_1_bits_ldq_idx,
                io_core_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_1_bits_pdst,
                io_core_dis_uops_1_bits_prs1,
                io_core_dis_uops_1_bits_prs2,
                io_core_dis_uops_1_bits_prs3,
  input         io_core_dis_uops_1_bits_prs1_busy,
                io_core_dis_uops_1_bits_prs2_busy,
                io_core_dis_uops_1_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_1_bits_stale_pdst,
  input         io_core_dis_uops_1_bits_exception,
  input  [63:0] io_core_dis_uops_1_bits_exc_cause,
  input         io_core_dis_uops_1_bits_bypassable,
  input  [4:0]  io_core_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_1_bits_mem_size,
  input         io_core_dis_uops_1_bits_mem_signed,
                io_core_dis_uops_1_bits_is_fence,
                io_core_dis_uops_1_bits_is_fencei,
                io_core_dis_uops_1_bits_is_amo,
                io_core_dis_uops_1_bits_uses_ldq,
                io_core_dis_uops_1_bits_uses_stq,
                io_core_dis_uops_1_bits_is_sys_pc2epc,
                io_core_dis_uops_1_bits_is_unique,
                io_core_dis_uops_1_bits_flush_on_commit,
                io_core_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_1_bits_ldst,
                io_core_dis_uops_1_bits_lrs1,
                io_core_dis_uops_1_bits_lrs2,
                io_core_dis_uops_1_bits_lrs3,
  input         io_core_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_1_bits_dst_rtype,
                io_core_dis_uops_1_bits_lrs1_rtype,
                io_core_dis_uops_1_bits_lrs2_rtype,
  input         io_core_dis_uops_1_bits_frs3_en,
                io_core_dis_uops_1_bits_fp_val,
                io_core_dis_uops_1_bits_fp_single,
                io_core_dis_uops_1_bits_xcpt_pf_if,
                io_core_dis_uops_1_bits_xcpt_ae_if,
                io_core_dis_uops_1_bits_xcpt_ma_if,
                io_core_dis_uops_1_bits_bp_debug_if,
                io_core_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_1_bits_debug_fsrc,
                io_core_dis_uops_1_bits_debug_tsrc,
  input         io_core_fp_stdata_valid,
  input  [11:0] io_core_fp_stdata_bits_uop_br_mask,
  input  [5:0]  io_core_fp_stdata_bits_uop_rob_idx,
  input  [3:0]  io_core_fp_stdata_bits_uop_stq_idx,
  input  [63:0] io_core_fp_stdata_bits_data,
  input         io_core_commit_valids_0,
                io_core_commit_valids_1,
                io_core_commit_uops_0_uses_ldq,
                io_core_commit_uops_0_uses_stq,
                io_core_commit_uops_1_uses_ldq,
                io_core_commit_uops_1_uses_stq,
                io_core_commit_load_at_rob_head,
                io_core_fence_dmem,
  input  [11:0] io_core_brupdate_b1_resolve_mask,
                io_core_brupdate_b1_mispredict_mask,
  input  [3:0]  io_core_brupdate_b2_uop_ldq_idx,
                io_core_brupdate_b2_uop_stq_idx,
  input         io_core_brupdate_b2_mispredict,
  input  [5:0]  io_core_rob_head_idx,
  input         io_core_exception,
                io_dmem_req_ready,
                io_dmem_resp_0_valid,
  input  [3:0]  io_dmem_resp_0_bits_uop_ldq_idx,
                io_dmem_resp_0_bits_uop_stq_idx,
  input         io_dmem_resp_0_bits_uop_is_amo,
                io_dmem_resp_0_bits_uop_uses_ldq,
                io_dmem_resp_0_bits_uop_uses_stq,
  input  [63:0] io_dmem_resp_0_bits_data,
  input         io_dmem_resp_0_bits_is_hella,
                io_dmem_nack_0_valid,
  input  [3:0]  io_dmem_nack_0_bits_uop_ldq_idx,
                io_dmem_nack_0_bits_uop_stq_idx,
  input         io_dmem_nack_0_bits_uop_uses_ldq,
                io_dmem_nack_0_bits_uop_uses_stq,
                io_dmem_nack_0_bits_is_hella,
                io_dmem_release_valid,
  input  [31:0] io_dmem_release_bits_address,
  input         io_dmem_ordered,
                io_hellacache_req_valid,
  input  [39:0] io_hellacache_req_bits_addr,
  input         io_hellacache_s1_kill,
  output        io_ptw_req_valid,
                io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  output        io_core_exe_0_iresp_valid,
  output [5:0]  io_core_exe_0_iresp_bits_uop_rob_idx,
  output [6:0]  io_core_exe_0_iresp_bits_uop_pdst,
  output        io_core_exe_0_iresp_bits_uop_is_amo,
                io_core_exe_0_iresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_iresp_bits_uop_dst_rtype,
  output [63:0] io_core_exe_0_iresp_bits_data,
  output        io_core_exe_0_fresp_valid,
  output [6:0]  io_core_exe_0_fresp_bits_uop_uopc,
  output [11:0] io_core_exe_0_fresp_bits_uop_br_mask,
  output [5:0]  io_core_exe_0_fresp_bits_uop_rob_idx,
  output [3:0]  io_core_exe_0_fresp_bits_uop_stq_idx,
  output [6:0]  io_core_exe_0_fresp_bits_uop_pdst,
  output [1:0]  io_core_exe_0_fresp_bits_uop_mem_size,
  output        io_core_exe_0_fresp_bits_uop_is_amo,
                io_core_exe_0_fresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_fresp_bits_uop_dst_rtype,
  output        io_core_exe_0_fresp_bits_uop_fp_val,
  output [64:0] io_core_exe_0_fresp_bits_data,
  output [3:0]  io_core_dis_ldq_idx_0,
                io_core_dis_ldq_idx_1,
                io_core_dis_stq_idx_0,
                io_core_dis_stq_idx_1,
  output        io_core_ldq_full_0,
                io_core_ldq_full_1,
                io_core_stq_full_0,
                io_core_stq_full_1,
                io_core_fp_stdata_ready,
                io_core_clr_bsy_0_valid,
  output [5:0]  io_core_clr_bsy_0_bits,
  output        io_core_clr_bsy_1_valid,
  output [5:0]  io_core_clr_bsy_1_bits,
  output        io_core_spec_ld_wakeup_0_valid,
  output [6:0]  io_core_spec_ld_wakeup_0_bits,
  output        io_core_ld_miss,
                io_core_fencei_rdy,
                io_core_lxcpt_valid,
  output [11:0] io_core_lxcpt_bits_uop_br_mask,
  output [5:0]  io_core_lxcpt_bits_uop_rob_idx,
  output [4:0]  io_core_lxcpt_bits_cause,
  output [39:0] io_core_lxcpt_bits_badvaddr,
  output        io_core_perf_tlbMiss,
                io_dmem_req_valid,
                io_dmem_req_bits_0_valid,
  output [6:0]  io_dmem_req_bits_0_bits_uop_uopc,
  output [31:0] io_dmem_req_bits_0_bits_uop_inst,
                io_dmem_req_bits_0_bits_uop_debug_inst,
  output        io_dmem_req_bits_0_bits_uop_is_rvc,
  output [39:0] io_dmem_req_bits_0_bits_uop_debug_pc,
  output [2:0]  io_dmem_req_bits_0_bits_uop_iq_type,
  output [9:0]  io_dmem_req_bits_0_bits_uop_fu_code,
  output [3:0]  io_dmem_req_bits_0_bits_uop_ctrl_br_type,
  output [1:0]  io_dmem_req_bits_0_bits_uop_ctrl_op1_sel,
  output [2:0]  io_dmem_req_bits_0_bits_uop_ctrl_op2_sel,
                io_dmem_req_bits_0_bits_uop_ctrl_imm_sel,
  output [3:0]  io_dmem_req_bits_0_bits_uop_ctrl_op_fcn,
  output        io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd,
  output        io_dmem_req_bits_0_bits_uop_ctrl_is_load,
                io_dmem_req_bits_0_bits_uop_ctrl_is_sta,
                io_dmem_req_bits_0_bits_uop_ctrl_is_std,
  output [1:0]  io_dmem_req_bits_0_bits_uop_iw_state,
  output        io_dmem_req_bits_0_bits_uop_iw_p1_poisoned,
                io_dmem_req_bits_0_bits_uop_iw_p2_poisoned,
                io_dmem_req_bits_0_bits_uop_is_br,
                io_dmem_req_bits_0_bits_uop_is_jalr,
                io_dmem_req_bits_0_bits_uop_is_jal,
                io_dmem_req_bits_0_bits_uop_is_sfb,
  output [11:0] io_dmem_req_bits_0_bits_uop_br_mask,
  output [3:0]  io_dmem_req_bits_0_bits_uop_br_tag,
  output [4:0]  io_dmem_req_bits_0_bits_uop_ftq_idx,
  output        io_dmem_req_bits_0_bits_uop_edge_inst,
  output [5:0]  io_dmem_req_bits_0_bits_uop_pc_lob,
  output        io_dmem_req_bits_0_bits_uop_taken,
  output [19:0] io_dmem_req_bits_0_bits_uop_imm_packed,
  output [11:0] io_dmem_req_bits_0_bits_uop_csr_addr,
  output [5:0]  io_dmem_req_bits_0_bits_uop_rob_idx,
  output [3:0]  io_dmem_req_bits_0_bits_uop_ldq_idx,
                io_dmem_req_bits_0_bits_uop_stq_idx,
  output [1:0]  io_dmem_req_bits_0_bits_uop_rxq_idx,
  output [6:0]  io_dmem_req_bits_0_bits_uop_pdst,
                io_dmem_req_bits_0_bits_uop_prs1,
                io_dmem_req_bits_0_bits_uop_prs2,
                io_dmem_req_bits_0_bits_uop_prs3,
  output [4:0]  io_dmem_req_bits_0_bits_uop_ppred,
  output        io_dmem_req_bits_0_bits_uop_prs1_busy,
                io_dmem_req_bits_0_bits_uop_prs2_busy,
                io_dmem_req_bits_0_bits_uop_prs3_busy,
                io_dmem_req_bits_0_bits_uop_ppred_busy,
  output [6:0]  io_dmem_req_bits_0_bits_uop_stale_pdst,
  output        io_dmem_req_bits_0_bits_uop_exception,
  output [63:0] io_dmem_req_bits_0_bits_uop_exc_cause,
  output        io_dmem_req_bits_0_bits_uop_bypassable,
  output [4:0]  io_dmem_req_bits_0_bits_uop_mem_cmd,
  output [1:0]  io_dmem_req_bits_0_bits_uop_mem_size,
  output        io_dmem_req_bits_0_bits_uop_mem_signed,
                io_dmem_req_bits_0_bits_uop_is_fence,
                io_dmem_req_bits_0_bits_uop_is_fencei,
                io_dmem_req_bits_0_bits_uop_is_amo,
                io_dmem_req_bits_0_bits_uop_uses_ldq,
                io_dmem_req_bits_0_bits_uop_uses_stq,
                io_dmem_req_bits_0_bits_uop_is_sys_pc2epc,
                io_dmem_req_bits_0_bits_uop_is_unique,
                io_dmem_req_bits_0_bits_uop_flush_on_commit,
                io_dmem_req_bits_0_bits_uop_ldst_is_rs1,
  output [5:0]  io_dmem_req_bits_0_bits_uop_ldst,
                io_dmem_req_bits_0_bits_uop_lrs1,
                io_dmem_req_bits_0_bits_uop_lrs2,
                io_dmem_req_bits_0_bits_uop_lrs3,
  output        io_dmem_req_bits_0_bits_uop_ldst_val,
  output [1:0]  io_dmem_req_bits_0_bits_uop_dst_rtype,
                io_dmem_req_bits_0_bits_uop_lrs1_rtype,
                io_dmem_req_bits_0_bits_uop_lrs2_rtype,
  output        io_dmem_req_bits_0_bits_uop_frs3_en,
                io_dmem_req_bits_0_bits_uop_fp_val,
                io_dmem_req_bits_0_bits_uop_fp_single,
                io_dmem_req_bits_0_bits_uop_xcpt_pf_if,
                io_dmem_req_bits_0_bits_uop_xcpt_ae_if,
                io_dmem_req_bits_0_bits_uop_xcpt_ma_if,
                io_dmem_req_bits_0_bits_uop_bp_debug_if,
                io_dmem_req_bits_0_bits_uop_bp_xcpt_if,
  output [1:0]  io_dmem_req_bits_0_bits_uop_debug_fsrc,
                io_dmem_req_bits_0_bits_uop_debug_tsrc,
  output [39:0] io_dmem_req_bits_0_bits_addr,
  output [63:0] io_dmem_req_bits_0_bits_data,
  output        io_dmem_req_bits_0_bits_is_hella,
                io_dmem_s1_kill_0,
                io_dmem_release_ready,
                io_dmem_force_order,
                io_hellacache_req_ready,
                io_hellacache_s2_nack,
                io_hellacache_resp_valid,
                io_hellacache_s2_xcpt_ae_ld
);

  wire              _GEN;	// lsu.scala:1527:34, :1533:38, :1550:43, :1553:38, :1560:40, :1576:42
  wire              store_needs_order;	// lsu.scala:1495:3, :1496:64
  wire              nacking_loads_15;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_14;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_13;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_12;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_11;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_10;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_9;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_8;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_7;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_6;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_5;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_4;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_3;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_2;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_1;	// lsu.scala:1284:5, :1287:7
  wire              nacking_loads_0;	// lsu.scala:1284:5, :1287:7
  wire              block_load_wakeup;	// lsu.scala:1199:80, :1210:43, :1211:25
  wire              _GEN_0;	// lsu.scala:820:26
  wire              _GEN_1;	// lsu.scala:803:26
  reg               mem_xcpt_valids_0;	// lsu.scala:667:32
  wire              _will_fire_store_commit_0_T_2;	// lsu.scala:538:31
  wire [3:0]        _forwarding_age_logic_0_io_forwarding_idx;	// lsu.scala:1178:57
  wire              _dtlb_io_miss_rdy;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_miss;	// lsu.scala:249:20
  wire [31:0]       _dtlb_io_resp_0_paddr;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_pf_ld;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_pf_st;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ae_ld;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ae_st;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ma_ld;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_ma_st;	// lsu.scala:249:20
  wire              _dtlb_io_resp_0_cacheable;	// lsu.scala:249:20
  wire              _dtlb_io_ptw_req_valid;	// lsu.scala:249:20
  reg               ldq_0_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_0_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_0_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_0_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_0_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_0_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_0_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_0_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_0_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_0_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_0_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_0_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_0_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_0_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_0_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_0_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_0_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_0_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_0_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_0_bits_executed;	// lsu.scala:210:16
  reg               ldq_0_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_0_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_0_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_0_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_0_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_0_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_1_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_1_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_1_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_1_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_1_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_1_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_1_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_1_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_1_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_1_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_1_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_1_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_1_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_1_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_1_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_1_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_1_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_1_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_1_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_1_bits_executed;	// lsu.scala:210:16
  reg               ldq_1_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_1_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_1_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_1_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_1_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_1_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_2_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_2_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_2_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_2_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_2_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_2_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_2_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_2_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_2_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_2_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_2_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_2_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_2_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_2_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_2_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_2_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_2_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_2_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_2_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_2_bits_executed;	// lsu.scala:210:16
  reg               ldq_2_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_2_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_2_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_2_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_2_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_2_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_3_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_3_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_3_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_3_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_3_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_3_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_3_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_3_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_3_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_3_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_3_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_3_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_3_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_3_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_3_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_3_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_3_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_3_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_3_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_3_bits_executed;	// lsu.scala:210:16
  reg               ldq_3_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_3_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_3_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_3_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_3_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_3_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_4_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_4_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_4_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_4_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_4_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_4_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_4_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_4_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_4_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_4_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_4_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_4_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_4_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_4_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_4_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_4_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_4_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_4_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_4_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_4_bits_executed;	// lsu.scala:210:16
  reg               ldq_4_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_4_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_4_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_4_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_4_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_4_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_5_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_5_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_5_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_5_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_5_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_5_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_5_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_5_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_5_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_5_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_5_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_5_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_5_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_5_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_5_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_5_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_5_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_5_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_5_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_5_bits_executed;	// lsu.scala:210:16
  reg               ldq_5_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_5_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_5_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_5_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_5_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_5_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_6_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_6_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_6_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_6_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_6_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_6_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_6_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_6_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_6_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_6_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_6_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_6_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_6_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_6_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_6_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_6_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_6_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_6_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_6_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_6_bits_executed;	// lsu.scala:210:16
  reg               ldq_6_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_6_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_6_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_6_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_6_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_6_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_7_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_7_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_7_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_7_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_7_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_7_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_7_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_7_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_7_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_7_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_7_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_7_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_7_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_7_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_7_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_7_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_7_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_7_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_7_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_7_bits_executed;	// lsu.scala:210:16
  reg               ldq_7_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_7_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_7_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_7_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_7_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_7_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_8_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_8_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_8_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_8_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_8_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_8_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_8_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_8_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_8_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_8_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_8_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_8_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_8_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_8_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_8_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_8_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_8_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_8_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_8_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_8_bits_executed;	// lsu.scala:210:16
  reg               ldq_8_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_8_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_8_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_8_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_8_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_8_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_9_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_9_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_9_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_9_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_9_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_9_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_9_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_9_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_9_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_9_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_9_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_9_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_9_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_9_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_9_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_9_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_9_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_9_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_9_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_9_bits_executed;	// lsu.scala:210:16
  reg               ldq_9_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_9_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_9_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_9_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_9_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_9_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_10_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_10_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_10_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_10_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_10_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_10_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_10_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_10_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_10_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_10_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_10_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_10_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_10_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_10_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_10_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_10_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_10_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_10_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_10_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_10_bits_executed;	// lsu.scala:210:16
  reg               ldq_10_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_10_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_10_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_10_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_10_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_10_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_11_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_11_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_11_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_11_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_11_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_11_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_11_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_11_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_11_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_11_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_11_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_11_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_11_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_11_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_11_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_11_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_11_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_11_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_11_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_11_bits_executed;	// lsu.scala:210:16
  reg               ldq_11_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_11_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_11_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_11_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_11_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_11_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_12_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_12_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_12_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_12_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_12_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_12_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_12_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_12_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_12_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_12_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_12_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_12_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_12_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_12_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_12_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_12_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_12_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_12_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_12_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_12_bits_executed;	// lsu.scala:210:16
  reg               ldq_12_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_12_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_12_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_12_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_12_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_12_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_13_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_13_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_13_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_13_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_13_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_13_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_13_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_13_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_13_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_13_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_13_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_13_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_13_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_13_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_13_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_13_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_13_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_13_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_13_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_13_bits_executed;	// lsu.scala:210:16
  reg               ldq_13_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_13_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_13_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_13_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_13_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_13_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_14_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_14_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_14_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_14_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_14_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_14_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_14_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_14_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_14_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_14_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_14_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_14_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_14_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_14_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_14_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_14_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_14_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_14_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_14_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_14_bits_executed;	// lsu.scala:210:16
  reg               ldq_14_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_14_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_14_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_14_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_14_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_14_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               ldq_15_valid;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_uopc;	// lsu.scala:210:16
  reg  [31:0]       ldq_15_bits_uop_inst;	// lsu.scala:210:16
  reg  [31:0]       ldq_15_bits_uop_debug_inst;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_rvc;	// lsu.scala:210:16
  reg  [39:0]       ldq_15_bits_uop_debug_pc;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_iq_type;	// lsu.scala:210:16
  reg  [9:0]        ldq_15_bits_uop_fu_code;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_ctrl_br_type;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_ctrl_op1_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_ctrl_op2_sel;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_ctrl_imm_sel;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_ctrl_op_fcn;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_fcn_dw;	// lsu.scala:210:16
  reg  [2:0]        ldq_15_bits_uop_ctrl_csr_cmd;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_is_load;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_is_sta;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ctrl_is_std;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_iw_state;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_iw_p1_poisoned;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_iw_p2_poisoned;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_br;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_jalr;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_jal;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_sfb;	// lsu.scala:210:16
  reg  [11:0]       ldq_15_bits_uop_br_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_br_tag;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_ftq_idx;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_edge_inst;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_pc_lob;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_taken;	// lsu.scala:210:16
  reg  [19:0]       ldq_15_bits_uop_imm_packed;	// lsu.scala:210:16
  reg  [11:0]       ldq_15_bits_uop_csr_addr;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_rob_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_ldq_idx;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_uop_stq_idx;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_rxq_idx;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_pdst;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_prs1;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_prs2;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_prs3;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_ppred;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_prs1_busy;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_prs2_busy;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_prs3_busy;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ppred_busy;	// lsu.scala:210:16
  reg  [6:0]        ldq_15_bits_uop_stale_pdst;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_exception;	// lsu.scala:210:16
  reg  [63:0]       ldq_15_bits_uop_exc_cause;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_bypassable;	// lsu.scala:210:16
  reg  [4:0]        ldq_15_bits_uop_mem_cmd;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_mem_size;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_mem_signed;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_fence;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_fencei;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_amo;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_uses_ldq;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_uses_stq;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_sys_pc2epc;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_is_unique;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_flush_on_commit;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ldst_is_rs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_ldst;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_lrs1;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_lrs2;	// lsu.scala:210:16
  reg  [5:0]        ldq_15_bits_uop_lrs3;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_ldst_val;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_dst_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_lrs1_rtype;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_lrs2_rtype;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_frs3_en;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_fp_val;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_fp_single;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_xcpt_pf_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_xcpt_ae_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_xcpt_ma_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_bp_debug_if;	// lsu.scala:210:16
  reg               ldq_15_bits_uop_bp_xcpt_if;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_debug_fsrc;	// lsu.scala:210:16
  reg  [1:0]        ldq_15_bits_uop_debug_tsrc;	// lsu.scala:210:16
  reg               ldq_15_bits_addr_valid;	// lsu.scala:210:16
  reg  [39:0]       ldq_15_bits_addr_bits;	// lsu.scala:210:16
  reg               ldq_15_bits_addr_is_virtual;	// lsu.scala:210:16
  reg               ldq_15_bits_addr_is_uncacheable;	// lsu.scala:210:16
  reg               ldq_15_bits_executed;	// lsu.scala:210:16
  reg               ldq_15_bits_succeeded;	// lsu.scala:210:16
  reg               ldq_15_bits_order_fail;	// lsu.scala:210:16
  reg               ldq_15_bits_observed;	// lsu.scala:210:16
  reg  [15:0]       ldq_15_bits_st_dep_mask;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_youngest_stq_idx;	// lsu.scala:210:16
  reg               ldq_15_bits_forward_std_val;	// lsu.scala:210:16
  reg  [3:0]        ldq_15_bits_forward_stq_idx;	// lsu.scala:210:16
  reg               stq_0_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_0_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_0_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_0_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_0_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_0_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_0_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_0_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_0_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_0_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_0_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_0_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_0_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_0_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_0_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_0_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_0_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_0_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_0_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_0_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_0_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_0_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_0_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_0_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_0_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_0_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_0_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_0_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_0_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_0_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_0_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_0_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_0_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_0_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_0_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_0_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_0_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_0_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_0_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_0_bits_data_bits;	// lsu.scala:211:16
  reg               stq_0_bits_committed;	// lsu.scala:211:16
  reg               stq_0_bits_succeeded;	// lsu.scala:211:16
  reg               stq_1_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_1_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_1_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_1_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_1_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_1_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_1_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_1_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_1_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_1_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_1_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_1_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_1_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_1_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_1_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_1_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_1_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_1_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_1_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_1_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_1_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_1_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_1_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_1_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_1_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_1_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_1_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_1_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_1_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_1_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_1_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_1_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_1_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_1_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_1_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_1_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_1_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_1_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_1_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_1_bits_data_bits;	// lsu.scala:211:16
  reg               stq_1_bits_committed;	// lsu.scala:211:16
  reg               stq_1_bits_succeeded;	// lsu.scala:211:16
  reg               stq_2_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_2_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_2_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_2_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_2_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_2_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_2_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_2_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_2_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_2_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_2_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_2_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_2_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_2_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_2_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_2_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_2_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_2_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_2_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_2_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_2_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_2_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_2_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_2_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_2_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_2_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_2_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_2_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_2_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_2_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_2_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_2_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_2_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_2_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_2_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_2_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_2_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_2_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_2_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_2_bits_data_bits;	// lsu.scala:211:16
  reg               stq_2_bits_committed;	// lsu.scala:211:16
  reg               stq_2_bits_succeeded;	// lsu.scala:211:16
  reg               stq_3_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_3_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_3_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_3_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_3_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_3_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_3_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_3_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_3_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_3_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_3_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_3_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_3_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_3_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_3_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_3_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_3_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_3_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_3_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_3_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_3_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_3_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_3_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_3_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_3_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_3_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_3_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_3_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_3_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_3_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_3_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_3_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_3_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_3_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_3_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_3_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_3_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_3_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_3_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_3_bits_data_bits;	// lsu.scala:211:16
  reg               stq_3_bits_committed;	// lsu.scala:211:16
  reg               stq_3_bits_succeeded;	// lsu.scala:211:16
  reg               stq_4_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_4_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_4_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_4_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_4_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_4_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_4_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_4_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_4_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_4_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_4_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_4_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_4_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_4_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_4_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_4_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_4_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_4_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_4_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_4_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_4_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_4_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_4_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_4_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_4_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_4_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_4_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_4_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_4_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_4_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_4_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_4_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_4_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_4_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_4_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_4_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_4_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_4_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_4_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_4_bits_data_bits;	// lsu.scala:211:16
  reg               stq_4_bits_committed;	// lsu.scala:211:16
  reg               stq_4_bits_succeeded;	// lsu.scala:211:16
  reg               stq_5_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_5_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_5_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_5_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_5_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_5_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_5_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_5_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_5_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_5_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_5_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_5_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_5_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_5_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_5_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_5_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_5_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_5_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_5_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_5_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_5_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_5_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_5_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_5_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_5_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_5_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_5_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_5_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_5_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_5_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_5_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_5_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_5_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_5_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_5_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_5_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_5_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_5_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_5_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_5_bits_data_bits;	// lsu.scala:211:16
  reg               stq_5_bits_committed;	// lsu.scala:211:16
  reg               stq_5_bits_succeeded;	// lsu.scala:211:16
  reg               stq_6_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_6_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_6_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_6_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_6_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_6_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_6_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_6_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_6_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_6_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_6_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_6_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_6_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_6_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_6_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_6_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_6_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_6_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_6_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_6_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_6_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_6_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_6_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_6_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_6_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_6_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_6_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_6_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_6_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_6_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_6_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_6_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_6_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_6_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_6_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_6_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_6_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_6_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_6_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_6_bits_data_bits;	// lsu.scala:211:16
  reg               stq_6_bits_committed;	// lsu.scala:211:16
  reg               stq_6_bits_succeeded;	// lsu.scala:211:16
  reg               stq_7_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_7_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_7_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_7_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_7_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_7_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_7_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_7_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_7_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_7_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_7_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_7_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_7_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_7_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_7_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_7_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_7_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_7_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_7_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_7_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_7_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_7_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_7_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_7_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_7_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_7_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_7_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_7_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_7_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_7_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_7_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_7_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_7_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_7_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_7_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_7_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_7_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_7_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_7_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_7_bits_data_bits;	// lsu.scala:211:16
  reg               stq_7_bits_committed;	// lsu.scala:211:16
  reg               stq_7_bits_succeeded;	// lsu.scala:211:16
  reg               stq_8_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_8_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_8_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_8_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_8_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_8_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_8_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_8_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_8_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_8_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_8_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_8_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_8_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_8_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_8_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_8_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_8_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_8_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_8_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_8_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_8_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_8_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_8_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_8_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_8_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_8_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_8_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_8_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_8_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_8_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_8_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_8_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_8_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_8_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_8_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_8_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_8_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_8_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_8_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_8_bits_data_bits;	// lsu.scala:211:16
  reg               stq_8_bits_committed;	// lsu.scala:211:16
  reg               stq_8_bits_succeeded;	// lsu.scala:211:16
  reg               stq_9_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_9_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_9_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_9_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_9_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_9_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_9_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_9_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_9_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_9_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_9_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_9_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_9_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_9_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_9_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_9_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_9_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_9_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_9_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_9_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_9_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_9_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_9_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_9_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_9_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_9_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_9_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_9_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_9_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_9_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_9_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_9_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_9_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_9_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_9_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_9_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_9_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_9_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_9_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_9_bits_data_bits;	// lsu.scala:211:16
  reg               stq_9_bits_committed;	// lsu.scala:211:16
  reg               stq_9_bits_succeeded;	// lsu.scala:211:16
  reg               stq_10_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_10_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_10_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_10_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_10_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_10_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_10_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_10_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_10_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_10_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_10_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_10_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_10_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_10_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_10_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_10_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_10_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_10_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_10_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_10_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_10_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_10_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_10_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_10_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_10_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_10_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_10_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_10_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_10_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_10_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_10_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_10_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_10_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_10_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_10_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_10_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_10_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_10_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_10_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_10_bits_data_bits;	// lsu.scala:211:16
  reg               stq_10_bits_committed;	// lsu.scala:211:16
  reg               stq_10_bits_succeeded;	// lsu.scala:211:16
  reg               stq_11_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_11_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_11_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_11_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_11_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_11_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_11_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_11_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_11_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_11_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_11_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_11_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_11_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_11_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_11_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_11_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_11_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_11_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_11_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_11_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_11_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_11_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_11_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_11_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_11_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_11_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_11_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_11_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_11_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_11_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_11_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_11_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_11_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_11_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_11_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_11_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_11_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_11_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_11_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_11_bits_data_bits;	// lsu.scala:211:16
  reg               stq_11_bits_committed;	// lsu.scala:211:16
  reg               stq_11_bits_succeeded;	// lsu.scala:211:16
  reg               stq_12_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_12_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_12_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_12_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_12_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_12_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_12_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_12_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_12_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_12_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_12_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_12_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_12_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_12_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_12_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_12_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_12_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_12_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_12_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_12_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_12_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_12_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_12_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_12_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_12_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_12_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_12_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_12_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_12_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_12_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_12_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_12_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_12_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_12_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_12_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_12_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_12_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_12_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_12_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_12_bits_data_bits;	// lsu.scala:211:16
  reg               stq_12_bits_committed;	// lsu.scala:211:16
  reg               stq_12_bits_succeeded;	// lsu.scala:211:16
  reg               stq_13_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_13_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_13_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_13_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_13_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_13_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_13_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_13_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_13_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_13_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_13_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_13_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_13_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_13_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_13_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_13_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_13_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_13_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_13_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_13_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_13_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_13_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_13_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_13_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_13_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_13_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_13_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_13_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_13_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_13_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_13_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_13_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_13_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_13_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_13_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_13_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_13_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_13_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_13_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_13_bits_data_bits;	// lsu.scala:211:16
  reg               stq_13_bits_committed;	// lsu.scala:211:16
  reg               stq_13_bits_succeeded;	// lsu.scala:211:16
  reg               stq_14_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_14_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_14_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_14_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_14_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_14_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_14_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_14_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_14_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_14_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_14_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_14_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_14_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_14_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_14_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_14_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_14_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_14_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_14_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_14_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_14_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_14_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_14_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_14_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_14_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_14_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_14_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_14_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_14_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_14_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_14_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_14_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_14_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_14_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_14_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_14_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_14_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_14_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_14_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_14_bits_data_bits;	// lsu.scala:211:16
  reg               stq_14_bits_committed;	// lsu.scala:211:16
  reg               stq_14_bits_succeeded;	// lsu.scala:211:16
  reg               stq_15_valid;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_uopc;	// lsu.scala:211:16
  reg  [31:0]       stq_15_bits_uop_inst;	// lsu.scala:211:16
  reg  [31:0]       stq_15_bits_uop_debug_inst;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_rvc;	// lsu.scala:211:16
  reg  [39:0]       stq_15_bits_uop_debug_pc;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_iq_type;	// lsu.scala:211:16
  reg  [9:0]        stq_15_bits_uop_fu_code;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_ctrl_br_type;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_ctrl_op1_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_ctrl_op2_sel;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_ctrl_imm_sel;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_ctrl_op_fcn;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_fcn_dw;	// lsu.scala:211:16
  reg  [2:0]        stq_15_bits_uop_ctrl_csr_cmd;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_is_load;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_is_sta;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ctrl_is_std;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_iw_state;	// lsu.scala:211:16
  reg               stq_15_bits_uop_iw_p1_poisoned;	// lsu.scala:211:16
  reg               stq_15_bits_uop_iw_p2_poisoned;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_br;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_jalr;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_jal;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_sfb;	// lsu.scala:211:16
  reg  [11:0]       stq_15_bits_uop_br_mask;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_br_tag;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_ftq_idx;	// lsu.scala:211:16
  reg               stq_15_bits_uop_edge_inst;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_pc_lob;	// lsu.scala:211:16
  reg               stq_15_bits_uop_taken;	// lsu.scala:211:16
  reg  [19:0]       stq_15_bits_uop_imm_packed;	// lsu.scala:211:16
  reg  [11:0]       stq_15_bits_uop_csr_addr;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_rob_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_ldq_idx;	// lsu.scala:211:16
  reg  [3:0]        stq_15_bits_uop_stq_idx;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_rxq_idx;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_pdst;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_prs1;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_prs2;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_prs3;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_ppred;	// lsu.scala:211:16
  reg               stq_15_bits_uop_prs1_busy;	// lsu.scala:211:16
  reg               stq_15_bits_uop_prs2_busy;	// lsu.scala:211:16
  reg               stq_15_bits_uop_prs3_busy;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ppred_busy;	// lsu.scala:211:16
  reg  [6:0]        stq_15_bits_uop_stale_pdst;	// lsu.scala:211:16
  reg               stq_15_bits_uop_exception;	// lsu.scala:211:16
  reg  [63:0]       stq_15_bits_uop_exc_cause;	// lsu.scala:211:16
  reg               stq_15_bits_uop_bypassable;	// lsu.scala:211:16
  reg  [4:0]        stq_15_bits_uop_mem_cmd;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_mem_size;	// lsu.scala:211:16
  reg               stq_15_bits_uop_mem_signed;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_fence;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_fencei;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_amo;	// lsu.scala:211:16
  reg               stq_15_bits_uop_uses_ldq;	// lsu.scala:211:16
  reg               stq_15_bits_uop_uses_stq;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_sys_pc2epc;	// lsu.scala:211:16
  reg               stq_15_bits_uop_is_unique;	// lsu.scala:211:16
  reg               stq_15_bits_uop_flush_on_commit;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ldst_is_rs1;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_ldst;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_lrs1;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_lrs2;	// lsu.scala:211:16
  reg  [5:0]        stq_15_bits_uop_lrs3;	// lsu.scala:211:16
  reg               stq_15_bits_uop_ldst_val;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_dst_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_lrs1_rtype;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_lrs2_rtype;	// lsu.scala:211:16
  reg               stq_15_bits_uop_frs3_en;	// lsu.scala:211:16
  reg               stq_15_bits_uop_fp_val;	// lsu.scala:211:16
  reg               stq_15_bits_uop_fp_single;	// lsu.scala:211:16
  reg               stq_15_bits_uop_xcpt_pf_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_xcpt_ae_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_xcpt_ma_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_bp_debug_if;	// lsu.scala:211:16
  reg               stq_15_bits_uop_bp_xcpt_if;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_debug_fsrc;	// lsu.scala:211:16
  reg  [1:0]        stq_15_bits_uop_debug_tsrc;	// lsu.scala:211:16
  reg               stq_15_bits_addr_valid;	// lsu.scala:211:16
  reg  [39:0]       stq_15_bits_addr_bits;	// lsu.scala:211:16
  reg               stq_15_bits_addr_is_virtual;	// lsu.scala:211:16
  reg               stq_15_bits_data_valid;	// lsu.scala:211:16
  reg  [63:0]       stq_15_bits_data_bits;	// lsu.scala:211:16
  reg               stq_15_bits_committed;	// lsu.scala:211:16
  reg               stq_15_bits_succeeded;	// lsu.scala:211:16
  reg  [3:0]        ldq_head;	// lsu.scala:215:29
  reg  [3:0]        ldq_tail;	// lsu.scala:216:29
  reg  [3:0]        stq_head;	// lsu.scala:217:29
  reg  [3:0]        stq_tail;	// lsu.scala:218:29
  reg  [3:0]        stq_commit_head;	// lsu.scala:219:29
  reg  [3:0]        stq_execute_head;	// lsu.scala:220:29
  wire [15:0]       _GEN_2 =
    {{stq_15_valid},
     {stq_14_valid},
     {stq_13_valid},
     {stq_12_valid},
     {stq_11_valid},
     {stq_10_valid},
     {stq_9_valid},
     {stq_8_valid},
     {stq_7_valid},
     {stq_6_valid},
     {stq_5_valid},
     {stq_4_valid},
     {stq_3_valid},
     {stq_2_valid},
     {stq_1_valid},
     {stq_0_valid}};	// lsu.scala:211:16, :224:42
  wire              _GEN_3 = _GEN_2[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [15:0][6:0]  _GEN_4 =
    {{stq_15_bits_uop_uopc},
     {stq_14_bits_uop_uopc},
     {stq_13_bits_uop_uopc},
     {stq_12_bits_uop_uopc},
     {stq_11_bits_uop_uopc},
     {stq_10_bits_uop_uopc},
     {stq_9_bits_uop_uopc},
     {stq_8_bits_uop_uopc},
     {stq_7_bits_uop_uopc},
     {stq_6_bits_uop_uopc},
     {stq_5_bits_uop_uopc},
     {stq_4_bits_uop_uopc},
     {stq_3_bits_uop_uopc},
     {stq_2_bits_uop_uopc},
     {stq_1_bits_uop_uopc},
     {stq_0_bits_uop_uopc}};	// lsu.scala:211:16, :224:42
  wire [15:0][31:0] _GEN_5 =
    {{stq_15_bits_uop_inst},
     {stq_14_bits_uop_inst},
     {stq_13_bits_uop_inst},
     {stq_12_bits_uop_inst},
     {stq_11_bits_uop_inst},
     {stq_10_bits_uop_inst},
     {stq_9_bits_uop_inst},
     {stq_8_bits_uop_inst},
     {stq_7_bits_uop_inst},
     {stq_6_bits_uop_inst},
     {stq_5_bits_uop_inst},
     {stq_4_bits_uop_inst},
     {stq_3_bits_uop_inst},
     {stq_2_bits_uop_inst},
     {stq_1_bits_uop_inst},
     {stq_0_bits_uop_inst}};	// lsu.scala:211:16, :224:42
  wire [15:0][31:0] _GEN_6 =
    {{stq_15_bits_uop_debug_inst},
     {stq_14_bits_uop_debug_inst},
     {stq_13_bits_uop_debug_inst},
     {stq_12_bits_uop_debug_inst},
     {stq_11_bits_uop_debug_inst},
     {stq_10_bits_uop_debug_inst},
     {stq_9_bits_uop_debug_inst},
     {stq_8_bits_uop_debug_inst},
     {stq_7_bits_uop_debug_inst},
     {stq_6_bits_uop_debug_inst},
     {stq_5_bits_uop_debug_inst},
     {stq_4_bits_uop_debug_inst},
     {stq_3_bits_uop_debug_inst},
     {stq_2_bits_uop_debug_inst},
     {stq_1_bits_uop_debug_inst},
     {stq_0_bits_uop_debug_inst}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_7 =
    {{stq_15_bits_uop_is_rvc},
     {stq_14_bits_uop_is_rvc},
     {stq_13_bits_uop_is_rvc},
     {stq_12_bits_uop_is_rvc},
     {stq_11_bits_uop_is_rvc},
     {stq_10_bits_uop_is_rvc},
     {stq_9_bits_uop_is_rvc},
     {stq_8_bits_uop_is_rvc},
     {stq_7_bits_uop_is_rvc},
     {stq_6_bits_uop_is_rvc},
     {stq_5_bits_uop_is_rvc},
     {stq_4_bits_uop_is_rvc},
     {stq_3_bits_uop_is_rvc},
     {stq_2_bits_uop_is_rvc},
     {stq_1_bits_uop_is_rvc},
     {stq_0_bits_uop_is_rvc}};	// lsu.scala:211:16, :224:42
  wire [15:0][39:0] _GEN_8 =
    {{stq_15_bits_uop_debug_pc},
     {stq_14_bits_uop_debug_pc},
     {stq_13_bits_uop_debug_pc},
     {stq_12_bits_uop_debug_pc},
     {stq_11_bits_uop_debug_pc},
     {stq_10_bits_uop_debug_pc},
     {stq_9_bits_uop_debug_pc},
     {stq_8_bits_uop_debug_pc},
     {stq_7_bits_uop_debug_pc},
     {stq_6_bits_uop_debug_pc},
     {stq_5_bits_uop_debug_pc},
     {stq_4_bits_uop_debug_pc},
     {stq_3_bits_uop_debug_pc},
     {stq_2_bits_uop_debug_pc},
     {stq_1_bits_uop_debug_pc},
     {stq_0_bits_uop_debug_pc}};	// lsu.scala:211:16, :224:42
  wire [15:0][2:0]  _GEN_9 =
    {{stq_15_bits_uop_iq_type},
     {stq_14_bits_uop_iq_type},
     {stq_13_bits_uop_iq_type},
     {stq_12_bits_uop_iq_type},
     {stq_11_bits_uop_iq_type},
     {stq_10_bits_uop_iq_type},
     {stq_9_bits_uop_iq_type},
     {stq_8_bits_uop_iq_type},
     {stq_7_bits_uop_iq_type},
     {stq_6_bits_uop_iq_type},
     {stq_5_bits_uop_iq_type},
     {stq_4_bits_uop_iq_type},
     {stq_3_bits_uop_iq_type},
     {stq_2_bits_uop_iq_type},
     {stq_1_bits_uop_iq_type},
     {stq_0_bits_uop_iq_type}};	// lsu.scala:211:16, :224:42
  wire [15:0][9:0]  _GEN_10 =
    {{stq_15_bits_uop_fu_code},
     {stq_14_bits_uop_fu_code},
     {stq_13_bits_uop_fu_code},
     {stq_12_bits_uop_fu_code},
     {stq_11_bits_uop_fu_code},
     {stq_10_bits_uop_fu_code},
     {stq_9_bits_uop_fu_code},
     {stq_8_bits_uop_fu_code},
     {stq_7_bits_uop_fu_code},
     {stq_6_bits_uop_fu_code},
     {stq_5_bits_uop_fu_code},
     {stq_4_bits_uop_fu_code},
     {stq_3_bits_uop_fu_code},
     {stq_2_bits_uop_fu_code},
     {stq_1_bits_uop_fu_code},
     {stq_0_bits_uop_fu_code}};	// lsu.scala:211:16, :224:42
  wire [15:0][3:0]  _GEN_11 =
    {{stq_15_bits_uop_ctrl_br_type},
     {stq_14_bits_uop_ctrl_br_type},
     {stq_13_bits_uop_ctrl_br_type},
     {stq_12_bits_uop_ctrl_br_type},
     {stq_11_bits_uop_ctrl_br_type},
     {stq_10_bits_uop_ctrl_br_type},
     {stq_9_bits_uop_ctrl_br_type},
     {stq_8_bits_uop_ctrl_br_type},
     {stq_7_bits_uop_ctrl_br_type},
     {stq_6_bits_uop_ctrl_br_type},
     {stq_5_bits_uop_ctrl_br_type},
     {stq_4_bits_uop_ctrl_br_type},
     {stq_3_bits_uop_ctrl_br_type},
     {stq_2_bits_uop_ctrl_br_type},
     {stq_1_bits_uop_ctrl_br_type},
     {stq_0_bits_uop_ctrl_br_type}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_12 =
    {{stq_15_bits_uop_ctrl_op1_sel},
     {stq_14_bits_uop_ctrl_op1_sel},
     {stq_13_bits_uop_ctrl_op1_sel},
     {stq_12_bits_uop_ctrl_op1_sel},
     {stq_11_bits_uop_ctrl_op1_sel},
     {stq_10_bits_uop_ctrl_op1_sel},
     {stq_9_bits_uop_ctrl_op1_sel},
     {stq_8_bits_uop_ctrl_op1_sel},
     {stq_7_bits_uop_ctrl_op1_sel},
     {stq_6_bits_uop_ctrl_op1_sel},
     {stq_5_bits_uop_ctrl_op1_sel},
     {stq_4_bits_uop_ctrl_op1_sel},
     {stq_3_bits_uop_ctrl_op1_sel},
     {stq_2_bits_uop_ctrl_op1_sel},
     {stq_1_bits_uop_ctrl_op1_sel},
     {stq_0_bits_uop_ctrl_op1_sel}};	// lsu.scala:211:16, :224:42
  wire [15:0][2:0]  _GEN_13 =
    {{stq_15_bits_uop_ctrl_op2_sel},
     {stq_14_bits_uop_ctrl_op2_sel},
     {stq_13_bits_uop_ctrl_op2_sel},
     {stq_12_bits_uop_ctrl_op2_sel},
     {stq_11_bits_uop_ctrl_op2_sel},
     {stq_10_bits_uop_ctrl_op2_sel},
     {stq_9_bits_uop_ctrl_op2_sel},
     {stq_8_bits_uop_ctrl_op2_sel},
     {stq_7_bits_uop_ctrl_op2_sel},
     {stq_6_bits_uop_ctrl_op2_sel},
     {stq_5_bits_uop_ctrl_op2_sel},
     {stq_4_bits_uop_ctrl_op2_sel},
     {stq_3_bits_uop_ctrl_op2_sel},
     {stq_2_bits_uop_ctrl_op2_sel},
     {stq_1_bits_uop_ctrl_op2_sel},
     {stq_0_bits_uop_ctrl_op2_sel}};	// lsu.scala:211:16, :224:42
  wire [15:0][2:0]  _GEN_14 =
    {{stq_15_bits_uop_ctrl_imm_sel},
     {stq_14_bits_uop_ctrl_imm_sel},
     {stq_13_bits_uop_ctrl_imm_sel},
     {stq_12_bits_uop_ctrl_imm_sel},
     {stq_11_bits_uop_ctrl_imm_sel},
     {stq_10_bits_uop_ctrl_imm_sel},
     {stq_9_bits_uop_ctrl_imm_sel},
     {stq_8_bits_uop_ctrl_imm_sel},
     {stq_7_bits_uop_ctrl_imm_sel},
     {stq_6_bits_uop_ctrl_imm_sel},
     {stq_5_bits_uop_ctrl_imm_sel},
     {stq_4_bits_uop_ctrl_imm_sel},
     {stq_3_bits_uop_ctrl_imm_sel},
     {stq_2_bits_uop_ctrl_imm_sel},
     {stq_1_bits_uop_ctrl_imm_sel},
     {stq_0_bits_uop_ctrl_imm_sel}};	// lsu.scala:211:16, :224:42
  wire [15:0][3:0]  _GEN_15 =
    {{stq_15_bits_uop_ctrl_op_fcn},
     {stq_14_bits_uop_ctrl_op_fcn},
     {stq_13_bits_uop_ctrl_op_fcn},
     {stq_12_bits_uop_ctrl_op_fcn},
     {stq_11_bits_uop_ctrl_op_fcn},
     {stq_10_bits_uop_ctrl_op_fcn},
     {stq_9_bits_uop_ctrl_op_fcn},
     {stq_8_bits_uop_ctrl_op_fcn},
     {stq_7_bits_uop_ctrl_op_fcn},
     {stq_6_bits_uop_ctrl_op_fcn},
     {stq_5_bits_uop_ctrl_op_fcn},
     {stq_4_bits_uop_ctrl_op_fcn},
     {stq_3_bits_uop_ctrl_op_fcn},
     {stq_2_bits_uop_ctrl_op_fcn},
     {stq_1_bits_uop_ctrl_op_fcn},
     {stq_0_bits_uop_ctrl_op_fcn}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_16 =
    {{stq_15_bits_uop_ctrl_fcn_dw},
     {stq_14_bits_uop_ctrl_fcn_dw},
     {stq_13_bits_uop_ctrl_fcn_dw},
     {stq_12_bits_uop_ctrl_fcn_dw},
     {stq_11_bits_uop_ctrl_fcn_dw},
     {stq_10_bits_uop_ctrl_fcn_dw},
     {stq_9_bits_uop_ctrl_fcn_dw},
     {stq_8_bits_uop_ctrl_fcn_dw},
     {stq_7_bits_uop_ctrl_fcn_dw},
     {stq_6_bits_uop_ctrl_fcn_dw},
     {stq_5_bits_uop_ctrl_fcn_dw},
     {stq_4_bits_uop_ctrl_fcn_dw},
     {stq_3_bits_uop_ctrl_fcn_dw},
     {stq_2_bits_uop_ctrl_fcn_dw},
     {stq_1_bits_uop_ctrl_fcn_dw},
     {stq_0_bits_uop_ctrl_fcn_dw}};	// lsu.scala:211:16, :224:42
  wire [15:0][2:0]  _GEN_17 =
    {{stq_15_bits_uop_ctrl_csr_cmd},
     {stq_14_bits_uop_ctrl_csr_cmd},
     {stq_13_bits_uop_ctrl_csr_cmd},
     {stq_12_bits_uop_ctrl_csr_cmd},
     {stq_11_bits_uop_ctrl_csr_cmd},
     {stq_10_bits_uop_ctrl_csr_cmd},
     {stq_9_bits_uop_ctrl_csr_cmd},
     {stq_8_bits_uop_ctrl_csr_cmd},
     {stq_7_bits_uop_ctrl_csr_cmd},
     {stq_6_bits_uop_ctrl_csr_cmd},
     {stq_5_bits_uop_ctrl_csr_cmd},
     {stq_4_bits_uop_ctrl_csr_cmd},
     {stq_3_bits_uop_ctrl_csr_cmd},
     {stq_2_bits_uop_ctrl_csr_cmd},
     {stq_1_bits_uop_ctrl_csr_cmd},
     {stq_0_bits_uop_ctrl_csr_cmd}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_18 =
    {{stq_15_bits_uop_ctrl_is_load},
     {stq_14_bits_uop_ctrl_is_load},
     {stq_13_bits_uop_ctrl_is_load},
     {stq_12_bits_uop_ctrl_is_load},
     {stq_11_bits_uop_ctrl_is_load},
     {stq_10_bits_uop_ctrl_is_load},
     {stq_9_bits_uop_ctrl_is_load},
     {stq_8_bits_uop_ctrl_is_load},
     {stq_7_bits_uop_ctrl_is_load},
     {stq_6_bits_uop_ctrl_is_load},
     {stq_5_bits_uop_ctrl_is_load},
     {stq_4_bits_uop_ctrl_is_load},
     {stq_3_bits_uop_ctrl_is_load},
     {stq_2_bits_uop_ctrl_is_load},
     {stq_1_bits_uop_ctrl_is_load},
     {stq_0_bits_uop_ctrl_is_load}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_19 =
    {{stq_15_bits_uop_ctrl_is_sta},
     {stq_14_bits_uop_ctrl_is_sta},
     {stq_13_bits_uop_ctrl_is_sta},
     {stq_12_bits_uop_ctrl_is_sta},
     {stq_11_bits_uop_ctrl_is_sta},
     {stq_10_bits_uop_ctrl_is_sta},
     {stq_9_bits_uop_ctrl_is_sta},
     {stq_8_bits_uop_ctrl_is_sta},
     {stq_7_bits_uop_ctrl_is_sta},
     {stq_6_bits_uop_ctrl_is_sta},
     {stq_5_bits_uop_ctrl_is_sta},
     {stq_4_bits_uop_ctrl_is_sta},
     {stq_3_bits_uop_ctrl_is_sta},
     {stq_2_bits_uop_ctrl_is_sta},
     {stq_1_bits_uop_ctrl_is_sta},
     {stq_0_bits_uop_ctrl_is_sta}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_20 =
    {{stq_15_bits_uop_ctrl_is_std},
     {stq_14_bits_uop_ctrl_is_std},
     {stq_13_bits_uop_ctrl_is_std},
     {stq_12_bits_uop_ctrl_is_std},
     {stq_11_bits_uop_ctrl_is_std},
     {stq_10_bits_uop_ctrl_is_std},
     {stq_9_bits_uop_ctrl_is_std},
     {stq_8_bits_uop_ctrl_is_std},
     {stq_7_bits_uop_ctrl_is_std},
     {stq_6_bits_uop_ctrl_is_std},
     {stq_5_bits_uop_ctrl_is_std},
     {stq_4_bits_uop_ctrl_is_std},
     {stq_3_bits_uop_ctrl_is_std},
     {stq_2_bits_uop_ctrl_is_std},
     {stq_1_bits_uop_ctrl_is_std},
     {stq_0_bits_uop_ctrl_is_std}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_21 =
    {{stq_15_bits_uop_iw_state},
     {stq_14_bits_uop_iw_state},
     {stq_13_bits_uop_iw_state},
     {stq_12_bits_uop_iw_state},
     {stq_11_bits_uop_iw_state},
     {stq_10_bits_uop_iw_state},
     {stq_9_bits_uop_iw_state},
     {stq_8_bits_uop_iw_state},
     {stq_7_bits_uop_iw_state},
     {stq_6_bits_uop_iw_state},
     {stq_5_bits_uop_iw_state},
     {stq_4_bits_uop_iw_state},
     {stq_3_bits_uop_iw_state},
     {stq_2_bits_uop_iw_state},
     {stq_1_bits_uop_iw_state},
     {stq_0_bits_uop_iw_state}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_22 =
    {{stq_15_bits_uop_iw_p1_poisoned},
     {stq_14_bits_uop_iw_p1_poisoned},
     {stq_13_bits_uop_iw_p1_poisoned},
     {stq_12_bits_uop_iw_p1_poisoned},
     {stq_11_bits_uop_iw_p1_poisoned},
     {stq_10_bits_uop_iw_p1_poisoned},
     {stq_9_bits_uop_iw_p1_poisoned},
     {stq_8_bits_uop_iw_p1_poisoned},
     {stq_7_bits_uop_iw_p1_poisoned},
     {stq_6_bits_uop_iw_p1_poisoned},
     {stq_5_bits_uop_iw_p1_poisoned},
     {stq_4_bits_uop_iw_p1_poisoned},
     {stq_3_bits_uop_iw_p1_poisoned},
     {stq_2_bits_uop_iw_p1_poisoned},
     {stq_1_bits_uop_iw_p1_poisoned},
     {stq_0_bits_uop_iw_p1_poisoned}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_23 =
    {{stq_15_bits_uop_iw_p2_poisoned},
     {stq_14_bits_uop_iw_p2_poisoned},
     {stq_13_bits_uop_iw_p2_poisoned},
     {stq_12_bits_uop_iw_p2_poisoned},
     {stq_11_bits_uop_iw_p2_poisoned},
     {stq_10_bits_uop_iw_p2_poisoned},
     {stq_9_bits_uop_iw_p2_poisoned},
     {stq_8_bits_uop_iw_p2_poisoned},
     {stq_7_bits_uop_iw_p2_poisoned},
     {stq_6_bits_uop_iw_p2_poisoned},
     {stq_5_bits_uop_iw_p2_poisoned},
     {stq_4_bits_uop_iw_p2_poisoned},
     {stq_3_bits_uop_iw_p2_poisoned},
     {stq_2_bits_uop_iw_p2_poisoned},
     {stq_1_bits_uop_iw_p2_poisoned},
     {stq_0_bits_uop_iw_p2_poisoned}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_24 =
    {{stq_15_bits_uop_is_br},
     {stq_14_bits_uop_is_br},
     {stq_13_bits_uop_is_br},
     {stq_12_bits_uop_is_br},
     {stq_11_bits_uop_is_br},
     {stq_10_bits_uop_is_br},
     {stq_9_bits_uop_is_br},
     {stq_8_bits_uop_is_br},
     {stq_7_bits_uop_is_br},
     {stq_6_bits_uop_is_br},
     {stq_5_bits_uop_is_br},
     {stq_4_bits_uop_is_br},
     {stq_3_bits_uop_is_br},
     {stq_2_bits_uop_is_br},
     {stq_1_bits_uop_is_br},
     {stq_0_bits_uop_is_br}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_25 =
    {{stq_15_bits_uop_is_jalr},
     {stq_14_bits_uop_is_jalr},
     {stq_13_bits_uop_is_jalr},
     {stq_12_bits_uop_is_jalr},
     {stq_11_bits_uop_is_jalr},
     {stq_10_bits_uop_is_jalr},
     {stq_9_bits_uop_is_jalr},
     {stq_8_bits_uop_is_jalr},
     {stq_7_bits_uop_is_jalr},
     {stq_6_bits_uop_is_jalr},
     {stq_5_bits_uop_is_jalr},
     {stq_4_bits_uop_is_jalr},
     {stq_3_bits_uop_is_jalr},
     {stq_2_bits_uop_is_jalr},
     {stq_1_bits_uop_is_jalr},
     {stq_0_bits_uop_is_jalr}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_26 =
    {{stq_15_bits_uop_is_jal},
     {stq_14_bits_uop_is_jal},
     {stq_13_bits_uop_is_jal},
     {stq_12_bits_uop_is_jal},
     {stq_11_bits_uop_is_jal},
     {stq_10_bits_uop_is_jal},
     {stq_9_bits_uop_is_jal},
     {stq_8_bits_uop_is_jal},
     {stq_7_bits_uop_is_jal},
     {stq_6_bits_uop_is_jal},
     {stq_5_bits_uop_is_jal},
     {stq_4_bits_uop_is_jal},
     {stq_3_bits_uop_is_jal},
     {stq_2_bits_uop_is_jal},
     {stq_1_bits_uop_is_jal},
     {stq_0_bits_uop_is_jal}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_27 =
    {{stq_15_bits_uop_is_sfb},
     {stq_14_bits_uop_is_sfb},
     {stq_13_bits_uop_is_sfb},
     {stq_12_bits_uop_is_sfb},
     {stq_11_bits_uop_is_sfb},
     {stq_10_bits_uop_is_sfb},
     {stq_9_bits_uop_is_sfb},
     {stq_8_bits_uop_is_sfb},
     {stq_7_bits_uop_is_sfb},
     {stq_6_bits_uop_is_sfb},
     {stq_5_bits_uop_is_sfb},
     {stq_4_bits_uop_is_sfb},
     {stq_3_bits_uop_is_sfb},
     {stq_2_bits_uop_is_sfb},
     {stq_1_bits_uop_is_sfb},
     {stq_0_bits_uop_is_sfb}};	// lsu.scala:211:16, :224:42
  wire [15:0][11:0] _GEN_28 =
    {{stq_15_bits_uop_br_mask},
     {stq_14_bits_uop_br_mask},
     {stq_13_bits_uop_br_mask},
     {stq_12_bits_uop_br_mask},
     {stq_11_bits_uop_br_mask},
     {stq_10_bits_uop_br_mask},
     {stq_9_bits_uop_br_mask},
     {stq_8_bits_uop_br_mask},
     {stq_7_bits_uop_br_mask},
     {stq_6_bits_uop_br_mask},
     {stq_5_bits_uop_br_mask},
     {stq_4_bits_uop_br_mask},
     {stq_3_bits_uop_br_mask},
     {stq_2_bits_uop_br_mask},
     {stq_1_bits_uop_br_mask},
     {stq_0_bits_uop_br_mask}};	// lsu.scala:211:16, :224:42
  wire [15:0][3:0]  _GEN_29 =
    {{stq_15_bits_uop_br_tag},
     {stq_14_bits_uop_br_tag},
     {stq_13_bits_uop_br_tag},
     {stq_12_bits_uop_br_tag},
     {stq_11_bits_uop_br_tag},
     {stq_10_bits_uop_br_tag},
     {stq_9_bits_uop_br_tag},
     {stq_8_bits_uop_br_tag},
     {stq_7_bits_uop_br_tag},
     {stq_6_bits_uop_br_tag},
     {stq_5_bits_uop_br_tag},
     {stq_4_bits_uop_br_tag},
     {stq_3_bits_uop_br_tag},
     {stq_2_bits_uop_br_tag},
     {stq_1_bits_uop_br_tag},
     {stq_0_bits_uop_br_tag}};	// lsu.scala:211:16, :224:42
  wire [15:0][4:0]  _GEN_30 =
    {{stq_15_bits_uop_ftq_idx},
     {stq_14_bits_uop_ftq_idx},
     {stq_13_bits_uop_ftq_idx},
     {stq_12_bits_uop_ftq_idx},
     {stq_11_bits_uop_ftq_idx},
     {stq_10_bits_uop_ftq_idx},
     {stq_9_bits_uop_ftq_idx},
     {stq_8_bits_uop_ftq_idx},
     {stq_7_bits_uop_ftq_idx},
     {stq_6_bits_uop_ftq_idx},
     {stq_5_bits_uop_ftq_idx},
     {stq_4_bits_uop_ftq_idx},
     {stq_3_bits_uop_ftq_idx},
     {stq_2_bits_uop_ftq_idx},
     {stq_1_bits_uop_ftq_idx},
     {stq_0_bits_uop_ftq_idx}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_31 =
    {{stq_15_bits_uop_edge_inst},
     {stq_14_bits_uop_edge_inst},
     {stq_13_bits_uop_edge_inst},
     {stq_12_bits_uop_edge_inst},
     {stq_11_bits_uop_edge_inst},
     {stq_10_bits_uop_edge_inst},
     {stq_9_bits_uop_edge_inst},
     {stq_8_bits_uop_edge_inst},
     {stq_7_bits_uop_edge_inst},
     {stq_6_bits_uop_edge_inst},
     {stq_5_bits_uop_edge_inst},
     {stq_4_bits_uop_edge_inst},
     {stq_3_bits_uop_edge_inst},
     {stq_2_bits_uop_edge_inst},
     {stq_1_bits_uop_edge_inst},
     {stq_0_bits_uop_edge_inst}};	// lsu.scala:211:16, :224:42
  wire [15:0][5:0]  _GEN_32 =
    {{stq_15_bits_uop_pc_lob},
     {stq_14_bits_uop_pc_lob},
     {stq_13_bits_uop_pc_lob},
     {stq_12_bits_uop_pc_lob},
     {stq_11_bits_uop_pc_lob},
     {stq_10_bits_uop_pc_lob},
     {stq_9_bits_uop_pc_lob},
     {stq_8_bits_uop_pc_lob},
     {stq_7_bits_uop_pc_lob},
     {stq_6_bits_uop_pc_lob},
     {stq_5_bits_uop_pc_lob},
     {stq_4_bits_uop_pc_lob},
     {stq_3_bits_uop_pc_lob},
     {stq_2_bits_uop_pc_lob},
     {stq_1_bits_uop_pc_lob},
     {stq_0_bits_uop_pc_lob}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_33 =
    {{stq_15_bits_uop_taken},
     {stq_14_bits_uop_taken},
     {stq_13_bits_uop_taken},
     {stq_12_bits_uop_taken},
     {stq_11_bits_uop_taken},
     {stq_10_bits_uop_taken},
     {stq_9_bits_uop_taken},
     {stq_8_bits_uop_taken},
     {stq_7_bits_uop_taken},
     {stq_6_bits_uop_taken},
     {stq_5_bits_uop_taken},
     {stq_4_bits_uop_taken},
     {stq_3_bits_uop_taken},
     {stq_2_bits_uop_taken},
     {stq_1_bits_uop_taken},
     {stq_0_bits_uop_taken}};	// lsu.scala:211:16, :224:42
  wire [15:0][19:0] _GEN_34 =
    {{stq_15_bits_uop_imm_packed},
     {stq_14_bits_uop_imm_packed},
     {stq_13_bits_uop_imm_packed},
     {stq_12_bits_uop_imm_packed},
     {stq_11_bits_uop_imm_packed},
     {stq_10_bits_uop_imm_packed},
     {stq_9_bits_uop_imm_packed},
     {stq_8_bits_uop_imm_packed},
     {stq_7_bits_uop_imm_packed},
     {stq_6_bits_uop_imm_packed},
     {stq_5_bits_uop_imm_packed},
     {stq_4_bits_uop_imm_packed},
     {stq_3_bits_uop_imm_packed},
     {stq_2_bits_uop_imm_packed},
     {stq_1_bits_uop_imm_packed},
     {stq_0_bits_uop_imm_packed}};	// lsu.scala:211:16, :224:42
  wire [15:0][11:0] _GEN_35 =
    {{stq_15_bits_uop_csr_addr},
     {stq_14_bits_uop_csr_addr},
     {stq_13_bits_uop_csr_addr},
     {stq_12_bits_uop_csr_addr},
     {stq_11_bits_uop_csr_addr},
     {stq_10_bits_uop_csr_addr},
     {stq_9_bits_uop_csr_addr},
     {stq_8_bits_uop_csr_addr},
     {stq_7_bits_uop_csr_addr},
     {stq_6_bits_uop_csr_addr},
     {stq_5_bits_uop_csr_addr},
     {stq_4_bits_uop_csr_addr},
     {stq_3_bits_uop_csr_addr},
     {stq_2_bits_uop_csr_addr},
     {stq_1_bits_uop_csr_addr},
     {stq_0_bits_uop_csr_addr}};	// lsu.scala:211:16, :224:42
  wire [15:0][5:0]  _GEN_36 =
    {{stq_15_bits_uop_rob_idx},
     {stq_14_bits_uop_rob_idx},
     {stq_13_bits_uop_rob_idx},
     {stq_12_bits_uop_rob_idx},
     {stq_11_bits_uop_rob_idx},
     {stq_10_bits_uop_rob_idx},
     {stq_9_bits_uop_rob_idx},
     {stq_8_bits_uop_rob_idx},
     {stq_7_bits_uop_rob_idx},
     {stq_6_bits_uop_rob_idx},
     {stq_5_bits_uop_rob_idx},
     {stq_4_bits_uop_rob_idx},
     {stq_3_bits_uop_rob_idx},
     {stq_2_bits_uop_rob_idx},
     {stq_1_bits_uop_rob_idx},
     {stq_0_bits_uop_rob_idx}};	// lsu.scala:211:16, :224:42
  wire [15:0][3:0]  _GEN_37 =
    {{stq_15_bits_uop_ldq_idx},
     {stq_14_bits_uop_ldq_idx},
     {stq_13_bits_uop_ldq_idx},
     {stq_12_bits_uop_ldq_idx},
     {stq_11_bits_uop_ldq_idx},
     {stq_10_bits_uop_ldq_idx},
     {stq_9_bits_uop_ldq_idx},
     {stq_8_bits_uop_ldq_idx},
     {stq_7_bits_uop_ldq_idx},
     {stq_6_bits_uop_ldq_idx},
     {stq_5_bits_uop_ldq_idx},
     {stq_4_bits_uop_ldq_idx},
     {stq_3_bits_uop_ldq_idx},
     {stq_2_bits_uop_ldq_idx},
     {stq_1_bits_uop_ldq_idx},
     {stq_0_bits_uop_ldq_idx}};	// lsu.scala:211:16, :224:42
  wire [15:0][3:0]  _GEN_38 =
    {{stq_15_bits_uop_stq_idx},
     {stq_14_bits_uop_stq_idx},
     {stq_13_bits_uop_stq_idx},
     {stq_12_bits_uop_stq_idx},
     {stq_11_bits_uop_stq_idx},
     {stq_10_bits_uop_stq_idx},
     {stq_9_bits_uop_stq_idx},
     {stq_8_bits_uop_stq_idx},
     {stq_7_bits_uop_stq_idx},
     {stq_6_bits_uop_stq_idx},
     {stq_5_bits_uop_stq_idx},
     {stq_4_bits_uop_stq_idx},
     {stq_3_bits_uop_stq_idx},
     {stq_2_bits_uop_stq_idx},
     {stq_1_bits_uop_stq_idx},
     {stq_0_bits_uop_stq_idx}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_39 =
    {{stq_15_bits_uop_rxq_idx},
     {stq_14_bits_uop_rxq_idx},
     {stq_13_bits_uop_rxq_idx},
     {stq_12_bits_uop_rxq_idx},
     {stq_11_bits_uop_rxq_idx},
     {stq_10_bits_uop_rxq_idx},
     {stq_9_bits_uop_rxq_idx},
     {stq_8_bits_uop_rxq_idx},
     {stq_7_bits_uop_rxq_idx},
     {stq_6_bits_uop_rxq_idx},
     {stq_5_bits_uop_rxq_idx},
     {stq_4_bits_uop_rxq_idx},
     {stq_3_bits_uop_rxq_idx},
     {stq_2_bits_uop_rxq_idx},
     {stq_1_bits_uop_rxq_idx},
     {stq_0_bits_uop_rxq_idx}};	// lsu.scala:211:16, :224:42
  wire [15:0][6:0]  _GEN_40 =
    {{stq_15_bits_uop_pdst},
     {stq_14_bits_uop_pdst},
     {stq_13_bits_uop_pdst},
     {stq_12_bits_uop_pdst},
     {stq_11_bits_uop_pdst},
     {stq_10_bits_uop_pdst},
     {stq_9_bits_uop_pdst},
     {stq_8_bits_uop_pdst},
     {stq_7_bits_uop_pdst},
     {stq_6_bits_uop_pdst},
     {stq_5_bits_uop_pdst},
     {stq_4_bits_uop_pdst},
     {stq_3_bits_uop_pdst},
     {stq_2_bits_uop_pdst},
     {stq_1_bits_uop_pdst},
     {stq_0_bits_uop_pdst}};	// lsu.scala:211:16, :224:42
  wire [15:0][6:0]  _GEN_41 =
    {{stq_15_bits_uop_prs1},
     {stq_14_bits_uop_prs1},
     {stq_13_bits_uop_prs1},
     {stq_12_bits_uop_prs1},
     {stq_11_bits_uop_prs1},
     {stq_10_bits_uop_prs1},
     {stq_9_bits_uop_prs1},
     {stq_8_bits_uop_prs1},
     {stq_7_bits_uop_prs1},
     {stq_6_bits_uop_prs1},
     {stq_5_bits_uop_prs1},
     {stq_4_bits_uop_prs1},
     {stq_3_bits_uop_prs1},
     {stq_2_bits_uop_prs1},
     {stq_1_bits_uop_prs1},
     {stq_0_bits_uop_prs1}};	// lsu.scala:211:16, :224:42
  wire [15:0][6:0]  _GEN_42 =
    {{stq_15_bits_uop_prs2},
     {stq_14_bits_uop_prs2},
     {stq_13_bits_uop_prs2},
     {stq_12_bits_uop_prs2},
     {stq_11_bits_uop_prs2},
     {stq_10_bits_uop_prs2},
     {stq_9_bits_uop_prs2},
     {stq_8_bits_uop_prs2},
     {stq_7_bits_uop_prs2},
     {stq_6_bits_uop_prs2},
     {stq_5_bits_uop_prs2},
     {stq_4_bits_uop_prs2},
     {stq_3_bits_uop_prs2},
     {stq_2_bits_uop_prs2},
     {stq_1_bits_uop_prs2},
     {stq_0_bits_uop_prs2}};	// lsu.scala:211:16, :224:42
  wire [15:0][6:0]  _GEN_43 =
    {{stq_15_bits_uop_prs3},
     {stq_14_bits_uop_prs3},
     {stq_13_bits_uop_prs3},
     {stq_12_bits_uop_prs3},
     {stq_11_bits_uop_prs3},
     {stq_10_bits_uop_prs3},
     {stq_9_bits_uop_prs3},
     {stq_8_bits_uop_prs3},
     {stq_7_bits_uop_prs3},
     {stq_6_bits_uop_prs3},
     {stq_5_bits_uop_prs3},
     {stq_4_bits_uop_prs3},
     {stq_3_bits_uop_prs3},
     {stq_2_bits_uop_prs3},
     {stq_1_bits_uop_prs3},
     {stq_0_bits_uop_prs3}};	// lsu.scala:211:16, :224:42
  wire [15:0][4:0]  _GEN_44 =
    {{stq_15_bits_uop_ppred},
     {stq_14_bits_uop_ppred},
     {stq_13_bits_uop_ppred},
     {stq_12_bits_uop_ppred},
     {stq_11_bits_uop_ppred},
     {stq_10_bits_uop_ppred},
     {stq_9_bits_uop_ppred},
     {stq_8_bits_uop_ppred},
     {stq_7_bits_uop_ppred},
     {stq_6_bits_uop_ppred},
     {stq_5_bits_uop_ppred},
     {stq_4_bits_uop_ppred},
     {stq_3_bits_uop_ppred},
     {stq_2_bits_uop_ppred},
     {stq_1_bits_uop_ppred},
     {stq_0_bits_uop_ppred}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_45 =
    {{stq_15_bits_uop_prs1_busy},
     {stq_14_bits_uop_prs1_busy},
     {stq_13_bits_uop_prs1_busy},
     {stq_12_bits_uop_prs1_busy},
     {stq_11_bits_uop_prs1_busy},
     {stq_10_bits_uop_prs1_busy},
     {stq_9_bits_uop_prs1_busy},
     {stq_8_bits_uop_prs1_busy},
     {stq_7_bits_uop_prs1_busy},
     {stq_6_bits_uop_prs1_busy},
     {stq_5_bits_uop_prs1_busy},
     {stq_4_bits_uop_prs1_busy},
     {stq_3_bits_uop_prs1_busy},
     {stq_2_bits_uop_prs1_busy},
     {stq_1_bits_uop_prs1_busy},
     {stq_0_bits_uop_prs1_busy}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_46 =
    {{stq_15_bits_uop_prs2_busy},
     {stq_14_bits_uop_prs2_busy},
     {stq_13_bits_uop_prs2_busy},
     {stq_12_bits_uop_prs2_busy},
     {stq_11_bits_uop_prs2_busy},
     {stq_10_bits_uop_prs2_busy},
     {stq_9_bits_uop_prs2_busy},
     {stq_8_bits_uop_prs2_busy},
     {stq_7_bits_uop_prs2_busy},
     {stq_6_bits_uop_prs2_busy},
     {stq_5_bits_uop_prs2_busy},
     {stq_4_bits_uop_prs2_busy},
     {stq_3_bits_uop_prs2_busy},
     {stq_2_bits_uop_prs2_busy},
     {stq_1_bits_uop_prs2_busy},
     {stq_0_bits_uop_prs2_busy}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_47 =
    {{stq_15_bits_uop_prs3_busy},
     {stq_14_bits_uop_prs3_busy},
     {stq_13_bits_uop_prs3_busy},
     {stq_12_bits_uop_prs3_busy},
     {stq_11_bits_uop_prs3_busy},
     {stq_10_bits_uop_prs3_busy},
     {stq_9_bits_uop_prs3_busy},
     {stq_8_bits_uop_prs3_busy},
     {stq_7_bits_uop_prs3_busy},
     {stq_6_bits_uop_prs3_busy},
     {stq_5_bits_uop_prs3_busy},
     {stq_4_bits_uop_prs3_busy},
     {stq_3_bits_uop_prs3_busy},
     {stq_2_bits_uop_prs3_busy},
     {stq_1_bits_uop_prs3_busy},
     {stq_0_bits_uop_prs3_busy}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_48 =
    {{stq_15_bits_uop_ppred_busy},
     {stq_14_bits_uop_ppred_busy},
     {stq_13_bits_uop_ppred_busy},
     {stq_12_bits_uop_ppred_busy},
     {stq_11_bits_uop_ppred_busy},
     {stq_10_bits_uop_ppred_busy},
     {stq_9_bits_uop_ppred_busy},
     {stq_8_bits_uop_ppred_busy},
     {stq_7_bits_uop_ppred_busy},
     {stq_6_bits_uop_ppred_busy},
     {stq_5_bits_uop_ppred_busy},
     {stq_4_bits_uop_ppred_busy},
     {stq_3_bits_uop_ppred_busy},
     {stq_2_bits_uop_ppred_busy},
     {stq_1_bits_uop_ppred_busy},
     {stq_0_bits_uop_ppred_busy}};	// lsu.scala:211:16, :224:42
  wire [15:0][6:0]  _GEN_49 =
    {{stq_15_bits_uop_stale_pdst},
     {stq_14_bits_uop_stale_pdst},
     {stq_13_bits_uop_stale_pdst},
     {stq_12_bits_uop_stale_pdst},
     {stq_11_bits_uop_stale_pdst},
     {stq_10_bits_uop_stale_pdst},
     {stq_9_bits_uop_stale_pdst},
     {stq_8_bits_uop_stale_pdst},
     {stq_7_bits_uop_stale_pdst},
     {stq_6_bits_uop_stale_pdst},
     {stq_5_bits_uop_stale_pdst},
     {stq_4_bits_uop_stale_pdst},
     {stq_3_bits_uop_stale_pdst},
     {stq_2_bits_uop_stale_pdst},
     {stq_1_bits_uop_stale_pdst},
     {stq_0_bits_uop_stale_pdst}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_50 =
    {{stq_15_bits_uop_exception},
     {stq_14_bits_uop_exception},
     {stq_13_bits_uop_exception},
     {stq_12_bits_uop_exception},
     {stq_11_bits_uop_exception},
     {stq_10_bits_uop_exception},
     {stq_9_bits_uop_exception},
     {stq_8_bits_uop_exception},
     {stq_7_bits_uop_exception},
     {stq_6_bits_uop_exception},
     {stq_5_bits_uop_exception},
     {stq_4_bits_uop_exception},
     {stq_3_bits_uop_exception},
     {stq_2_bits_uop_exception},
     {stq_1_bits_uop_exception},
     {stq_0_bits_uop_exception}};	// lsu.scala:211:16, :224:42
  wire              _GEN_51 = _GEN_50[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [15:0][63:0] _GEN_52 =
    {{stq_15_bits_uop_exc_cause},
     {stq_14_bits_uop_exc_cause},
     {stq_13_bits_uop_exc_cause},
     {stq_12_bits_uop_exc_cause},
     {stq_11_bits_uop_exc_cause},
     {stq_10_bits_uop_exc_cause},
     {stq_9_bits_uop_exc_cause},
     {stq_8_bits_uop_exc_cause},
     {stq_7_bits_uop_exc_cause},
     {stq_6_bits_uop_exc_cause},
     {stq_5_bits_uop_exc_cause},
     {stq_4_bits_uop_exc_cause},
     {stq_3_bits_uop_exc_cause},
     {stq_2_bits_uop_exc_cause},
     {stq_1_bits_uop_exc_cause},
     {stq_0_bits_uop_exc_cause}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_53 =
    {{stq_15_bits_uop_bypassable},
     {stq_14_bits_uop_bypassable},
     {stq_13_bits_uop_bypassable},
     {stq_12_bits_uop_bypassable},
     {stq_11_bits_uop_bypassable},
     {stq_10_bits_uop_bypassable},
     {stq_9_bits_uop_bypassable},
     {stq_8_bits_uop_bypassable},
     {stq_7_bits_uop_bypassable},
     {stq_6_bits_uop_bypassable},
     {stq_5_bits_uop_bypassable},
     {stq_4_bits_uop_bypassable},
     {stq_3_bits_uop_bypassable},
     {stq_2_bits_uop_bypassable},
     {stq_1_bits_uop_bypassable},
     {stq_0_bits_uop_bypassable}};	// lsu.scala:211:16, :224:42
  wire [15:0][4:0]  _GEN_54 =
    {{stq_15_bits_uop_mem_cmd},
     {stq_14_bits_uop_mem_cmd},
     {stq_13_bits_uop_mem_cmd},
     {stq_12_bits_uop_mem_cmd},
     {stq_11_bits_uop_mem_cmd},
     {stq_10_bits_uop_mem_cmd},
     {stq_9_bits_uop_mem_cmd},
     {stq_8_bits_uop_mem_cmd},
     {stq_7_bits_uop_mem_cmd},
     {stq_6_bits_uop_mem_cmd},
     {stq_5_bits_uop_mem_cmd},
     {stq_4_bits_uop_mem_cmd},
     {stq_3_bits_uop_mem_cmd},
     {stq_2_bits_uop_mem_cmd},
     {stq_1_bits_uop_mem_cmd},
     {stq_0_bits_uop_mem_cmd}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_55 =
    {{stq_15_bits_uop_mem_size},
     {stq_14_bits_uop_mem_size},
     {stq_13_bits_uop_mem_size},
     {stq_12_bits_uop_mem_size},
     {stq_11_bits_uop_mem_size},
     {stq_10_bits_uop_mem_size},
     {stq_9_bits_uop_mem_size},
     {stq_8_bits_uop_mem_size},
     {stq_7_bits_uop_mem_size},
     {stq_6_bits_uop_mem_size},
     {stq_5_bits_uop_mem_size},
     {stq_4_bits_uop_mem_size},
     {stq_3_bits_uop_mem_size},
     {stq_2_bits_uop_mem_size},
     {stq_1_bits_uop_mem_size},
     {stq_0_bits_uop_mem_size}};	// lsu.scala:211:16, :224:42
  wire [1:0]        _GEN_56 = _GEN_55[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [15:0]       _GEN_57 =
    {{stq_15_bits_uop_mem_signed},
     {stq_14_bits_uop_mem_signed},
     {stq_13_bits_uop_mem_signed},
     {stq_12_bits_uop_mem_signed},
     {stq_11_bits_uop_mem_signed},
     {stq_10_bits_uop_mem_signed},
     {stq_9_bits_uop_mem_signed},
     {stq_8_bits_uop_mem_signed},
     {stq_7_bits_uop_mem_signed},
     {stq_6_bits_uop_mem_signed},
     {stq_5_bits_uop_mem_signed},
     {stq_4_bits_uop_mem_signed},
     {stq_3_bits_uop_mem_signed},
     {stq_2_bits_uop_mem_signed},
     {stq_1_bits_uop_mem_signed},
     {stq_0_bits_uop_mem_signed}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_58 =
    {{stq_15_bits_uop_is_fence},
     {stq_14_bits_uop_is_fence},
     {stq_13_bits_uop_is_fence},
     {stq_12_bits_uop_is_fence},
     {stq_11_bits_uop_is_fence},
     {stq_10_bits_uop_is_fence},
     {stq_9_bits_uop_is_fence},
     {stq_8_bits_uop_is_fence},
     {stq_7_bits_uop_is_fence},
     {stq_6_bits_uop_is_fence},
     {stq_5_bits_uop_is_fence},
     {stq_4_bits_uop_is_fence},
     {stq_3_bits_uop_is_fence},
     {stq_2_bits_uop_is_fence},
     {stq_1_bits_uop_is_fence},
     {stq_0_bits_uop_is_fence}};	// lsu.scala:211:16, :224:42
  wire              _GEN_59 = _GEN_58[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [15:0]       _GEN_60 =
    {{stq_15_bits_uop_is_fencei},
     {stq_14_bits_uop_is_fencei},
     {stq_13_bits_uop_is_fencei},
     {stq_12_bits_uop_is_fencei},
     {stq_11_bits_uop_is_fencei},
     {stq_10_bits_uop_is_fencei},
     {stq_9_bits_uop_is_fencei},
     {stq_8_bits_uop_is_fencei},
     {stq_7_bits_uop_is_fencei},
     {stq_6_bits_uop_is_fencei},
     {stq_5_bits_uop_is_fencei},
     {stq_4_bits_uop_is_fencei},
     {stq_3_bits_uop_is_fencei},
     {stq_2_bits_uop_is_fencei},
     {stq_1_bits_uop_is_fencei},
     {stq_0_bits_uop_is_fencei}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_61 =
    {{stq_15_bits_uop_is_amo},
     {stq_14_bits_uop_is_amo},
     {stq_13_bits_uop_is_amo},
     {stq_12_bits_uop_is_amo},
     {stq_11_bits_uop_is_amo},
     {stq_10_bits_uop_is_amo},
     {stq_9_bits_uop_is_amo},
     {stq_8_bits_uop_is_amo},
     {stq_7_bits_uop_is_amo},
     {stq_6_bits_uop_is_amo},
     {stq_5_bits_uop_is_amo},
     {stq_4_bits_uop_is_amo},
     {stq_3_bits_uop_is_amo},
     {stq_2_bits_uop_is_amo},
     {stq_1_bits_uop_is_amo},
     {stq_0_bits_uop_is_amo}};	// lsu.scala:211:16, :224:42
  wire              _GEN_62 = _GEN_61[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [15:0]       _GEN_63 =
    {{stq_15_bits_uop_uses_ldq},
     {stq_14_bits_uop_uses_ldq},
     {stq_13_bits_uop_uses_ldq},
     {stq_12_bits_uop_uses_ldq},
     {stq_11_bits_uop_uses_ldq},
     {stq_10_bits_uop_uses_ldq},
     {stq_9_bits_uop_uses_ldq},
     {stq_8_bits_uop_uses_ldq},
     {stq_7_bits_uop_uses_ldq},
     {stq_6_bits_uop_uses_ldq},
     {stq_5_bits_uop_uses_ldq},
     {stq_4_bits_uop_uses_ldq},
     {stq_3_bits_uop_uses_ldq},
     {stq_2_bits_uop_uses_ldq},
     {stq_1_bits_uop_uses_ldq},
     {stq_0_bits_uop_uses_ldq}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_64 =
    {{stq_15_bits_uop_uses_stq},
     {stq_14_bits_uop_uses_stq},
     {stq_13_bits_uop_uses_stq},
     {stq_12_bits_uop_uses_stq},
     {stq_11_bits_uop_uses_stq},
     {stq_10_bits_uop_uses_stq},
     {stq_9_bits_uop_uses_stq},
     {stq_8_bits_uop_uses_stq},
     {stq_7_bits_uop_uses_stq},
     {stq_6_bits_uop_uses_stq},
     {stq_5_bits_uop_uses_stq},
     {stq_4_bits_uop_uses_stq},
     {stq_3_bits_uop_uses_stq},
     {stq_2_bits_uop_uses_stq},
     {stq_1_bits_uop_uses_stq},
     {stq_0_bits_uop_uses_stq}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_65 =
    {{stq_15_bits_uop_is_sys_pc2epc},
     {stq_14_bits_uop_is_sys_pc2epc},
     {stq_13_bits_uop_is_sys_pc2epc},
     {stq_12_bits_uop_is_sys_pc2epc},
     {stq_11_bits_uop_is_sys_pc2epc},
     {stq_10_bits_uop_is_sys_pc2epc},
     {stq_9_bits_uop_is_sys_pc2epc},
     {stq_8_bits_uop_is_sys_pc2epc},
     {stq_7_bits_uop_is_sys_pc2epc},
     {stq_6_bits_uop_is_sys_pc2epc},
     {stq_5_bits_uop_is_sys_pc2epc},
     {stq_4_bits_uop_is_sys_pc2epc},
     {stq_3_bits_uop_is_sys_pc2epc},
     {stq_2_bits_uop_is_sys_pc2epc},
     {stq_1_bits_uop_is_sys_pc2epc},
     {stq_0_bits_uop_is_sys_pc2epc}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_66 =
    {{stq_15_bits_uop_is_unique},
     {stq_14_bits_uop_is_unique},
     {stq_13_bits_uop_is_unique},
     {stq_12_bits_uop_is_unique},
     {stq_11_bits_uop_is_unique},
     {stq_10_bits_uop_is_unique},
     {stq_9_bits_uop_is_unique},
     {stq_8_bits_uop_is_unique},
     {stq_7_bits_uop_is_unique},
     {stq_6_bits_uop_is_unique},
     {stq_5_bits_uop_is_unique},
     {stq_4_bits_uop_is_unique},
     {stq_3_bits_uop_is_unique},
     {stq_2_bits_uop_is_unique},
     {stq_1_bits_uop_is_unique},
     {stq_0_bits_uop_is_unique}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_67 =
    {{stq_15_bits_uop_flush_on_commit},
     {stq_14_bits_uop_flush_on_commit},
     {stq_13_bits_uop_flush_on_commit},
     {stq_12_bits_uop_flush_on_commit},
     {stq_11_bits_uop_flush_on_commit},
     {stq_10_bits_uop_flush_on_commit},
     {stq_9_bits_uop_flush_on_commit},
     {stq_8_bits_uop_flush_on_commit},
     {stq_7_bits_uop_flush_on_commit},
     {stq_6_bits_uop_flush_on_commit},
     {stq_5_bits_uop_flush_on_commit},
     {stq_4_bits_uop_flush_on_commit},
     {stq_3_bits_uop_flush_on_commit},
     {stq_2_bits_uop_flush_on_commit},
     {stq_1_bits_uop_flush_on_commit},
     {stq_0_bits_uop_flush_on_commit}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_68 =
    {{stq_15_bits_uop_ldst_is_rs1},
     {stq_14_bits_uop_ldst_is_rs1},
     {stq_13_bits_uop_ldst_is_rs1},
     {stq_12_bits_uop_ldst_is_rs1},
     {stq_11_bits_uop_ldst_is_rs1},
     {stq_10_bits_uop_ldst_is_rs1},
     {stq_9_bits_uop_ldst_is_rs1},
     {stq_8_bits_uop_ldst_is_rs1},
     {stq_7_bits_uop_ldst_is_rs1},
     {stq_6_bits_uop_ldst_is_rs1},
     {stq_5_bits_uop_ldst_is_rs1},
     {stq_4_bits_uop_ldst_is_rs1},
     {stq_3_bits_uop_ldst_is_rs1},
     {stq_2_bits_uop_ldst_is_rs1},
     {stq_1_bits_uop_ldst_is_rs1},
     {stq_0_bits_uop_ldst_is_rs1}};	// lsu.scala:211:16, :224:42
  wire [15:0][5:0]  _GEN_69 =
    {{stq_15_bits_uop_ldst},
     {stq_14_bits_uop_ldst},
     {stq_13_bits_uop_ldst},
     {stq_12_bits_uop_ldst},
     {stq_11_bits_uop_ldst},
     {stq_10_bits_uop_ldst},
     {stq_9_bits_uop_ldst},
     {stq_8_bits_uop_ldst},
     {stq_7_bits_uop_ldst},
     {stq_6_bits_uop_ldst},
     {stq_5_bits_uop_ldst},
     {stq_4_bits_uop_ldst},
     {stq_3_bits_uop_ldst},
     {stq_2_bits_uop_ldst},
     {stq_1_bits_uop_ldst},
     {stq_0_bits_uop_ldst}};	// lsu.scala:211:16, :224:42
  wire [15:0][5:0]  _GEN_70 =
    {{stq_15_bits_uop_lrs1},
     {stq_14_bits_uop_lrs1},
     {stq_13_bits_uop_lrs1},
     {stq_12_bits_uop_lrs1},
     {stq_11_bits_uop_lrs1},
     {stq_10_bits_uop_lrs1},
     {stq_9_bits_uop_lrs1},
     {stq_8_bits_uop_lrs1},
     {stq_7_bits_uop_lrs1},
     {stq_6_bits_uop_lrs1},
     {stq_5_bits_uop_lrs1},
     {stq_4_bits_uop_lrs1},
     {stq_3_bits_uop_lrs1},
     {stq_2_bits_uop_lrs1},
     {stq_1_bits_uop_lrs1},
     {stq_0_bits_uop_lrs1}};	// lsu.scala:211:16, :224:42
  wire [15:0][5:0]  _GEN_71 =
    {{stq_15_bits_uop_lrs2},
     {stq_14_bits_uop_lrs2},
     {stq_13_bits_uop_lrs2},
     {stq_12_bits_uop_lrs2},
     {stq_11_bits_uop_lrs2},
     {stq_10_bits_uop_lrs2},
     {stq_9_bits_uop_lrs2},
     {stq_8_bits_uop_lrs2},
     {stq_7_bits_uop_lrs2},
     {stq_6_bits_uop_lrs2},
     {stq_5_bits_uop_lrs2},
     {stq_4_bits_uop_lrs2},
     {stq_3_bits_uop_lrs2},
     {stq_2_bits_uop_lrs2},
     {stq_1_bits_uop_lrs2},
     {stq_0_bits_uop_lrs2}};	// lsu.scala:211:16, :224:42
  wire [15:0][5:0]  _GEN_72 =
    {{stq_15_bits_uop_lrs3},
     {stq_14_bits_uop_lrs3},
     {stq_13_bits_uop_lrs3},
     {stq_12_bits_uop_lrs3},
     {stq_11_bits_uop_lrs3},
     {stq_10_bits_uop_lrs3},
     {stq_9_bits_uop_lrs3},
     {stq_8_bits_uop_lrs3},
     {stq_7_bits_uop_lrs3},
     {stq_6_bits_uop_lrs3},
     {stq_5_bits_uop_lrs3},
     {stq_4_bits_uop_lrs3},
     {stq_3_bits_uop_lrs3},
     {stq_2_bits_uop_lrs3},
     {stq_1_bits_uop_lrs3},
     {stq_0_bits_uop_lrs3}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_73 =
    {{stq_15_bits_uop_ldst_val},
     {stq_14_bits_uop_ldst_val},
     {stq_13_bits_uop_ldst_val},
     {stq_12_bits_uop_ldst_val},
     {stq_11_bits_uop_ldst_val},
     {stq_10_bits_uop_ldst_val},
     {stq_9_bits_uop_ldst_val},
     {stq_8_bits_uop_ldst_val},
     {stq_7_bits_uop_ldst_val},
     {stq_6_bits_uop_ldst_val},
     {stq_5_bits_uop_ldst_val},
     {stq_4_bits_uop_ldst_val},
     {stq_3_bits_uop_ldst_val},
     {stq_2_bits_uop_ldst_val},
     {stq_1_bits_uop_ldst_val},
     {stq_0_bits_uop_ldst_val}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_74 =
    {{stq_15_bits_uop_dst_rtype},
     {stq_14_bits_uop_dst_rtype},
     {stq_13_bits_uop_dst_rtype},
     {stq_12_bits_uop_dst_rtype},
     {stq_11_bits_uop_dst_rtype},
     {stq_10_bits_uop_dst_rtype},
     {stq_9_bits_uop_dst_rtype},
     {stq_8_bits_uop_dst_rtype},
     {stq_7_bits_uop_dst_rtype},
     {stq_6_bits_uop_dst_rtype},
     {stq_5_bits_uop_dst_rtype},
     {stq_4_bits_uop_dst_rtype},
     {stq_3_bits_uop_dst_rtype},
     {stq_2_bits_uop_dst_rtype},
     {stq_1_bits_uop_dst_rtype},
     {stq_0_bits_uop_dst_rtype}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_75 =
    {{stq_15_bits_uop_lrs1_rtype},
     {stq_14_bits_uop_lrs1_rtype},
     {stq_13_bits_uop_lrs1_rtype},
     {stq_12_bits_uop_lrs1_rtype},
     {stq_11_bits_uop_lrs1_rtype},
     {stq_10_bits_uop_lrs1_rtype},
     {stq_9_bits_uop_lrs1_rtype},
     {stq_8_bits_uop_lrs1_rtype},
     {stq_7_bits_uop_lrs1_rtype},
     {stq_6_bits_uop_lrs1_rtype},
     {stq_5_bits_uop_lrs1_rtype},
     {stq_4_bits_uop_lrs1_rtype},
     {stq_3_bits_uop_lrs1_rtype},
     {stq_2_bits_uop_lrs1_rtype},
     {stq_1_bits_uop_lrs1_rtype},
     {stq_0_bits_uop_lrs1_rtype}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_76 =
    {{stq_15_bits_uop_lrs2_rtype},
     {stq_14_bits_uop_lrs2_rtype},
     {stq_13_bits_uop_lrs2_rtype},
     {stq_12_bits_uop_lrs2_rtype},
     {stq_11_bits_uop_lrs2_rtype},
     {stq_10_bits_uop_lrs2_rtype},
     {stq_9_bits_uop_lrs2_rtype},
     {stq_8_bits_uop_lrs2_rtype},
     {stq_7_bits_uop_lrs2_rtype},
     {stq_6_bits_uop_lrs2_rtype},
     {stq_5_bits_uop_lrs2_rtype},
     {stq_4_bits_uop_lrs2_rtype},
     {stq_3_bits_uop_lrs2_rtype},
     {stq_2_bits_uop_lrs2_rtype},
     {stq_1_bits_uop_lrs2_rtype},
     {stq_0_bits_uop_lrs2_rtype}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_77 =
    {{stq_15_bits_uop_frs3_en},
     {stq_14_bits_uop_frs3_en},
     {stq_13_bits_uop_frs3_en},
     {stq_12_bits_uop_frs3_en},
     {stq_11_bits_uop_frs3_en},
     {stq_10_bits_uop_frs3_en},
     {stq_9_bits_uop_frs3_en},
     {stq_8_bits_uop_frs3_en},
     {stq_7_bits_uop_frs3_en},
     {stq_6_bits_uop_frs3_en},
     {stq_5_bits_uop_frs3_en},
     {stq_4_bits_uop_frs3_en},
     {stq_3_bits_uop_frs3_en},
     {stq_2_bits_uop_frs3_en},
     {stq_1_bits_uop_frs3_en},
     {stq_0_bits_uop_frs3_en}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_78 =
    {{stq_15_bits_uop_fp_val},
     {stq_14_bits_uop_fp_val},
     {stq_13_bits_uop_fp_val},
     {stq_12_bits_uop_fp_val},
     {stq_11_bits_uop_fp_val},
     {stq_10_bits_uop_fp_val},
     {stq_9_bits_uop_fp_val},
     {stq_8_bits_uop_fp_val},
     {stq_7_bits_uop_fp_val},
     {stq_6_bits_uop_fp_val},
     {stq_5_bits_uop_fp_val},
     {stq_4_bits_uop_fp_val},
     {stq_3_bits_uop_fp_val},
     {stq_2_bits_uop_fp_val},
     {stq_1_bits_uop_fp_val},
     {stq_0_bits_uop_fp_val}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_79 =
    {{stq_15_bits_uop_fp_single},
     {stq_14_bits_uop_fp_single},
     {stq_13_bits_uop_fp_single},
     {stq_12_bits_uop_fp_single},
     {stq_11_bits_uop_fp_single},
     {stq_10_bits_uop_fp_single},
     {stq_9_bits_uop_fp_single},
     {stq_8_bits_uop_fp_single},
     {stq_7_bits_uop_fp_single},
     {stq_6_bits_uop_fp_single},
     {stq_5_bits_uop_fp_single},
     {stq_4_bits_uop_fp_single},
     {stq_3_bits_uop_fp_single},
     {stq_2_bits_uop_fp_single},
     {stq_1_bits_uop_fp_single},
     {stq_0_bits_uop_fp_single}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_80 =
    {{stq_15_bits_uop_xcpt_pf_if},
     {stq_14_bits_uop_xcpt_pf_if},
     {stq_13_bits_uop_xcpt_pf_if},
     {stq_12_bits_uop_xcpt_pf_if},
     {stq_11_bits_uop_xcpt_pf_if},
     {stq_10_bits_uop_xcpt_pf_if},
     {stq_9_bits_uop_xcpt_pf_if},
     {stq_8_bits_uop_xcpt_pf_if},
     {stq_7_bits_uop_xcpt_pf_if},
     {stq_6_bits_uop_xcpt_pf_if},
     {stq_5_bits_uop_xcpt_pf_if},
     {stq_4_bits_uop_xcpt_pf_if},
     {stq_3_bits_uop_xcpt_pf_if},
     {stq_2_bits_uop_xcpt_pf_if},
     {stq_1_bits_uop_xcpt_pf_if},
     {stq_0_bits_uop_xcpt_pf_if}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_81 =
    {{stq_15_bits_uop_xcpt_ae_if},
     {stq_14_bits_uop_xcpt_ae_if},
     {stq_13_bits_uop_xcpt_ae_if},
     {stq_12_bits_uop_xcpt_ae_if},
     {stq_11_bits_uop_xcpt_ae_if},
     {stq_10_bits_uop_xcpt_ae_if},
     {stq_9_bits_uop_xcpt_ae_if},
     {stq_8_bits_uop_xcpt_ae_if},
     {stq_7_bits_uop_xcpt_ae_if},
     {stq_6_bits_uop_xcpt_ae_if},
     {stq_5_bits_uop_xcpt_ae_if},
     {stq_4_bits_uop_xcpt_ae_if},
     {stq_3_bits_uop_xcpt_ae_if},
     {stq_2_bits_uop_xcpt_ae_if},
     {stq_1_bits_uop_xcpt_ae_if},
     {stq_0_bits_uop_xcpt_ae_if}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_82 =
    {{stq_15_bits_uop_xcpt_ma_if},
     {stq_14_bits_uop_xcpt_ma_if},
     {stq_13_bits_uop_xcpt_ma_if},
     {stq_12_bits_uop_xcpt_ma_if},
     {stq_11_bits_uop_xcpt_ma_if},
     {stq_10_bits_uop_xcpt_ma_if},
     {stq_9_bits_uop_xcpt_ma_if},
     {stq_8_bits_uop_xcpt_ma_if},
     {stq_7_bits_uop_xcpt_ma_if},
     {stq_6_bits_uop_xcpt_ma_if},
     {stq_5_bits_uop_xcpt_ma_if},
     {stq_4_bits_uop_xcpt_ma_if},
     {stq_3_bits_uop_xcpt_ma_if},
     {stq_2_bits_uop_xcpt_ma_if},
     {stq_1_bits_uop_xcpt_ma_if},
     {stq_0_bits_uop_xcpt_ma_if}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_83 =
    {{stq_15_bits_uop_bp_debug_if},
     {stq_14_bits_uop_bp_debug_if},
     {stq_13_bits_uop_bp_debug_if},
     {stq_12_bits_uop_bp_debug_if},
     {stq_11_bits_uop_bp_debug_if},
     {stq_10_bits_uop_bp_debug_if},
     {stq_9_bits_uop_bp_debug_if},
     {stq_8_bits_uop_bp_debug_if},
     {stq_7_bits_uop_bp_debug_if},
     {stq_6_bits_uop_bp_debug_if},
     {stq_5_bits_uop_bp_debug_if},
     {stq_4_bits_uop_bp_debug_if},
     {stq_3_bits_uop_bp_debug_if},
     {stq_2_bits_uop_bp_debug_if},
     {stq_1_bits_uop_bp_debug_if},
     {stq_0_bits_uop_bp_debug_if}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_84 =
    {{stq_15_bits_uop_bp_xcpt_if},
     {stq_14_bits_uop_bp_xcpt_if},
     {stq_13_bits_uop_bp_xcpt_if},
     {stq_12_bits_uop_bp_xcpt_if},
     {stq_11_bits_uop_bp_xcpt_if},
     {stq_10_bits_uop_bp_xcpt_if},
     {stq_9_bits_uop_bp_xcpt_if},
     {stq_8_bits_uop_bp_xcpt_if},
     {stq_7_bits_uop_bp_xcpt_if},
     {stq_6_bits_uop_bp_xcpt_if},
     {stq_5_bits_uop_bp_xcpt_if},
     {stq_4_bits_uop_bp_xcpt_if},
     {stq_3_bits_uop_bp_xcpt_if},
     {stq_2_bits_uop_bp_xcpt_if},
     {stq_1_bits_uop_bp_xcpt_if},
     {stq_0_bits_uop_bp_xcpt_if}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_85 =
    {{stq_15_bits_uop_debug_fsrc},
     {stq_14_bits_uop_debug_fsrc},
     {stq_13_bits_uop_debug_fsrc},
     {stq_12_bits_uop_debug_fsrc},
     {stq_11_bits_uop_debug_fsrc},
     {stq_10_bits_uop_debug_fsrc},
     {stq_9_bits_uop_debug_fsrc},
     {stq_8_bits_uop_debug_fsrc},
     {stq_7_bits_uop_debug_fsrc},
     {stq_6_bits_uop_debug_fsrc},
     {stq_5_bits_uop_debug_fsrc},
     {stq_4_bits_uop_debug_fsrc},
     {stq_3_bits_uop_debug_fsrc},
     {stq_2_bits_uop_debug_fsrc},
     {stq_1_bits_uop_debug_fsrc},
     {stq_0_bits_uop_debug_fsrc}};	// lsu.scala:211:16, :224:42
  wire [15:0][1:0]  _GEN_86 =
    {{stq_15_bits_uop_debug_tsrc},
     {stq_14_bits_uop_debug_tsrc},
     {stq_13_bits_uop_debug_tsrc},
     {stq_12_bits_uop_debug_tsrc},
     {stq_11_bits_uop_debug_tsrc},
     {stq_10_bits_uop_debug_tsrc},
     {stq_9_bits_uop_debug_tsrc},
     {stq_8_bits_uop_debug_tsrc},
     {stq_7_bits_uop_debug_tsrc},
     {stq_6_bits_uop_debug_tsrc},
     {stq_5_bits_uop_debug_tsrc},
     {stq_4_bits_uop_debug_tsrc},
     {stq_3_bits_uop_debug_tsrc},
     {stq_2_bits_uop_debug_tsrc},
     {stq_1_bits_uop_debug_tsrc},
     {stq_0_bits_uop_debug_tsrc}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_87 =
    {{stq_15_bits_addr_valid},
     {stq_14_bits_addr_valid},
     {stq_13_bits_addr_valid},
     {stq_12_bits_addr_valid},
     {stq_11_bits_addr_valid},
     {stq_10_bits_addr_valid},
     {stq_9_bits_addr_valid},
     {stq_8_bits_addr_valid},
     {stq_7_bits_addr_valid},
     {stq_6_bits_addr_valid},
     {stq_5_bits_addr_valid},
     {stq_4_bits_addr_valid},
     {stq_3_bits_addr_valid},
     {stq_2_bits_addr_valid},
     {stq_1_bits_addr_valid},
     {stq_0_bits_addr_valid}};	// lsu.scala:211:16, :224:42
  wire [15:0][39:0] _GEN_88 =
    {{stq_15_bits_addr_bits},
     {stq_14_bits_addr_bits},
     {stq_13_bits_addr_bits},
     {stq_12_bits_addr_bits},
     {stq_11_bits_addr_bits},
     {stq_10_bits_addr_bits},
     {stq_9_bits_addr_bits},
     {stq_8_bits_addr_bits},
     {stq_7_bits_addr_bits},
     {stq_6_bits_addr_bits},
     {stq_5_bits_addr_bits},
     {stq_4_bits_addr_bits},
     {stq_3_bits_addr_bits},
     {stq_2_bits_addr_bits},
     {stq_1_bits_addr_bits},
     {stq_0_bits_addr_bits}};	// lsu.scala:211:16, :224:42
  wire [39:0]       _GEN_89 = _GEN_88[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [15:0]       _GEN_90 =
    {{stq_15_bits_addr_is_virtual},
     {stq_14_bits_addr_is_virtual},
     {stq_13_bits_addr_is_virtual},
     {stq_12_bits_addr_is_virtual},
     {stq_11_bits_addr_is_virtual},
     {stq_10_bits_addr_is_virtual},
     {stq_9_bits_addr_is_virtual},
     {stq_8_bits_addr_is_virtual},
     {stq_7_bits_addr_is_virtual},
     {stq_6_bits_addr_is_virtual},
     {stq_5_bits_addr_is_virtual},
     {stq_4_bits_addr_is_virtual},
     {stq_3_bits_addr_is_virtual},
     {stq_2_bits_addr_is_virtual},
     {stq_1_bits_addr_is_virtual},
     {stq_0_bits_addr_is_virtual}};	// lsu.scala:211:16, :224:42
  wire [15:0]       _GEN_91 =
    {{stq_15_bits_data_valid},
     {stq_14_bits_data_valid},
     {stq_13_bits_data_valid},
     {stq_12_bits_data_valid},
     {stq_11_bits_data_valid},
     {stq_10_bits_data_valid},
     {stq_9_bits_data_valid},
     {stq_8_bits_data_valid},
     {stq_7_bits_data_valid},
     {stq_6_bits_data_valid},
     {stq_5_bits_data_valid},
     {stq_4_bits_data_valid},
     {stq_3_bits_data_valid},
     {stq_2_bits_data_valid},
     {stq_1_bits_data_valid},
     {stq_0_bits_data_valid}};	// lsu.scala:211:16, :224:42
  wire [15:0][63:0] _GEN_92 =
    {{stq_15_bits_data_bits},
     {stq_14_bits_data_bits},
     {stq_13_bits_data_bits},
     {stq_12_bits_data_bits},
     {stq_11_bits_data_bits},
     {stq_10_bits_data_bits},
     {stq_9_bits_data_bits},
     {stq_8_bits_data_bits},
     {stq_7_bits_data_bits},
     {stq_6_bits_data_bits},
     {stq_5_bits_data_bits},
     {stq_4_bits_data_bits},
     {stq_3_bits_data_bits},
     {stq_2_bits_data_bits},
     {stq_1_bits_data_bits},
     {stq_0_bits_data_bits}};	// lsu.scala:211:16, :224:42
  wire [63:0]       _GEN_93 = _GEN_92[stq_execute_head];	// lsu.scala:220:29, :224:42
  wire [15:0]       _GEN_94 =
    {{stq_15_bits_committed},
     {stq_14_bits_committed},
     {stq_13_bits_committed},
     {stq_12_bits_committed},
     {stq_11_bits_committed},
     {stq_10_bits_committed},
     {stq_9_bits_committed},
     {stq_8_bits_committed},
     {stq_7_bits_committed},
     {stq_6_bits_committed},
     {stq_5_bits_committed},
     {stq_4_bits_committed},
     {stq_3_bits_committed},
     {stq_2_bits_committed},
     {stq_1_bits_committed},
     {stq_0_bits_committed}};	// lsu.scala:211:16, :224:42
  reg  [2:0]        hella_state;	// lsu.scala:242:38
  reg  [39:0]       hella_req_addr;	// lsu.scala:243:34
  reg  [4:0]        hella_req_cmd;	// lsu.scala:243:34
  reg  [1:0]        hella_req_size;	// lsu.scala:243:34
  reg               hella_req_signed;	// lsu.scala:243:34
  reg               hella_req_phys;	// lsu.scala:243:34
  reg  [63:0]       hella_data_data;	// lsu.scala:244:34
  reg  [31:0]       hella_paddr;	// lsu.scala:245:34
  reg               hella_xcpt_ma_ld;	// lsu.scala:246:34
  reg               hella_xcpt_ma_st;	// lsu.scala:246:34
  reg               hella_xcpt_pf_ld;	// lsu.scala:246:34
  reg               hella_xcpt_pf_st;	// lsu.scala:246:34
  reg               hella_xcpt_ae_ld;	// lsu.scala:246:34
  reg               hella_xcpt_ae_st;	// lsu.scala:246:34
  reg  [15:0]       live_store_mask;	// lsu.scala:259:32
  wire [3:0]        _GEN_95 = ldq_tail + 4'h1;	// lsu.scala:216:29, :305:44, util.scala:203:14
  wire [3:0]        _GEN_96 = stq_tail + 4'h1;	// lsu.scala:218:29, :305:44, util.scala:203:14
  wire              dis_ld_val =
    io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_ldq
    & ~io_core_dis_uops_0_bits_exception;	// lsu.scala:301:{85,88}
  wire              dis_st_val =
    io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_stq
    & ~io_core_dis_uops_0_bits_exception;	// lsu.scala:301:88, :302:85
  wire [15:0]       _GEN_97 =
    {{ldq_15_valid},
     {ldq_14_valid},
     {ldq_13_valid},
     {ldq_12_valid},
     {ldq_11_valid},
     {ldq_10_valid},
     {ldq_9_valid},
     {ldq_8_valid},
     {ldq_7_valid},
     {ldq_6_valid},
     {ldq_5_valid},
     {ldq_4_valid},
     {ldq_3_valid},
     {ldq_2_valid},
     {ldq_1_valid},
     {ldq_0_valid}};	// lsu.scala:210:16, :305:44
  wire [3:0]        _GEN_98 = dis_ld_val ? _GEN_95 : ldq_tail;	// lsu.scala:216:29, :301:85, :333:21, util.scala:203:14
  wire [3:0]        _GEN_99 = dis_st_val ? _GEN_96 : stq_tail;	// lsu.scala:218:29, :302:85, :338:21, util.scala:203:14
  wire [3:0]        _GEN_100 = _GEN_98 + 4'h1;	// lsu.scala:305:44, :333:21, util.scala:203:14
  wire [3:0]        _GEN_101 = _GEN_99 + 4'h1;	// lsu.scala:305:44, :338:21, util.scala:203:14
  wire              dis_ld_val_1 =
    io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_ldq
    & ~io_core_dis_uops_1_bits_exception;	// lsu.scala:301:{85,88}
  wire              dis_st_val_1 =
    io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_stq
    & ~io_core_dis_uops_1_bits_exception;	// lsu.scala:301:88, :302:85
  reg               p1_block_load_mask_0;	// lsu.scala:398:35
  reg               p1_block_load_mask_1;	// lsu.scala:398:35
  reg               p1_block_load_mask_2;	// lsu.scala:398:35
  reg               p1_block_load_mask_3;	// lsu.scala:398:35
  reg               p1_block_load_mask_4;	// lsu.scala:398:35
  reg               p1_block_load_mask_5;	// lsu.scala:398:35
  reg               p1_block_load_mask_6;	// lsu.scala:398:35
  reg               p1_block_load_mask_7;	// lsu.scala:398:35
  reg               p1_block_load_mask_8;	// lsu.scala:398:35
  reg               p1_block_load_mask_9;	// lsu.scala:398:35
  reg               p1_block_load_mask_10;	// lsu.scala:398:35
  reg               p1_block_load_mask_11;	// lsu.scala:398:35
  reg               p1_block_load_mask_12;	// lsu.scala:398:35
  reg               p1_block_load_mask_13;	// lsu.scala:398:35
  reg               p1_block_load_mask_14;	// lsu.scala:398:35
  reg               p1_block_load_mask_15;	// lsu.scala:398:35
  reg               p2_block_load_mask_0;	// lsu.scala:399:35
  reg               p2_block_load_mask_1;	// lsu.scala:399:35
  reg               p2_block_load_mask_2;	// lsu.scala:399:35
  reg               p2_block_load_mask_3;	// lsu.scala:399:35
  reg               p2_block_load_mask_4;	// lsu.scala:399:35
  reg               p2_block_load_mask_5;	// lsu.scala:399:35
  reg               p2_block_load_mask_6;	// lsu.scala:399:35
  reg               p2_block_load_mask_7;	// lsu.scala:399:35
  reg               p2_block_load_mask_8;	// lsu.scala:399:35
  reg               p2_block_load_mask_9;	// lsu.scala:399:35
  reg               p2_block_load_mask_10;	// lsu.scala:399:35
  reg               p2_block_load_mask_11;	// lsu.scala:399:35
  reg               p2_block_load_mask_12;	// lsu.scala:399:35
  reg               p2_block_load_mask_13;	// lsu.scala:399:35
  reg               p2_block_load_mask_14;	// lsu.scala:399:35
  reg               p2_block_load_mask_15;	// lsu.scala:399:35
  wire [15:0][11:0] _GEN_102 =
    {{ldq_15_bits_uop_br_mask},
     {ldq_14_bits_uop_br_mask},
     {ldq_13_bits_uop_br_mask},
     {ldq_12_bits_uop_br_mask},
     {ldq_11_bits_uop_br_mask},
     {ldq_10_bits_uop_br_mask},
     {ldq_9_bits_uop_br_mask},
     {ldq_8_bits_uop_br_mask},
     {ldq_7_bits_uop_br_mask},
     {ldq_6_bits_uop_br_mask},
     {ldq_5_bits_uop_br_mask},
     {ldq_4_bits_uop_br_mask},
     {ldq_3_bits_uop_br_mask},
     {ldq_2_bits_uop_br_mask},
     {ldq_1_bits_uop_br_mask},
     {ldq_0_bits_uop_br_mask}};	// lsu.scala:210:16, :264:49
  wire [15:0][3:0]  _GEN_103 =
    {{ldq_15_bits_uop_stq_idx},
     {ldq_14_bits_uop_stq_idx},
     {ldq_13_bits_uop_stq_idx},
     {ldq_12_bits_uop_stq_idx},
     {ldq_11_bits_uop_stq_idx},
     {ldq_10_bits_uop_stq_idx},
     {ldq_9_bits_uop_stq_idx},
     {ldq_8_bits_uop_stq_idx},
     {ldq_7_bits_uop_stq_idx},
     {ldq_6_bits_uop_stq_idx},
     {ldq_5_bits_uop_stq_idx},
     {ldq_4_bits_uop_stq_idx},
     {ldq_3_bits_uop_stq_idx},
     {ldq_2_bits_uop_stq_idx},
     {ldq_1_bits_uop_stq_idx},
     {ldq_0_bits_uop_stq_idx}};	// lsu.scala:210:16, :264:49
  wire [15:0][1:0]  _GEN_104 =
    {{ldq_15_bits_uop_mem_size},
     {ldq_14_bits_uop_mem_size},
     {ldq_13_bits_uop_mem_size},
     {ldq_12_bits_uop_mem_size},
     {ldq_11_bits_uop_mem_size},
     {ldq_10_bits_uop_mem_size},
     {ldq_9_bits_uop_mem_size},
     {ldq_8_bits_uop_mem_size},
     {ldq_7_bits_uop_mem_size},
     {ldq_6_bits_uop_mem_size},
     {ldq_5_bits_uop_mem_size},
     {ldq_4_bits_uop_mem_size},
     {ldq_3_bits_uop_mem_size},
     {ldq_2_bits_uop_mem_size},
     {ldq_1_bits_uop_mem_size},
     {ldq_0_bits_uop_mem_size}};	// lsu.scala:210:16, :264:49
  wire [15:0]       _GEN_105 =
    {{ldq_15_bits_addr_valid},
     {ldq_14_bits_addr_valid},
     {ldq_13_bits_addr_valid},
     {ldq_12_bits_addr_valid},
     {ldq_11_bits_addr_valid},
     {ldq_10_bits_addr_valid},
     {ldq_9_bits_addr_valid},
     {ldq_8_bits_addr_valid},
     {ldq_7_bits_addr_valid},
     {ldq_6_bits_addr_valid},
     {ldq_5_bits_addr_valid},
     {ldq_4_bits_addr_valid},
     {ldq_3_bits_addr_valid},
     {ldq_2_bits_addr_valid},
     {ldq_1_bits_addr_valid},
     {ldq_0_bits_addr_valid}};	// lsu.scala:210:16, :264:49
  wire [15:0]       _GEN_106 =
    {{ldq_15_bits_executed},
     {ldq_14_bits_executed},
     {ldq_13_bits_executed},
     {ldq_12_bits_executed},
     {ldq_11_bits_executed},
     {ldq_10_bits_executed},
     {ldq_9_bits_executed},
     {ldq_8_bits_executed},
     {ldq_7_bits_executed},
     {ldq_6_bits_executed},
     {ldq_5_bits_executed},
     {ldq_4_bits_executed},
     {ldq_3_bits_executed},
     {ldq_2_bits_executed},
     {ldq_1_bits_executed},
     {ldq_0_bits_executed}};	// lsu.scala:210:16, :264:49
  wire [15:0][15:0] _GEN_107 =
    {{ldq_15_bits_st_dep_mask},
     {ldq_14_bits_st_dep_mask},
     {ldq_13_bits_st_dep_mask},
     {ldq_12_bits_st_dep_mask},
     {ldq_11_bits_st_dep_mask},
     {ldq_10_bits_st_dep_mask},
     {ldq_9_bits_st_dep_mask},
     {ldq_8_bits_st_dep_mask},
     {ldq_7_bits_st_dep_mask},
     {ldq_6_bits_st_dep_mask},
     {ldq_5_bits_st_dep_mask},
     {ldq_4_bits_st_dep_mask},
     {ldq_3_bits_st_dep_mask},
     {ldq_2_bits_st_dep_mask},
     {ldq_1_bits_st_dep_mask},
     {ldq_0_bits_st_dep_mask}};	// lsu.scala:210:16, :264:49
  reg  [3:0]        ldq_retry_idx;	// lsu.scala:415:30
  reg  [3:0]        stq_retry_idx;	// lsu.scala:422:30
  reg  [3:0]        ldq_wakeup_idx;	// lsu.scala:430:31
  wire              can_fire_load_incoming_0 =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_ctrl_is_load;	// lsu.scala:441:63
  wire              _can_fire_sta_incoming_T =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_ctrl_is_sta;	// lsu.scala:444:63
  wire [15:0][6:0]  _GEN_108 =
    {{ldq_15_bits_uop_uopc},
     {ldq_14_bits_uop_uopc},
     {ldq_13_bits_uop_uopc},
     {ldq_12_bits_uop_uopc},
     {ldq_11_bits_uop_uopc},
     {ldq_10_bits_uop_uopc},
     {ldq_9_bits_uop_uopc},
     {ldq_8_bits_uop_uopc},
     {ldq_7_bits_uop_uopc},
     {ldq_6_bits_uop_uopc},
     {ldq_5_bits_uop_uopc},
     {ldq_4_bits_uop_uopc},
     {ldq_3_bits_uop_uopc},
     {ldq_2_bits_uop_uopc},
     {ldq_1_bits_uop_uopc},
     {ldq_0_bits_uop_uopc}};	// lsu.scala:210:16, :465:79
  wire [15:0][31:0] _GEN_109 =
    {{ldq_15_bits_uop_inst},
     {ldq_14_bits_uop_inst},
     {ldq_13_bits_uop_inst},
     {ldq_12_bits_uop_inst},
     {ldq_11_bits_uop_inst},
     {ldq_10_bits_uop_inst},
     {ldq_9_bits_uop_inst},
     {ldq_8_bits_uop_inst},
     {ldq_7_bits_uop_inst},
     {ldq_6_bits_uop_inst},
     {ldq_5_bits_uop_inst},
     {ldq_4_bits_uop_inst},
     {ldq_3_bits_uop_inst},
     {ldq_2_bits_uop_inst},
     {ldq_1_bits_uop_inst},
     {ldq_0_bits_uop_inst}};	// lsu.scala:210:16, :465:79
  wire [15:0][31:0] _GEN_110 =
    {{ldq_15_bits_uop_debug_inst},
     {ldq_14_bits_uop_debug_inst},
     {ldq_13_bits_uop_debug_inst},
     {ldq_12_bits_uop_debug_inst},
     {ldq_11_bits_uop_debug_inst},
     {ldq_10_bits_uop_debug_inst},
     {ldq_9_bits_uop_debug_inst},
     {ldq_8_bits_uop_debug_inst},
     {ldq_7_bits_uop_debug_inst},
     {ldq_6_bits_uop_debug_inst},
     {ldq_5_bits_uop_debug_inst},
     {ldq_4_bits_uop_debug_inst},
     {ldq_3_bits_uop_debug_inst},
     {ldq_2_bits_uop_debug_inst},
     {ldq_1_bits_uop_debug_inst},
     {ldq_0_bits_uop_debug_inst}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_111 =
    {{ldq_15_bits_uop_is_rvc},
     {ldq_14_bits_uop_is_rvc},
     {ldq_13_bits_uop_is_rvc},
     {ldq_12_bits_uop_is_rvc},
     {ldq_11_bits_uop_is_rvc},
     {ldq_10_bits_uop_is_rvc},
     {ldq_9_bits_uop_is_rvc},
     {ldq_8_bits_uop_is_rvc},
     {ldq_7_bits_uop_is_rvc},
     {ldq_6_bits_uop_is_rvc},
     {ldq_5_bits_uop_is_rvc},
     {ldq_4_bits_uop_is_rvc},
     {ldq_3_bits_uop_is_rvc},
     {ldq_2_bits_uop_is_rvc},
     {ldq_1_bits_uop_is_rvc},
     {ldq_0_bits_uop_is_rvc}};	// lsu.scala:210:16, :465:79
  wire [15:0][39:0] _GEN_112 =
    {{ldq_15_bits_uop_debug_pc},
     {ldq_14_bits_uop_debug_pc},
     {ldq_13_bits_uop_debug_pc},
     {ldq_12_bits_uop_debug_pc},
     {ldq_11_bits_uop_debug_pc},
     {ldq_10_bits_uop_debug_pc},
     {ldq_9_bits_uop_debug_pc},
     {ldq_8_bits_uop_debug_pc},
     {ldq_7_bits_uop_debug_pc},
     {ldq_6_bits_uop_debug_pc},
     {ldq_5_bits_uop_debug_pc},
     {ldq_4_bits_uop_debug_pc},
     {ldq_3_bits_uop_debug_pc},
     {ldq_2_bits_uop_debug_pc},
     {ldq_1_bits_uop_debug_pc},
     {ldq_0_bits_uop_debug_pc}};	// lsu.scala:210:16, :465:79
  wire [15:0][2:0]  _GEN_113 =
    {{ldq_15_bits_uop_iq_type},
     {ldq_14_bits_uop_iq_type},
     {ldq_13_bits_uop_iq_type},
     {ldq_12_bits_uop_iq_type},
     {ldq_11_bits_uop_iq_type},
     {ldq_10_bits_uop_iq_type},
     {ldq_9_bits_uop_iq_type},
     {ldq_8_bits_uop_iq_type},
     {ldq_7_bits_uop_iq_type},
     {ldq_6_bits_uop_iq_type},
     {ldq_5_bits_uop_iq_type},
     {ldq_4_bits_uop_iq_type},
     {ldq_3_bits_uop_iq_type},
     {ldq_2_bits_uop_iq_type},
     {ldq_1_bits_uop_iq_type},
     {ldq_0_bits_uop_iq_type}};	// lsu.scala:210:16, :465:79
  wire [15:0][9:0]  _GEN_114 =
    {{ldq_15_bits_uop_fu_code},
     {ldq_14_bits_uop_fu_code},
     {ldq_13_bits_uop_fu_code},
     {ldq_12_bits_uop_fu_code},
     {ldq_11_bits_uop_fu_code},
     {ldq_10_bits_uop_fu_code},
     {ldq_9_bits_uop_fu_code},
     {ldq_8_bits_uop_fu_code},
     {ldq_7_bits_uop_fu_code},
     {ldq_6_bits_uop_fu_code},
     {ldq_5_bits_uop_fu_code},
     {ldq_4_bits_uop_fu_code},
     {ldq_3_bits_uop_fu_code},
     {ldq_2_bits_uop_fu_code},
     {ldq_1_bits_uop_fu_code},
     {ldq_0_bits_uop_fu_code}};	// lsu.scala:210:16, :465:79
  wire [15:0][3:0]  _GEN_115 =
    {{ldq_15_bits_uop_ctrl_br_type},
     {ldq_14_bits_uop_ctrl_br_type},
     {ldq_13_bits_uop_ctrl_br_type},
     {ldq_12_bits_uop_ctrl_br_type},
     {ldq_11_bits_uop_ctrl_br_type},
     {ldq_10_bits_uop_ctrl_br_type},
     {ldq_9_bits_uop_ctrl_br_type},
     {ldq_8_bits_uop_ctrl_br_type},
     {ldq_7_bits_uop_ctrl_br_type},
     {ldq_6_bits_uop_ctrl_br_type},
     {ldq_5_bits_uop_ctrl_br_type},
     {ldq_4_bits_uop_ctrl_br_type},
     {ldq_3_bits_uop_ctrl_br_type},
     {ldq_2_bits_uop_ctrl_br_type},
     {ldq_1_bits_uop_ctrl_br_type},
     {ldq_0_bits_uop_ctrl_br_type}};	// lsu.scala:210:16, :465:79
  wire [15:0][1:0]  _GEN_116 =
    {{ldq_15_bits_uop_ctrl_op1_sel},
     {ldq_14_bits_uop_ctrl_op1_sel},
     {ldq_13_bits_uop_ctrl_op1_sel},
     {ldq_12_bits_uop_ctrl_op1_sel},
     {ldq_11_bits_uop_ctrl_op1_sel},
     {ldq_10_bits_uop_ctrl_op1_sel},
     {ldq_9_bits_uop_ctrl_op1_sel},
     {ldq_8_bits_uop_ctrl_op1_sel},
     {ldq_7_bits_uop_ctrl_op1_sel},
     {ldq_6_bits_uop_ctrl_op1_sel},
     {ldq_5_bits_uop_ctrl_op1_sel},
     {ldq_4_bits_uop_ctrl_op1_sel},
     {ldq_3_bits_uop_ctrl_op1_sel},
     {ldq_2_bits_uop_ctrl_op1_sel},
     {ldq_1_bits_uop_ctrl_op1_sel},
     {ldq_0_bits_uop_ctrl_op1_sel}};	// lsu.scala:210:16, :465:79
  wire [15:0][2:0]  _GEN_117 =
    {{ldq_15_bits_uop_ctrl_op2_sel},
     {ldq_14_bits_uop_ctrl_op2_sel},
     {ldq_13_bits_uop_ctrl_op2_sel},
     {ldq_12_bits_uop_ctrl_op2_sel},
     {ldq_11_bits_uop_ctrl_op2_sel},
     {ldq_10_bits_uop_ctrl_op2_sel},
     {ldq_9_bits_uop_ctrl_op2_sel},
     {ldq_8_bits_uop_ctrl_op2_sel},
     {ldq_7_bits_uop_ctrl_op2_sel},
     {ldq_6_bits_uop_ctrl_op2_sel},
     {ldq_5_bits_uop_ctrl_op2_sel},
     {ldq_4_bits_uop_ctrl_op2_sel},
     {ldq_3_bits_uop_ctrl_op2_sel},
     {ldq_2_bits_uop_ctrl_op2_sel},
     {ldq_1_bits_uop_ctrl_op2_sel},
     {ldq_0_bits_uop_ctrl_op2_sel}};	// lsu.scala:210:16, :465:79
  wire [15:0][2:0]  _GEN_118 =
    {{ldq_15_bits_uop_ctrl_imm_sel},
     {ldq_14_bits_uop_ctrl_imm_sel},
     {ldq_13_bits_uop_ctrl_imm_sel},
     {ldq_12_bits_uop_ctrl_imm_sel},
     {ldq_11_bits_uop_ctrl_imm_sel},
     {ldq_10_bits_uop_ctrl_imm_sel},
     {ldq_9_bits_uop_ctrl_imm_sel},
     {ldq_8_bits_uop_ctrl_imm_sel},
     {ldq_7_bits_uop_ctrl_imm_sel},
     {ldq_6_bits_uop_ctrl_imm_sel},
     {ldq_5_bits_uop_ctrl_imm_sel},
     {ldq_4_bits_uop_ctrl_imm_sel},
     {ldq_3_bits_uop_ctrl_imm_sel},
     {ldq_2_bits_uop_ctrl_imm_sel},
     {ldq_1_bits_uop_ctrl_imm_sel},
     {ldq_0_bits_uop_ctrl_imm_sel}};	// lsu.scala:210:16, :465:79
  wire [15:0][3:0]  _GEN_119 =
    {{ldq_15_bits_uop_ctrl_op_fcn},
     {ldq_14_bits_uop_ctrl_op_fcn},
     {ldq_13_bits_uop_ctrl_op_fcn},
     {ldq_12_bits_uop_ctrl_op_fcn},
     {ldq_11_bits_uop_ctrl_op_fcn},
     {ldq_10_bits_uop_ctrl_op_fcn},
     {ldq_9_bits_uop_ctrl_op_fcn},
     {ldq_8_bits_uop_ctrl_op_fcn},
     {ldq_7_bits_uop_ctrl_op_fcn},
     {ldq_6_bits_uop_ctrl_op_fcn},
     {ldq_5_bits_uop_ctrl_op_fcn},
     {ldq_4_bits_uop_ctrl_op_fcn},
     {ldq_3_bits_uop_ctrl_op_fcn},
     {ldq_2_bits_uop_ctrl_op_fcn},
     {ldq_1_bits_uop_ctrl_op_fcn},
     {ldq_0_bits_uop_ctrl_op_fcn}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_120 =
    {{ldq_15_bits_uop_ctrl_fcn_dw},
     {ldq_14_bits_uop_ctrl_fcn_dw},
     {ldq_13_bits_uop_ctrl_fcn_dw},
     {ldq_12_bits_uop_ctrl_fcn_dw},
     {ldq_11_bits_uop_ctrl_fcn_dw},
     {ldq_10_bits_uop_ctrl_fcn_dw},
     {ldq_9_bits_uop_ctrl_fcn_dw},
     {ldq_8_bits_uop_ctrl_fcn_dw},
     {ldq_7_bits_uop_ctrl_fcn_dw},
     {ldq_6_bits_uop_ctrl_fcn_dw},
     {ldq_5_bits_uop_ctrl_fcn_dw},
     {ldq_4_bits_uop_ctrl_fcn_dw},
     {ldq_3_bits_uop_ctrl_fcn_dw},
     {ldq_2_bits_uop_ctrl_fcn_dw},
     {ldq_1_bits_uop_ctrl_fcn_dw},
     {ldq_0_bits_uop_ctrl_fcn_dw}};	// lsu.scala:210:16, :465:79
  wire [15:0][2:0]  _GEN_121 =
    {{ldq_15_bits_uop_ctrl_csr_cmd},
     {ldq_14_bits_uop_ctrl_csr_cmd},
     {ldq_13_bits_uop_ctrl_csr_cmd},
     {ldq_12_bits_uop_ctrl_csr_cmd},
     {ldq_11_bits_uop_ctrl_csr_cmd},
     {ldq_10_bits_uop_ctrl_csr_cmd},
     {ldq_9_bits_uop_ctrl_csr_cmd},
     {ldq_8_bits_uop_ctrl_csr_cmd},
     {ldq_7_bits_uop_ctrl_csr_cmd},
     {ldq_6_bits_uop_ctrl_csr_cmd},
     {ldq_5_bits_uop_ctrl_csr_cmd},
     {ldq_4_bits_uop_ctrl_csr_cmd},
     {ldq_3_bits_uop_ctrl_csr_cmd},
     {ldq_2_bits_uop_ctrl_csr_cmd},
     {ldq_1_bits_uop_ctrl_csr_cmd},
     {ldq_0_bits_uop_ctrl_csr_cmd}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_122 =
    {{ldq_15_bits_uop_ctrl_is_load},
     {ldq_14_bits_uop_ctrl_is_load},
     {ldq_13_bits_uop_ctrl_is_load},
     {ldq_12_bits_uop_ctrl_is_load},
     {ldq_11_bits_uop_ctrl_is_load},
     {ldq_10_bits_uop_ctrl_is_load},
     {ldq_9_bits_uop_ctrl_is_load},
     {ldq_8_bits_uop_ctrl_is_load},
     {ldq_7_bits_uop_ctrl_is_load},
     {ldq_6_bits_uop_ctrl_is_load},
     {ldq_5_bits_uop_ctrl_is_load},
     {ldq_4_bits_uop_ctrl_is_load},
     {ldq_3_bits_uop_ctrl_is_load},
     {ldq_2_bits_uop_ctrl_is_load},
     {ldq_1_bits_uop_ctrl_is_load},
     {ldq_0_bits_uop_ctrl_is_load}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_123 =
    {{ldq_15_bits_uop_ctrl_is_sta},
     {ldq_14_bits_uop_ctrl_is_sta},
     {ldq_13_bits_uop_ctrl_is_sta},
     {ldq_12_bits_uop_ctrl_is_sta},
     {ldq_11_bits_uop_ctrl_is_sta},
     {ldq_10_bits_uop_ctrl_is_sta},
     {ldq_9_bits_uop_ctrl_is_sta},
     {ldq_8_bits_uop_ctrl_is_sta},
     {ldq_7_bits_uop_ctrl_is_sta},
     {ldq_6_bits_uop_ctrl_is_sta},
     {ldq_5_bits_uop_ctrl_is_sta},
     {ldq_4_bits_uop_ctrl_is_sta},
     {ldq_3_bits_uop_ctrl_is_sta},
     {ldq_2_bits_uop_ctrl_is_sta},
     {ldq_1_bits_uop_ctrl_is_sta},
     {ldq_0_bits_uop_ctrl_is_sta}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_124 =
    {{ldq_15_bits_uop_ctrl_is_std},
     {ldq_14_bits_uop_ctrl_is_std},
     {ldq_13_bits_uop_ctrl_is_std},
     {ldq_12_bits_uop_ctrl_is_std},
     {ldq_11_bits_uop_ctrl_is_std},
     {ldq_10_bits_uop_ctrl_is_std},
     {ldq_9_bits_uop_ctrl_is_std},
     {ldq_8_bits_uop_ctrl_is_std},
     {ldq_7_bits_uop_ctrl_is_std},
     {ldq_6_bits_uop_ctrl_is_std},
     {ldq_5_bits_uop_ctrl_is_std},
     {ldq_4_bits_uop_ctrl_is_std},
     {ldq_3_bits_uop_ctrl_is_std},
     {ldq_2_bits_uop_ctrl_is_std},
     {ldq_1_bits_uop_ctrl_is_std},
     {ldq_0_bits_uop_ctrl_is_std}};	// lsu.scala:210:16, :465:79
  wire [15:0][1:0]  _GEN_125 =
    {{ldq_15_bits_uop_iw_state},
     {ldq_14_bits_uop_iw_state},
     {ldq_13_bits_uop_iw_state},
     {ldq_12_bits_uop_iw_state},
     {ldq_11_bits_uop_iw_state},
     {ldq_10_bits_uop_iw_state},
     {ldq_9_bits_uop_iw_state},
     {ldq_8_bits_uop_iw_state},
     {ldq_7_bits_uop_iw_state},
     {ldq_6_bits_uop_iw_state},
     {ldq_5_bits_uop_iw_state},
     {ldq_4_bits_uop_iw_state},
     {ldq_3_bits_uop_iw_state},
     {ldq_2_bits_uop_iw_state},
     {ldq_1_bits_uop_iw_state},
     {ldq_0_bits_uop_iw_state}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_126 =
    {{ldq_15_bits_uop_iw_p1_poisoned},
     {ldq_14_bits_uop_iw_p1_poisoned},
     {ldq_13_bits_uop_iw_p1_poisoned},
     {ldq_12_bits_uop_iw_p1_poisoned},
     {ldq_11_bits_uop_iw_p1_poisoned},
     {ldq_10_bits_uop_iw_p1_poisoned},
     {ldq_9_bits_uop_iw_p1_poisoned},
     {ldq_8_bits_uop_iw_p1_poisoned},
     {ldq_7_bits_uop_iw_p1_poisoned},
     {ldq_6_bits_uop_iw_p1_poisoned},
     {ldq_5_bits_uop_iw_p1_poisoned},
     {ldq_4_bits_uop_iw_p1_poisoned},
     {ldq_3_bits_uop_iw_p1_poisoned},
     {ldq_2_bits_uop_iw_p1_poisoned},
     {ldq_1_bits_uop_iw_p1_poisoned},
     {ldq_0_bits_uop_iw_p1_poisoned}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_127 =
    {{ldq_15_bits_uop_iw_p2_poisoned},
     {ldq_14_bits_uop_iw_p2_poisoned},
     {ldq_13_bits_uop_iw_p2_poisoned},
     {ldq_12_bits_uop_iw_p2_poisoned},
     {ldq_11_bits_uop_iw_p2_poisoned},
     {ldq_10_bits_uop_iw_p2_poisoned},
     {ldq_9_bits_uop_iw_p2_poisoned},
     {ldq_8_bits_uop_iw_p2_poisoned},
     {ldq_7_bits_uop_iw_p2_poisoned},
     {ldq_6_bits_uop_iw_p2_poisoned},
     {ldq_5_bits_uop_iw_p2_poisoned},
     {ldq_4_bits_uop_iw_p2_poisoned},
     {ldq_3_bits_uop_iw_p2_poisoned},
     {ldq_2_bits_uop_iw_p2_poisoned},
     {ldq_1_bits_uop_iw_p2_poisoned},
     {ldq_0_bits_uop_iw_p2_poisoned}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_128 =
    {{ldq_15_bits_uop_is_br},
     {ldq_14_bits_uop_is_br},
     {ldq_13_bits_uop_is_br},
     {ldq_12_bits_uop_is_br},
     {ldq_11_bits_uop_is_br},
     {ldq_10_bits_uop_is_br},
     {ldq_9_bits_uop_is_br},
     {ldq_8_bits_uop_is_br},
     {ldq_7_bits_uop_is_br},
     {ldq_6_bits_uop_is_br},
     {ldq_5_bits_uop_is_br},
     {ldq_4_bits_uop_is_br},
     {ldq_3_bits_uop_is_br},
     {ldq_2_bits_uop_is_br},
     {ldq_1_bits_uop_is_br},
     {ldq_0_bits_uop_is_br}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_129 =
    {{ldq_15_bits_uop_is_jalr},
     {ldq_14_bits_uop_is_jalr},
     {ldq_13_bits_uop_is_jalr},
     {ldq_12_bits_uop_is_jalr},
     {ldq_11_bits_uop_is_jalr},
     {ldq_10_bits_uop_is_jalr},
     {ldq_9_bits_uop_is_jalr},
     {ldq_8_bits_uop_is_jalr},
     {ldq_7_bits_uop_is_jalr},
     {ldq_6_bits_uop_is_jalr},
     {ldq_5_bits_uop_is_jalr},
     {ldq_4_bits_uop_is_jalr},
     {ldq_3_bits_uop_is_jalr},
     {ldq_2_bits_uop_is_jalr},
     {ldq_1_bits_uop_is_jalr},
     {ldq_0_bits_uop_is_jalr}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_130 =
    {{ldq_15_bits_uop_is_jal},
     {ldq_14_bits_uop_is_jal},
     {ldq_13_bits_uop_is_jal},
     {ldq_12_bits_uop_is_jal},
     {ldq_11_bits_uop_is_jal},
     {ldq_10_bits_uop_is_jal},
     {ldq_9_bits_uop_is_jal},
     {ldq_8_bits_uop_is_jal},
     {ldq_7_bits_uop_is_jal},
     {ldq_6_bits_uop_is_jal},
     {ldq_5_bits_uop_is_jal},
     {ldq_4_bits_uop_is_jal},
     {ldq_3_bits_uop_is_jal},
     {ldq_2_bits_uop_is_jal},
     {ldq_1_bits_uop_is_jal},
     {ldq_0_bits_uop_is_jal}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_131 =
    {{ldq_15_bits_uop_is_sfb},
     {ldq_14_bits_uop_is_sfb},
     {ldq_13_bits_uop_is_sfb},
     {ldq_12_bits_uop_is_sfb},
     {ldq_11_bits_uop_is_sfb},
     {ldq_10_bits_uop_is_sfb},
     {ldq_9_bits_uop_is_sfb},
     {ldq_8_bits_uop_is_sfb},
     {ldq_7_bits_uop_is_sfb},
     {ldq_6_bits_uop_is_sfb},
     {ldq_5_bits_uop_is_sfb},
     {ldq_4_bits_uop_is_sfb},
     {ldq_3_bits_uop_is_sfb},
     {ldq_2_bits_uop_is_sfb},
     {ldq_1_bits_uop_is_sfb},
     {ldq_0_bits_uop_is_sfb}};	// lsu.scala:210:16, :465:79
  wire [11:0]       _GEN_132 = _GEN_102[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79
  wire [15:0][3:0]  _GEN_133 =
    {{ldq_15_bits_uop_br_tag},
     {ldq_14_bits_uop_br_tag},
     {ldq_13_bits_uop_br_tag},
     {ldq_12_bits_uop_br_tag},
     {ldq_11_bits_uop_br_tag},
     {ldq_10_bits_uop_br_tag},
     {ldq_9_bits_uop_br_tag},
     {ldq_8_bits_uop_br_tag},
     {ldq_7_bits_uop_br_tag},
     {ldq_6_bits_uop_br_tag},
     {ldq_5_bits_uop_br_tag},
     {ldq_4_bits_uop_br_tag},
     {ldq_3_bits_uop_br_tag},
     {ldq_2_bits_uop_br_tag},
     {ldq_1_bits_uop_br_tag},
     {ldq_0_bits_uop_br_tag}};	// lsu.scala:210:16, :465:79
  wire [15:0][4:0]  _GEN_134 =
    {{ldq_15_bits_uop_ftq_idx},
     {ldq_14_bits_uop_ftq_idx},
     {ldq_13_bits_uop_ftq_idx},
     {ldq_12_bits_uop_ftq_idx},
     {ldq_11_bits_uop_ftq_idx},
     {ldq_10_bits_uop_ftq_idx},
     {ldq_9_bits_uop_ftq_idx},
     {ldq_8_bits_uop_ftq_idx},
     {ldq_7_bits_uop_ftq_idx},
     {ldq_6_bits_uop_ftq_idx},
     {ldq_5_bits_uop_ftq_idx},
     {ldq_4_bits_uop_ftq_idx},
     {ldq_3_bits_uop_ftq_idx},
     {ldq_2_bits_uop_ftq_idx},
     {ldq_1_bits_uop_ftq_idx},
     {ldq_0_bits_uop_ftq_idx}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_135 =
    {{ldq_15_bits_uop_edge_inst},
     {ldq_14_bits_uop_edge_inst},
     {ldq_13_bits_uop_edge_inst},
     {ldq_12_bits_uop_edge_inst},
     {ldq_11_bits_uop_edge_inst},
     {ldq_10_bits_uop_edge_inst},
     {ldq_9_bits_uop_edge_inst},
     {ldq_8_bits_uop_edge_inst},
     {ldq_7_bits_uop_edge_inst},
     {ldq_6_bits_uop_edge_inst},
     {ldq_5_bits_uop_edge_inst},
     {ldq_4_bits_uop_edge_inst},
     {ldq_3_bits_uop_edge_inst},
     {ldq_2_bits_uop_edge_inst},
     {ldq_1_bits_uop_edge_inst},
     {ldq_0_bits_uop_edge_inst}};	// lsu.scala:210:16, :465:79
  wire [15:0][5:0]  _GEN_136 =
    {{ldq_15_bits_uop_pc_lob},
     {ldq_14_bits_uop_pc_lob},
     {ldq_13_bits_uop_pc_lob},
     {ldq_12_bits_uop_pc_lob},
     {ldq_11_bits_uop_pc_lob},
     {ldq_10_bits_uop_pc_lob},
     {ldq_9_bits_uop_pc_lob},
     {ldq_8_bits_uop_pc_lob},
     {ldq_7_bits_uop_pc_lob},
     {ldq_6_bits_uop_pc_lob},
     {ldq_5_bits_uop_pc_lob},
     {ldq_4_bits_uop_pc_lob},
     {ldq_3_bits_uop_pc_lob},
     {ldq_2_bits_uop_pc_lob},
     {ldq_1_bits_uop_pc_lob},
     {ldq_0_bits_uop_pc_lob}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_137 =
    {{ldq_15_bits_uop_taken},
     {ldq_14_bits_uop_taken},
     {ldq_13_bits_uop_taken},
     {ldq_12_bits_uop_taken},
     {ldq_11_bits_uop_taken},
     {ldq_10_bits_uop_taken},
     {ldq_9_bits_uop_taken},
     {ldq_8_bits_uop_taken},
     {ldq_7_bits_uop_taken},
     {ldq_6_bits_uop_taken},
     {ldq_5_bits_uop_taken},
     {ldq_4_bits_uop_taken},
     {ldq_3_bits_uop_taken},
     {ldq_2_bits_uop_taken},
     {ldq_1_bits_uop_taken},
     {ldq_0_bits_uop_taken}};	// lsu.scala:210:16, :465:79
  wire [15:0][19:0] _GEN_138 =
    {{ldq_15_bits_uop_imm_packed},
     {ldq_14_bits_uop_imm_packed},
     {ldq_13_bits_uop_imm_packed},
     {ldq_12_bits_uop_imm_packed},
     {ldq_11_bits_uop_imm_packed},
     {ldq_10_bits_uop_imm_packed},
     {ldq_9_bits_uop_imm_packed},
     {ldq_8_bits_uop_imm_packed},
     {ldq_7_bits_uop_imm_packed},
     {ldq_6_bits_uop_imm_packed},
     {ldq_5_bits_uop_imm_packed},
     {ldq_4_bits_uop_imm_packed},
     {ldq_3_bits_uop_imm_packed},
     {ldq_2_bits_uop_imm_packed},
     {ldq_1_bits_uop_imm_packed},
     {ldq_0_bits_uop_imm_packed}};	// lsu.scala:210:16, :465:79
  wire [15:0][11:0] _GEN_139 =
    {{ldq_15_bits_uop_csr_addr},
     {ldq_14_bits_uop_csr_addr},
     {ldq_13_bits_uop_csr_addr},
     {ldq_12_bits_uop_csr_addr},
     {ldq_11_bits_uop_csr_addr},
     {ldq_10_bits_uop_csr_addr},
     {ldq_9_bits_uop_csr_addr},
     {ldq_8_bits_uop_csr_addr},
     {ldq_7_bits_uop_csr_addr},
     {ldq_6_bits_uop_csr_addr},
     {ldq_5_bits_uop_csr_addr},
     {ldq_4_bits_uop_csr_addr},
     {ldq_3_bits_uop_csr_addr},
     {ldq_2_bits_uop_csr_addr},
     {ldq_1_bits_uop_csr_addr},
     {ldq_0_bits_uop_csr_addr}};	// lsu.scala:210:16, :465:79
  wire [15:0][5:0]  _GEN_140 =
    {{ldq_15_bits_uop_rob_idx},
     {ldq_14_bits_uop_rob_idx},
     {ldq_13_bits_uop_rob_idx},
     {ldq_12_bits_uop_rob_idx},
     {ldq_11_bits_uop_rob_idx},
     {ldq_10_bits_uop_rob_idx},
     {ldq_9_bits_uop_rob_idx},
     {ldq_8_bits_uop_rob_idx},
     {ldq_7_bits_uop_rob_idx},
     {ldq_6_bits_uop_rob_idx},
     {ldq_5_bits_uop_rob_idx},
     {ldq_4_bits_uop_rob_idx},
     {ldq_3_bits_uop_rob_idx},
     {ldq_2_bits_uop_rob_idx},
     {ldq_1_bits_uop_rob_idx},
     {ldq_0_bits_uop_rob_idx}};	// lsu.scala:210:16, :465:79
  wire [5:0]        _GEN_141 = _GEN_140[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [15:0][3:0]  _GEN_142 =
    {{ldq_15_bits_uop_ldq_idx},
     {ldq_14_bits_uop_ldq_idx},
     {ldq_13_bits_uop_ldq_idx},
     {ldq_12_bits_uop_ldq_idx},
     {ldq_11_bits_uop_ldq_idx},
     {ldq_10_bits_uop_ldq_idx},
     {ldq_9_bits_uop_ldq_idx},
     {ldq_8_bits_uop_ldq_idx},
     {ldq_7_bits_uop_ldq_idx},
     {ldq_6_bits_uop_ldq_idx},
     {ldq_5_bits_uop_ldq_idx},
     {ldq_4_bits_uop_ldq_idx},
     {ldq_3_bits_uop_ldq_idx},
     {ldq_2_bits_uop_ldq_idx},
     {ldq_1_bits_uop_ldq_idx},
     {ldq_0_bits_uop_ldq_idx}};	// lsu.scala:210:16, :465:79
  wire [3:0]        _GEN_143 = _GEN_142[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [3:0]        mem_ldq_retry_e_out_bits_uop_stq_idx = _GEN_103[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79
  wire [15:0][1:0]  _GEN_144 =
    {{ldq_15_bits_uop_rxq_idx},
     {ldq_14_bits_uop_rxq_idx},
     {ldq_13_bits_uop_rxq_idx},
     {ldq_12_bits_uop_rxq_idx},
     {ldq_11_bits_uop_rxq_idx},
     {ldq_10_bits_uop_rxq_idx},
     {ldq_9_bits_uop_rxq_idx},
     {ldq_8_bits_uop_rxq_idx},
     {ldq_7_bits_uop_rxq_idx},
     {ldq_6_bits_uop_rxq_idx},
     {ldq_5_bits_uop_rxq_idx},
     {ldq_4_bits_uop_rxq_idx},
     {ldq_3_bits_uop_rxq_idx},
     {ldq_2_bits_uop_rxq_idx},
     {ldq_1_bits_uop_rxq_idx},
     {ldq_0_bits_uop_rxq_idx}};	// lsu.scala:210:16, :465:79
  wire [15:0][6:0]  _GEN_145 =
    {{ldq_15_bits_uop_pdst},
     {ldq_14_bits_uop_pdst},
     {ldq_13_bits_uop_pdst},
     {ldq_12_bits_uop_pdst},
     {ldq_11_bits_uop_pdst},
     {ldq_10_bits_uop_pdst},
     {ldq_9_bits_uop_pdst},
     {ldq_8_bits_uop_pdst},
     {ldq_7_bits_uop_pdst},
     {ldq_6_bits_uop_pdst},
     {ldq_5_bits_uop_pdst},
     {ldq_4_bits_uop_pdst},
     {ldq_3_bits_uop_pdst},
     {ldq_2_bits_uop_pdst},
     {ldq_1_bits_uop_pdst},
     {ldq_0_bits_uop_pdst}};	// lsu.scala:210:16, :465:79
  wire [6:0]        _GEN_146 = _GEN_145[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [15:0][6:0]  _GEN_147 =
    {{ldq_15_bits_uop_prs1},
     {ldq_14_bits_uop_prs1},
     {ldq_13_bits_uop_prs1},
     {ldq_12_bits_uop_prs1},
     {ldq_11_bits_uop_prs1},
     {ldq_10_bits_uop_prs1},
     {ldq_9_bits_uop_prs1},
     {ldq_8_bits_uop_prs1},
     {ldq_7_bits_uop_prs1},
     {ldq_6_bits_uop_prs1},
     {ldq_5_bits_uop_prs1},
     {ldq_4_bits_uop_prs1},
     {ldq_3_bits_uop_prs1},
     {ldq_2_bits_uop_prs1},
     {ldq_1_bits_uop_prs1},
     {ldq_0_bits_uop_prs1}};	// lsu.scala:210:16, :465:79
  wire [15:0][6:0]  _GEN_148 =
    {{ldq_15_bits_uop_prs2},
     {ldq_14_bits_uop_prs2},
     {ldq_13_bits_uop_prs2},
     {ldq_12_bits_uop_prs2},
     {ldq_11_bits_uop_prs2},
     {ldq_10_bits_uop_prs2},
     {ldq_9_bits_uop_prs2},
     {ldq_8_bits_uop_prs2},
     {ldq_7_bits_uop_prs2},
     {ldq_6_bits_uop_prs2},
     {ldq_5_bits_uop_prs2},
     {ldq_4_bits_uop_prs2},
     {ldq_3_bits_uop_prs2},
     {ldq_2_bits_uop_prs2},
     {ldq_1_bits_uop_prs2},
     {ldq_0_bits_uop_prs2}};	// lsu.scala:210:16, :465:79
  wire [15:0][6:0]  _GEN_149 =
    {{ldq_15_bits_uop_prs3},
     {ldq_14_bits_uop_prs3},
     {ldq_13_bits_uop_prs3},
     {ldq_12_bits_uop_prs3},
     {ldq_11_bits_uop_prs3},
     {ldq_10_bits_uop_prs3},
     {ldq_9_bits_uop_prs3},
     {ldq_8_bits_uop_prs3},
     {ldq_7_bits_uop_prs3},
     {ldq_6_bits_uop_prs3},
     {ldq_5_bits_uop_prs3},
     {ldq_4_bits_uop_prs3},
     {ldq_3_bits_uop_prs3},
     {ldq_2_bits_uop_prs3},
     {ldq_1_bits_uop_prs3},
     {ldq_0_bits_uop_prs3}};	// lsu.scala:210:16, :465:79
  wire [15:0][4:0]  _GEN_150 =
    {{ldq_15_bits_uop_ppred},
     {ldq_14_bits_uop_ppred},
     {ldq_13_bits_uop_ppred},
     {ldq_12_bits_uop_ppred},
     {ldq_11_bits_uop_ppred},
     {ldq_10_bits_uop_ppred},
     {ldq_9_bits_uop_ppred},
     {ldq_8_bits_uop_ppred},
     {ldq_7_bits_uop_ppred},
     {ldq_6_bits_uop_ppred},
     {ldq_5_bits_uop_ppred},
     {ldq_4_bits_uop_ppred},
     {ldq_3_bits_uop_ppred},
     {ldq_2_bits_uop_ppred},
     {ldq_1_bits_uop_ppred},
     {ldq_0_bits_uop_ppred}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_151 =
    {{ldq_15_bits_uop_prs1_busy},
     {ldq_14_bits_uop_prs1_busy},
     {ldq_13_bits_uop_prs1_busy},
     {ldq_12_bits_uop_prs1_busy},
     {ldq_11_bits_uop_prs1_busy},
     {ldq_10_bits_uop_prs1_busy},
     {ldq_9_bits_uop_prs1_busy},
     {ldq_8_bits_uop_prs1_busy},
     {ldq_7_bits_uop_prs1_busy},
     {ldq_6_bits_uop_prs1_busy},
     {ldq_5_bits_uop_prs1_busy},
     {ldq_4_bits_uop_prs1_busy},
     {ldq_3_bits_uop_prs1_busy},
     {ldq_2_bits_uop_prs1_busy},
     {ldq_1_bits_uop_prs1_busy},
     {ldq_0_bits_uop_prs1_busy}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_152 =
    {{ldq_15_bits_uop_prs2_busy},
     {ldq_14_bits_uop_prs2_busy},
     {ldq_13_bits_uop_prs2_busy},
     {ldq_12_bits_uop_prs2_busy},
     {ldq_11_bits_uop_prs2_busy},
     {ldq_10_bits_uop_prs2_busy},
     {ldq_9_bits_uop_prs2_busy},
     {ldq_8_bits_uop_prs2_busy},
     {ldq_7_bits_uop_prs2_busy},
     {ldq_6_bits_uop_prs2_busy},
     {ldq_5_bits_uop_prs2_busy},
     {ldq_4_bits_uop_prs2_busy},
     {ldq_3_bits_uop_prs2_busy},
     {ldq_2_bits_uop_prs2_busy},
     {ldq_1_bits_uop_prs2_busy},
     {ldq_0_bits_uop_prs2_busy}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_153 =
    {{ldq_15_bits_uop_prs3_busy},
     {ldq_14_bits_uop_prs3_busy},
     {ldq_13_bits_uop_prs3_busy},
     {ldq_12_bits_uop_prs3_busy},
     {ldq_11_bits_uop_prs3_busy},
     {ldq_10_bits_uop_prs3_busy},
     {ldq_9_bits_uop_prs3_busy},
     {ldq_8_bits_uop_prs3_busy},
     {ldq_7_bits_uop_prs3_busy},
     {ldq_6_bits_uop_prs3_busy},
     {ldq_5_bits_uop_prs3_busy},
     {ldq_4_bits_uop_prs3_busy},
     {ldq_3_bits_uop_prs3_busy},
     {ldq_2_bits_uop_prs3_busy},
     {ldq_1_bits_uop_prs3_busy},
     {ldq_0_bits_uop_prs3_busy}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_154 =
    {{ldq_15_bits_uop_ppred_busy},
     {ldq_14_bits_uop_ppred_busy},
     {ldq_13_bits_uop_ppred_busy},
     {ldq_12_bits_uop_ppred_busy},
     {ldq_11_bits_uop_ppred_busy},
     {ldq_10_bits_uop_ppred_busy},
     {ldq_9_bits_uop_ppred_busy},
     {ldq_8_bits_uop_ppred_busy},
     {ldq_7_bits_uop_ppred_busy},
     {ldq_6_bits_uop_ppred_busy},
     {ldq_5_bits_uop_ppred_busy},
     {ldq_4_bits_uop_ppred_busy},
     {ldq_3_bits_uop_ppred_busy},
     {ldq_2_bits_uop_ppred_busy},
     {ldq_1_bits_uop_ppred_busy},
     {ldq_0_bits_uop_ppred_busy}};	// lsu.scala:210:16, :465:79
  wire [15:0][6:0]  _GEN_155 =
    {{ldq_15_bits_uop_stale_pdst},
     {ldq_14_bits_uop_stale_pdst},
     {ldq_13_bits_uop_stale_pdst},
     {ldq_12_bits_uop_stale_pdst},
     {ldq_11_bits_uop_stale_pdst},
     {ldq_10_bits_uop_stale_pdst},
     {ldq_9_bits_uop_stale_pdst},
     {ldq_8_bits_uop_stale_pdst},
     {ldq_7_bits_uop_stale_pdst},
     {ldq_6_bits_uop_stale_pdst},
     {ldq_5_bits_uop_stale_pdst},
     {ldq_4_bits_uop_stale_pdst},
     {ldq_3_bits_uop_stale_pdst},
     {ldq_2_bits_uop_stale_pdst},
     {ldq_1_bits_uop_stale_pdst},
     {ldq_0_bits_uop_stale_pdst}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_156 =
    {{ldq_15_bits_uop_exception},
     {ldq_14_bits_uop_exception},
     {ldq_13_bits_uop_exception},
     {ldq_12_bits_uop_exception},
     {ldq_11_bits_uop_exception},
     {ldq_10_bits_uop_exception},
     {ldq_9_bits_uop_exception},
     {ldq_8_bits_uop_exception},
     {ldq_7_bits_uop_exception},
     {ldq_6_bits_uop_exception},
     {ldq_5_bits_uop_exception},
     {ldq_4_bits_uop_exception},
     {ldq_3_bits_uop_exception},
     {ldq_2_bits_uop_exception},
     {ldq_1_bits_uop_exception},
     {ldq_0_bits_uop_exception}};	// lsu.scala:210:16, :465:79
  wire [15:0][63:0] _GEN_157 =
    {{ldq_15_bits_uop_exc_cause},
     {ldq_14_bits_uop_exc_cause},
     {ldq_13_bits_uop_exc_cause},
     {ldq_12_bits_uop_exc_cause},
     {ldq_11_bits_uop_exc_cause},
     {ldq_10_bits_uop_exc_cause},
     {ldq_9_bits_uop_exc_cause},
     {ldq_8_bits_uop_exc_cause},
     {ldq_7_bits_uop_exc_cause},
     {ldq_6_bits_uop_exc_cause},
     {ldq_5_bits_uop_exc_cause},
     {ldq_4_bits_uop_exc_cause},
     {ldq_3_bits_uop_exc_cause},
     {ldq_2_bits_uop_exc_cause},
     {ldq_1_bits_uop_exc_cause},
     {ldq_0_bits_uop_exc_cause}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_158 =
    {{ldq_15_bits_uop_bypassable},
     {ldq_14_bits_uop_bypassable},
     {ldq_13_bits_uop_bypassable},
     {ldq_12_bits_uop_bypassable},
     {ldq_11_bits_uop_bypassable},
     {ldq_10_bits_uop_bypassable},
     {ldq_9_bits_uop_bypassable},
     {ldq_8_bits_uop_bypassable},
     {ldq_7_bits_uop_bypassable},
     {ldq_6_bits_uop_bypassable},
     {ldq_5_bits_uop_bypassable},
     {ldq_4_bits_uop_bypassable},
     {ldq_3_bits_uop_bypassable},
     {ldq_2_bits_uop_bypassable},
     {ldq_1_bits_uop_bypassable},
     {ldq_0_bits_uop_bypassable}};	// lsu.scala:210:16, :465:79
  wire [15:0][4:0]  _GEN_159 =
    {{ldq_15_bits_uop_mem_cmd},
     {ldq_14_bits_uop_mem_cmd},
     {ldq_13_bits_uop_mem_cmd},
     {ldq_12_bits_uop_mem_cmd},
     {ldq_11_bits_uop_mem_cmd},
     {ldq_10_bits_uop_mem_cmd},
     {ldq_9_bits_uop_mem_cmd},
     {ldq_8_bits_uop_mem_cmd},
     {ldq_7_bits_uop_mem_cmd},
     {ldq_6_bits_uop_mem_cmd},
     {ldq_5_bits_uop_mem_cmd},
     {ldq_4_bits_uop_mem_cmd},
     {ldq_3_bits_uop_mem_cmd},
     {ldq_2_bits_uop_mem_cmd},
     {ldq_1_bits_uop_mem_cmd},
     {ldq_0_bits_uop_mem_cmd}};	// lsu.scala:210:16, :465:79
  wire [1:0]        mem_ldq_retry_e_out_bits_uop_mem_size = _GEN_104[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79
  wire [15:0]       _GEN_160 =
    {{ldq_15_bits_uop_mem_signed},
     {ldq_14_bits_uop_mem_signed},
     {ldq_13_bits_uop_mem_signed},
     {ldq_12_bits_uop_mem_signed},
     {ldq_11_bits_uop_mem_signed},
     {ldq_10_bits_uop_mem_signed},
     {ldq_9_bits_uop_mem_signed},
     {ldq_8_bits_uop_mem_signed},
     {ldq_7_bits_uop_mem_signed},
     {ldq_6_bits_uop_mem_signed},
     {ldq_5_bits_uop_mem_signed},
     {ldq_4_bits_uop_mem_signed},
     {ldq_3_bits_uop_mem_signed},
     {ldq_2_bits_uop_mem_signed},
     {ldq_1_bits_uop_mem_signed},
     {ldq_0_bits_uop_mem_signed}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_161 =
    {{ldq_15_bits_uop_is_fence},
     {ldq_14_bits_uop_is_fence},
     {ldq_13_bits_uop_is_fence},
     {ldq_12_bits_uop_is_fence},
     {ldq_11_bits_uop_is_fence},
     {ldq_10_bits_uop_is_fence},
     {ldq_9_bits_uop_is_fence},
     {ldq_8_bits_uop_is_fence},
     {ldq_7_bits_uop_is_fence},
     {ldq_6_bits_uop_is_fence},
     {ldq_5_bits_uop_is_fence},
     {ldq_4_bits_uop_is_fence},
     {ldq_3_bits_uop_is_fence},
     {ldq_2_bits_uop_is_fence},
     {ldq_1_bits_uop_is_fence},
     {ldq_0_bits_uop_is_fence}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_162 =
    {{ldq_15_bits_uop_is_fencei},
     {ldq_14_bits_uop_is_fencei},
     {ldq_13_bits_uop_is_fencei},
     {ldq_12_bits_uop_is_fencei},
     {ldq_11_bits_uop_is_fencei},
     {ldq_10_bits_uop_is_fencei},
     {ldq_9_bits_uop_is_fencei},
     {ldq_8_bits_uop_is_fencei},
     {ldq_7_bits_uop_is_fencei},
     {ldq_6_bits_uop_is_fencei},
     {ldq_5_bits_uop_is_fencei},
     {ldq_4_bits_uop_is_fencei},
     {ldq_3_bits_uop_is_fencei},
     {ldq_2_bits_uop_is_fencei},
     {ldq_1_bits_uop_is_fencei},
     {ldq_0_bits_uop_is_fencei}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_163 =
    {{ldq_15_bits_uop_is_amo},
     {ldq_14_bits_uop_is_amo},
     {ldq_13_bits_uop_is_amo},
     {ldq_12_bits_uop_is_amo},
     {ldq_11_bits_uop_is_amo},
     {ldq_10_bits_uop_is_amo},
     {ldq_9_bits_uop_is_amo},
     {ldq_8_bits_uop_is_amo},
     {ldq_7_bits_uop_is_amo},
     {ldq_6_bits_uop_is_amo},
     {ldq_5_bits_uop_is_amo},
     {ldq_4_bits_uop_is_amo},
     {ldq_3_bits_uop_is_amo},
     {ldq_2_bits_uop_is_amo},
     {ldq_1_bits_uop_is_amo},
     {ldq_0_bits_uop_is_amo}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_164 =
    {{ldq_15_bits_uop_uses_ldq},
     {ldq_14_bits_uop_uses_ldq},
     {ldq_13_bits_uop_uses_ldq},
     {ldq_12_bits_uop_uses_ldq},
     {ldq_11_bits_uop_uses_ldq},
     {ldq_10_bits_uop_uses_ldq},
     {ldq_9_bits_uop_uses_ldq},
     {ldq_8_bits_uop_uses_ldq},
     {ldq_7_bits_uop_uses_ldq},
     {ldq_6_bits_uop_uses_ldq},
     {ldq_5_bits_uop_uses_ldq},
     {ldq_4_bits_uop_uses_ldq},
     {ldq_3_bits_uop_uses_ldq},
     {ldq_2_bits_uop_uses_ldq},
     {ldq_1_bits_uop_uses_ldq},
     {ldq_0_bits_uop_uses_ldq}};	// lsu.scala:210:16, :465:79
  wire              _GEN_165 = _GEN_164[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [15:0]       _GEN_166 =
    {{ldq_15_bits_uop_uses_stq},
     {ldq_14_bits_uop_uses_stq},
     {ldq_13_bits_uop_uses_stq},
     {ldq_12_bits_uop_uses_stq},
     {ldq_11_bits_uop_uses_stq},
     {ldq_10_bits_uop_uses_stq},
     {ldq_9_bits_uop_uses_stq},
     {ldq_8_bits_uop_uses_stq},
     {ldq_7_bits_uop_uses_stq},
     {ldq_6_bits_uop_uses_stq},
     {ldq_5_bits_uop_uses_stq},
     {ldq_4_bits_uop_uses_stq},
     {ldq_3_bits_uop_uses_stq},
     {ldq_2_bits_uop_uses_stq},
     {ldq_1_bits_uop_uses_stq},
     {ldq_0_bits_uop_uses_stq}};	// lsu.scala:210:16, :465:79
  wire              _GEN_167 = _GEN_166[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [15:0]       _GEN_168 =
    {{ldq_15_bits_uop_is_sys_pc2epc},
     {ldq_14_bits_uop_is_sys_pc2epc},
     {ldq_13_bits_uop_is_sys_pc2epc},
     {ldq_12_bits_uop_is_sys_pc2epc},
     {ldq_11_bits_uop_is_sys_pc2epc},
     {ldq_10_bits_uop_is_sys_pc2epc},
     {ldq_9_bits_uop_is_sys_pc2epc},
     {ldq_8_bits_uop_is_sys_pc2epc},
     {ldq_7_bits_uop_is_sys_pc2epc},
     {ldq_6_bits_uop_is_sys_pc2epc},
     {ldq_5_bits_uop_is_sys_pc2epc},
     {ldq_4_bits_uop_is_sys_pc2epc},
     {ldq_3_bits_uop_is_sys_pc2epc},
     {ldq_2_bits_uop_is_sys_pc2epc},
     {ldq_1_bits_uop_is_sys_pc2epc},
     {ldq_0_bits_uop_is_sys_pc2epc}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_169 =
    {{ldq_15_bits_uop_is_unique},
     {ldq_14_bits_uop_is_unique},
     {ldq_13_bits_uop_is_unique},
     {ldq_12_bits_uop_is_unique},
     {ldq_11_bits_uop_is_unique},
     {ldq_10_bits_uop_is_unique},
     {ldq_9_bits_uop_is_unique},
     {ldq_8_bits_uop_is_unique},
     {ldq_7_bits_uop_is_unique},
     {ldq_6_bits_uop_is_unique},
     {ldq_5_bits_uop_is_unique},
     {ldq_4_bits_uop_is_unique},
     {ldq_3_bits_uop_is_unique},
     {ldq_2_bits_uop_is_unique},
     {ldq_1_bits_uop_is_unique},
     {ldq_0_bits_uop_is_unique}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_170 =
    {{ldq_15_bits_uop_flush_on_commit},
     {ldq_14_bits_uop_flush_on_commit},
     {ldq_13_bits_uop_flush_on_commit},
     {ldq_12_bits_uop_flush_on_commit},
     {ldq_11_bits_uop_flush_on_commit},
     {ldq_10_bits_uop_flush_on_commit},
     {ldq_9_bits_uop_flush_on_commit},
     {ldq_8_bits_uop_flush_on_commit},
     {ldq_7_bits_uop_flush_on_commit},
     {ldq_6_bits_uop_flush_on_commit},
     {ldq_5_bits_uop_flush_on_commit},
     {ldq_4_bits_uop_flush_on_commit},
     {ldq_3_bits_uop_flush_on_commit},
     {ldq_2_bits_uop_flush_on_commit},
     {ldq_1_bits_uop_flush_on_commit},
     {ldq_0_bits_uop_flush_on_commit}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_171 =
    {{ldq_15_bits_uop_ldst_is_rs1},
     {ldq_14_bits_uop_ldst_is_rs1},
     {ldq_13_bits_uop_ldst_is_rs1},
     {ldq_12_bits_uop_ldst_is_rs1},
     {ldq_11_bits_uop_ldst_is_rs1},
     {ldq_10_bits_uop_ldst_is_rs1},
     {ldq_9_bits_uop_ldst_is_rs1},
     {ldq_8_bits_uop_ldst_is_rs1},
     {ldq_7_bits_uop_ldst_is_rs1},
     {ldq_6_bits_uop_ldst_is_rs1},
     {ldq_5_bits_uop_ldst_is_rs1},
     {ldq_4_bits_uop_ldst_is_rs1},
     {ldq_3_bits_uop_ldst_is_rs1},
     {ldq_2_bits_uop_ldst_is_rs1},
     {ldq_1_bits_uop_ldst_is_rs1},
     {ldq_0_bits_uop_ldst_is_rs1}};	// lsu.scala:210:16, :465:79
  wire [15:0][5:0]  _GEN_172 =
    {{ldq_15_bits_uop_ldst},
     {ldq_14_bits_uop_ldst},
     {ldq_13_bits_uop_ldst},
     {ldq_12_bits_uop_ldst},
     {ldq_11_bits_uop_ldst},
     {ldq_10_bits_uop_ldst},
     {ldq_9_bits_uop_ldst},
     {ldq_8_bits_uop_ldst},
     {ldq_7_bits_uop_ldst},
     {ldq_6_bits_uop_ldst},
     {ldq_5_bits_uop_ldst},
     {ldq_4_bits_uop_ldst},
     {ldq_3_bits_uop_ldst},
     {ldq_2_bits_uop_ldst},
     {ldq_1_bits_uop_ldst},
     {ldq_0_bits_uop_ldst}};	// lsu.scala:210:16, :465:79
  wire [15:0][5:0]  _GEN_173 =
    {{ldq_15_bits_uop_lrs1},
     {ldq_14_bits_uop_lrs1},
     {ldq_13_bits_uop_lrs1},
     {ldq_12_bits_uop_lrs1},
     {ldq_11_bits_uop_lrs1},
     {ldq_10_bits_uop_lrs1},
     {ldq_9_bits_uop_lrs1},
     {ldq_8_bits_uop_lrs1},
     {ldq_7_bits_uop_lrs1},
     {ldq_6_bits_uop_lrs1},
     {ldq_5_bits_uop_lrs1},
     {ldq_4_bits_uop_lrs1},
     {ldq_3_bits_uop_lrs1},
     {ldq_2_bits_uop_lrs1},
     {ldq_1_bits_uop_lrs1},
     {ldq_0_bits_uop_lrs1}};	// lsu.scala:210:16, :465:79
  wire [15:0][5:0]  _GEN_174 =
    {{ldq_15_bits_uop_lrs2},
     {ldq_14_bits_uop_lrs2},
     {ldq_13_bits_uop_lrs2},
     {ldq_12_bits_uop_lrs2},
     {ldq_11_bits_uop_lrs2},
     {ldq_10_bits_uop_lrs2},
     {ldq_9_bits_uop_lrs2},
     {ldq_8_bits_uop_lrs2},
     {ldq_7_bits_uop_lrs2},
     {ldq_6_bits_uop_lrs2},
     {ldq_5_bits_uop_lrs2},
     {ldq_4_bits_uop_lrs2},
     {ldq_3_bits_uop_lrs2},
     {ldq_2_bits_uop_lrs2},
     {ldq_1_bits_uop_lrs2},
     {ldq_0_bits_uop_lrs2}};	// lsu.scala:210:16, :465:79
  wire [15:0][5:0]  _GEN_175 =
    {{ldq_15_bits_uop_lrs3},
     {ldq_14_bits_uop_lrs3},
     {ldq_13_bits_uop_lrs3},
     {ldq_12_bits_uop_lrs3},
     {ldq_11_bits_uop_lrs3},
     {ldq_10_bits_uop_lrs3},
     {ldq_9_bits_uop_lrs3},
     {ldq_8_bits_uop_lrs3},
     {ldq_7_bits_uop_lrs3},
     {ldq_6_bits_uop_lrs3},
     {ldq_5_bits_uop_lrs3},
     {ldq_4_bits_uop_lrs3},
     {ldq_3_bits_uop_lrs3},
     {ldq_2_bits_uop_lrs3},
     {ldq_1_bits_uop_lrs3},
     {ldq_0_bits_uop_lrs3}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_176 =
    {{ldq_15_bits_uop_ldst_val},
     {ldq_14_bits_uop_ldst_val},
     {ldq_13_bits_uop_ldst_val},
     {ldq_12_bits_uop_ldst_val},
     {ldq_11_bits_uop_ldst_val},
     {ldq_10_bits_uop_ldst_val},
     {ldq_9_bits_uop_ldst_val},
     {ldq_8_bits_uop_ldst_val},
     {ldq_7_bits_uop_ldst_val},
     {ldq_6_bits_uop_ldst_val},
     {ldq_5_bits_uop_ldst_val},
     {ldq_4_bits_uop_ldst_val},
     {ldq_3_bits_uop_ldst_val},
     {ldq_2_bits_uop_ldst_val},
     {ldq_1_bits_uop_ldst_val},
     {ldq_0_bits_uop_ldst_val}};	// lsu.scala:210:16, :465:79
  wire [15:0][1:0]  _GEN_177 =
    {{ldq_15_bits_uop_dst_rtype},
     {ldq_14_bits_uop_dst_rtype},
     {ldq_13_bits_uop_dst_rtype},
     {ldq_12_bits_uop_dst_rtype},
     {ldq_11_bits_uop_dst_rtype},
     {ldq_10_bits_uop_dst_rtype},
     {ldq_9_bits_uop_dst_rtype},
     {ldq_8_bits_uop_dst_rtype},
     {ldq_7_bits_uop_dst_rtype},
     {ldq_6_bits_uop_dst_rtype},
     {ldq_5_bits_uop_dst_rtype},
     {ldq_4_bits_uop_dst_rtype},
     {ldq_3_bits_uop_dst_rtype},
     {ldq_2_bits_uop_dst_rtype},
     {ldq_1_bits_uop_dst_rtype},
     {ldq_0_bits_uop_dst_rtype}};	// lsu.scala:210:16, :465:79
  wire [15:0][1:0]  _GEN_178 =
    {{ldq_15_bits_uop_lrs1_rtype},
     {ldq_14_bits_uop_lrs1_rtype},
     {ldq_13_bits_uop_lrs1_rtype},
     {ldq_12_bits_uop_lrs1_rtype},
     {ldq_11_bits_uop_lrs1_rtype},
     {ldq_10_bits_uop_lrs1_rtype},
     {ldq_9_bits_uop_lrs1_rtype},
     {ldq_8_bits_uop_lrs1_rtype},
     {ldq_7_bits_uop_lrs1_rtype},
     {ldq_6_bits_uop_lrs1_rtype},
     {ldq_5_bits_uop_lrs1_rtype},
     {ldq_4_bits_uop_lrs1_rtype},
     {ldq_3_bits_uop_lrs1_rtype},
     {ldq_2_bits_uop_lrs1_rtype},
     {ldq_1_bits_uop_lrs1_rtype},
     {ldq_0_bits_uop_lrs1_rtype}};	// lsu.scala:210:16, :465:79
  wire [15:0][1:0]  _GEN_179 =
    {{ldq_15_bits_uop_lrs2_rtype},
     {ldq_14_bits_uop_lrs2_rtype},
     {ldq_13_bits_uop_lrs2_rtype},
     {ldq_12_bits_uop_lrs2_rtype},
     {ldq_11_bits_uop_lrs2_rtype},
     {ldq_10_bits_uop_lrs2_rtype},
     {ldq_9_bits_uop_lrs2_rtype},
     {ldq_8_bits_uop_lrs2_rtype},
     {ldq_7_bits_uop_lrs2_rtype},
     {ldq_6_bits_uop_lrs2_rtype},
     {ldq_5_bits_uop_lrs2_rtype},
     {ldq_4_bits_uop_lrs2_rtype},
     {ldq_3_bits_uop_lrs2_rtype},
     {ldq_2_bits_uop_lrs2_rtype},
     {ldq_1_bits_uop_lrs2_rtype},
     {ldq_0_bits_uop_lrs2_rtype}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_180 =
    {{ldq_15_bits_uop_frs3_en},
     {ldq_14_bits_uop_frs3_en},
     {ldq_13_bits_uop_frs3_en},
     {ldq_12_bits_uop_frs3_en},
     {ldq_11_bits_uop_frs3_en},
     {ldq_10_bits_uop_frs3_en},
     {ldq_9_bits_uop_frs3_en},
     {ldq_8_bits_uop_frs3_en},
     {ldq_7_bits_uop_frs3_en},
     {ldq_6_bits_uop_frs3_en},
     {ldq_5_bits_uop_frs3_en},
     {ldq_4_bits_uop_frs3_en},
     {ldq_3_bits_uop_frs3_en},
     {ldq_2_bits_uop_frs3_en},
     {ldq_1_bits_uop_frs3_en},
     {ldq_0_bits_uop_frs3_en}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_181 =
    {{ldq_15_bits_uop_fp_val},
     {ldq_14_bits_uop_fp_val},
     {ldq_13_bits_uop_fp_val},
     {ldq_12_bits_uop_fp_val},
     {ldq_11_bits_uop_fp_val},
     {ldq_10_bits_uop_fp_val},
     {ldq_9_bits_uop_fp_val},
     {ldq_8_bits_uop_fp_val},
     {ldq_7_bits_uop_fp_val},
     {ldq_6_bits_uop_fp_val},
     {ldq_5_bits_uop_fp_val},
     {ldq_4_bits_uop_fp_val},
     {ldq_3_bits_uop_fp_val},
     {ldq_2_bits_uop_fp_val},
     {ldq_1_bits_uop_fp_val},
     {ldq_0_bits_uop_fp_val}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_182 =
    {{ldq_15_bits_uop_fp_single},
     {ldq_14_bits_uop_fp_single},
     {ldq_13_bits_uop_fp_single},
     {ldq_12_bits_uop_fp_single},
     {ldq_11_bits_uop_fp_single},
     {ldq_10_bits_uop_fp_single},
     {ldq_9_bits_uop_fp_single},
     {ldq_8_bits_uop_fp_single},
     {ldq_7_bits_uop_fp_single},
     {ldq_6_bits_uop_fp_single},
     {ldq_5_bits_uop_fp_single},
     {ldq_4_bits_uop_fp_single},
     {ldq_3_bits_uop_fp_single},
     {ldq_2_bits_uop_fp_single},
     {ldq_1_bits_uop_fp_single},
     {ldq_0_bits_uop_fp_single}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_183 =
    {{ldq_15_bits_uop_xcpt_pf_if},
     {ldq_14_bits_uop_xcpt_pf_if},
     {ldq_13_bits_uop_xcpt_pf_if},
     {ldq_12_bits_uop_xcpt_pf_if},
     {ldq_11_bits_uop_xcpt_pf_if},
     {ldq_10_bits_uop_xcpt_pf_if},
     {ldq_9_bits_uop_xcpt_pf_if},
     {ldq_8_bits_uop_xcpt_pf_if},
     {ldq_7_bits_uop_xcpt_pf_if},
     {ldq_6_bits_uop_xcpt_pf_if},
     {ldq_5_bits_uop_xcpt_pf_if},
     {ldq_4_bits_uop_xcpt_pf_if},
     {ldq_3_bits_uop_xcpt_pf_if},
     {ldq_2_bits_uop_xcpt_pf_if},
     {ldq_1_bits_uop_xcpt_pf_if},
     {ldq_0_bits_uop_xcpt_pf_if}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_184 =
    {{ldq_15_bits_uop_xcpt_ae_if},
     {ldq_14_bits_uop_xcpt_ae_if},
     {ldq_13_bits_uop_xcpt_ae_if},
     {ldq_12_bits_uop_xcpt_ae_if},
     {ldq_11_bits_uop_xcpt_ae_if},
     {ldq_10_bits_uop_xcpt_ae_if},
     {ldq_9_bits_uop_xcpt_ae_if},
     {ldq_8_bits_uop_xcpt_ae_if},
     {ldq_7_bits_uop_xcpt_ae_if},
     {ldq_6_bits_uop_xcpt_ae_if},
     {ldq_5_bits_uop_xcpt_ae_if},
     {ldq_4_bits_uop_xcpt_ae_if},
     {ldq_3_bits_uop_xcpt_ae_if},
     {ldq_2_bits_uop_xcpt_ae_if},
     {ldq_1_bits_uop_xcpt_ae_if},
     {ldq_0_bits_uop_xcpt_ae_if}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_185 =
    {{ldq_15_bits_uop_xcpt_ma_if},
     {ldq_14_bits_uop_xcpt_ma_if},
     {ldq_13_bits_uop_xcpt_ma_if},
     {ldq_12_bits_uop_xcpt_ma_if},
     {ldq_11_bits_uop_xcpt_ma_if},
     {ldq_10_bits_uop_xcpt_ma_if},
     {ldq_9_bits_uop_xcpt_ma_if},
     {ldq_8_bits_uop_xcpt_ma_if},
     {ldq_7_bits_uop_xcpt_ma_if},
     {ldq_6_bits_uop_xcpt_ma_if},
     {ldq_5_bits_uop_xcpt_ma_if},
     {ldq_4_bits_uop_xcpt_ma_if},
     {ldq_3_bits_uop_xcpt_ma_if},
     {ldq_2_bits_uop_xcpt_ma_if},
     {ldq_1_bits_uop_xcpt_ma_if},
     {ldq_0_bits_uop_xcpt_ma_if}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_186 =
    {{ldq_15_bits_uop_bp_debug_if},
     {ldq_14_bits_uop_bp_debug_if},
     {ldq_13_bits_uop_bp_debug_if},
     {ldq_12_bits_uop_bp_debug_if},
     {ldq_11_bits_uop_bp_debug_if},
     {ldq_10_bits_uop_bp_debug_if},
     {ldq_9_bits_uop_bp_debug_if},
     {ldq_8_bits_uop_bp_debug_if},
     {ldq_7_bits_uop_bp_debug_if},
     {ldq_6_bits_uop_bp_debug_if},
     {ldq_5_bits_uop_bp_debug_if},
     {ldq_4_bits_uop_bp_debug_if},
     {ldq_3_bits_uop_bp_debug_if},
     {ldq_2_bits_uop_bp_debug_if},
     {ldq_1_bits_uop_bp_debug_if},
     {ldq_0_bits_uop_bp_debug_if}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_187 =
    {{ldq_15_bits_uop_bp_xcpt_if},
     {ldq_14_bits_uop_bp_xcpt_if},
     {ldq_13_bits_uop_bp_xcpt_if},
     {ldq_12_bits_uop_bp_xcpt_if},
     {ldq_11_bits_uop_bp_xcpt_if},
     {ldq_10_bits_uop_bp_xcpt_if},
     {ldq_9_bits_uop_bp_xcpt_if},
     {ldq_8_bits_uop_bp_xcpt_if},
     {ldq_7_bits_uop_bp_xcpt_if},
     {ldq_6_bits_uop_bp_xcpt_if},
     {ldq_5_bits_uop_bp_xcpt_if},
     {ldq_4_bits_uop_bp_xcpt_if},
     {ldq_3_bits_uop_bp_xcpt_if},
     {ldq_2_bits_uop_bp_xcpt_if},
     {ldq_1_bits_uop_bp_xcpt_if},
     {ldq_0_bits_uop_bp_xcpt_if}};	// lsu.scala:210:16, :465:79
  wire [15:0][1:0]  _GEN_188 =
    {{ldq_15_bits_uop_debug_fsrc},
     {ldq_14_bits_uop_debug_fsrc},
     {ldq_13_bits_uop_debug_fsrc},
     {ldq_12_bits_uop_debug_fsrc},
     {ldq_11_bits_uop_debug_fsrc},
     {ldq_10_bits_uop_debug_fsrc},
     {ldq_9_bits_uop_debug_fsrc},
     {ldq_8_bits_uop_debug_fsrc},
     {ldq_7_bits_uop_debug_fsrc},
     {ldq_6_bits_uop_debug_fsrc},
     {ldq_5_bits_uop_debug_fsrc},
     {ldq_4_bits_uop_debug_fsrc},
     {ldq_3_bits_uop_debug_fsrc},
     {ldq_2_bits_uop_debug_fsrc},
     {ldq_1_bits_uop_debug_fsrc},
     {ldq_0_bits_uop_debug_fsrc}};	// lsu.scala:210:16, :465:79
  wire [15:0][1:0]  _GEN_189 =
    {{ldq_15_bits_uop_debug_tsrc},
     {ldq_14_bits_uop_debug_tsrc},
     {ldq_13_bits_uop_debug_tsrc},
     {ldq_12_bits_uop_debug_tsrc},
     {ldq_11_bits_uop_debug_tsrc},
     {ldq_10_bits_uop_debug_tsrc},
     {ldq_9_bits_uop_debug_tsrc},
     {ldq_8_bits_uop_debug_tsrc},
     {ldq_7_bits_uop_debug_tsrc},
     {ldq_6_bits_uop_debug_tsrc},
     {ldq_5_bits_uop_debug_tsrc},
     {ldq_4_bits_uop_debug_tsrc},
     {ldq_3_bits_uop_debug_tsrc},
     {ldq_2_bits_uop_debug_tsrc},
     {ldq_1_bits_uop_debug_tsrc},
     {ldq_0_bits_uop_debug_tsrc}};	// lsu.scala:210:16, :465:79
  wire [15:0][39:0] _GEN_190 =
    {{ldq_15_bits_addr_bits},
     {ldq_14_bits_addr_bits},
     {ldq_13_bits_addr_bits},
     {ldq_12_bits_addr_bits},
     {ldq_11_bits_addr_bits},
     {ldq_10_bits_addr_bits},
     {ldq_9_bits_addr_bits},
     {ldq_8_bits_addr_bits},
     {ldq_7_bits_addr_bits},
     {ldq_6_bits_addr_bits},
     {ldq_5_bits_addr_bits},
     {ldq_4_bits_addr_bits},
     {ldq_3_bits_addr_bits},
     {ldq_2_bits_addr_bits},
     {ldq_1_bits_addr_bits},
     {ldq_0_bits_addr_bits}};	// lsu.scala:210:16, :465:79
  wire [39:0]       _GEN_191 = _GEN_190[ldq_retry_idx];	// lsu.scala:415:30, :465:79
  wire [15:0]       _GEN_192 =
    {{ldq_15_bits_addr_is_virtual},
     {ldq_14_bits_addr_is_virtual},
     {ldq_13_bits_addr_is_virtual},
     {ldq_12_bits_addr_is_virtual},
     {ldq_11_bits_addr_is_virtual},
     {ldq_10_bits_addr_is_virtual},
     {ldq_9_bits_addr_is_virtual},
     {ldq_8_bits_addr_is_virtual},
     {ldq_7_bits_addr_is_virtual},
     {ldq_6_bits_addr_is_virtual},
     {ldq_5_bits_addr_is_virtual},
     {ldq_4_bits_addr_is_virtual},
     {ldq_3_bits_addr_is_virtual},
     {ldq_2_bits_addr_is_virtual},
     {ldq_1_bits_addr_is_virtual},
     {ldq_0_bits_addr_is_virtual}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_193 =
    {{ldq_15_bits_order_fail},
     {ldq_14_bits_order_fail},
     {ldq_13_bits_order_fail},
     {ldq_12_bits_order_fail},
     {ldq_11_bits_order_fail},
     {ldq_10_bits_order_fail},
     {ldq_9_bits_order_fail},
     {ldq_8_bits_order_fail},
     {ldq_7_bits_order_fail},
     {ldq_6_bits_order_fail},
     {ldq_5_bits_order_fail},
     {ldq_4_bits_order_fail},
     {ldq_3_bits_order_fail},
     {ldq_2_bits_order_fail},
     {ldq_1_bits_order_fail},
     {ldq_0_bits_order_fail}};	// lsu.scala:210:16, :465:79
  wire [15:0]       _GEN_194 =
    {{p1_block_load_mask_15},
     {p1_block_load_mask_14},
     {p1_block_load_mask_13},
     {p1_block_load_mask_12},
     {p1_block_load_mask_11},
     {p1_block_load_mask_10},
     {p1_block_load_mask_9},
     {p1_block_load_mask_8},
     {p1_block_load_mask_7},
     {p1_block_load_mask_6},
     {p1_block_load_mask_5},
     {p1_block_load_mask_4},
     {p1_block_load_mask_3},
     {p1_block_load_mask_2},
     {p1_block_load_mask_1},
     {p1_block_load_mask_0}};	// lsu.scala:398:35, :468:33
  wire [15:0]       _GEN_195 =
    {{p2_block_load_mask_15},
     {p2_block_load_mask_14},
     {p2_block_load_mask_13},
     {p2_block_load_mask_12},
     {p2_block_load_mask_11},
     {p2_block_load_mask_10},
     {p2_block_load_mask_9},
     {p2_block_load_mask_8},
     {p2_block_load_mask_7},
     {p2_block_load_mask_6},
     {p2_block_load_mask_5},
     {p2_block_load_mask_4},
     {p2_block_load_mask_3},
     {p2_block_load_mask_2},
     {p2_block_load_mask_1},
     {p2_block_load_mask_0}};	// lsu.scala:399:35, :469:33
  reg               can_fire_load_retry_REG;	// lsu.scala:470:40
  wire              _GEN_196 = _GEN_2[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [11:0]       _GEN_197 = _GEN_28[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [5:0]        mem_stq_retry_e_out_bits_uop_rob_idx = _GEN_36[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [3:0]        _GEN_198 = _GEN_37[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [3:0]        mem_stq_retry_e_out_bits_uop_stq_idx = _GEN_38[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [6:0]        _GEN_199 = _GEN_40[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [1:0]        mem_stq_retry_e_out_bits_uop_mem_size = _GEN_55[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire              mem_stq_retry_e_out_bits_uop_is_amo = _GEN_61[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  wire [39:0]       _GEN_200 = _GEN_88[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79
  reg               can_fire_sta_retry_REG;	// lsu.scala:482:41
  wire              can_fire_store_commit_0 =
    _GEN_3 & ~_GEN_59 & ~mem_xcpt_valids_0 & ~_GEN_51
    & (_GEN_94[stq_execute_head] | _GEN_62 & _GEN_87[stq_execute_head]
       & ~_GEN_90[stq_execute_head] & _GEN_91[stq_execute_head]);	// lsu.scala:220:29, :224:42, :490:33, :491:33, :492:33, :493:79, :494:62, :496:{66,101}, :667:32
  wire [11:0]       _GEN_201 = _GEN_102[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [3:0]        mem_ldq_wakeup_e_out_bits_uop_stq_idx = _GEN_103[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [1:0]        mem_ldq_wakeup_e_out_bits_uop_mem_size = _GEN_104[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [39:0]       _GEN_202 = _GEN_190[ldq_wakeup_idx];	// lsu.scala:430:31, :465:79, :502:88
  wire              _GEN_203 = _GEN_192[ldq_wakeup_idx];	// lsu.scala:430:31, :465:79, :502:88
  wire [15:0]       _GEN_204 =
    {{ldq_15_bits_addr_is_uncacheable},
     {ldq_14_bits_addr_is_uncacheable},
     {ldq_13_bits_addr_is_uncacheable},
     {ldq_12_bits_addr_is_uncacheable},
     {ldq_11_bits_addr_is_uncacheable},
     {ldq_10_bits_addr_is_uncacheable},
     {ldq_9_bits_addr_is_uncacheable},
     {ldq_8_bits_addr_is_uncacheable},
     {ldq_7_bits_addr_is_uncacheable},
     {ldq_6_bits_addr_is_uncacheable},
     {ldq_5_bits_addr_is_uncacheable},
     {ldq_4_bits_addr_is_uncacheable},
     {ldq_3_bits_addr_is_uncacheable},
     {ldq_2_bits_addr_is_uncacheable},
     {ldq_1_bits_addr_is_uncacheable},
     {ldq_0_bits_addr_is_uncacheable}};	// lsu.scala:210:16, :502:88
  wire              _GEN_205 = _GEN_106[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire [15:0]       _GEN_206 =
    {{ldq_15_bits_succeeded},
     {ldq_14_bits_succeeded},
     {ldq_13_bits_succeeded},
     {ldq_12_bits_succeeded},
     {ldq_11_bits_succeeded},
     {ldq_10_bits_succeeded},
     {ldq_9_bits_succeeded},
     {ldq_8_bits_succeeded},
     {ldq_7_bits_succeeded},
     {ldq_6_bits_succeeded},
     {ldq_5_bits_succeeded},
     {ldq_4_bits_succeeded},
     {ldq_3_bits_succeeded},
     {ldq_2_bits_succeeded},
     {ldq_1_bits_succeeded},
     {ldq_0_bits_succeeded}};	// lsu.scala:210:16, :502:88
  wire [15:0]       mem_ldq_wakeup_e_out_bits_st_dep_mask = _GEN_107[ldq_wakeup_idx];	// lsu.scala:264:49, :430:31, :502:88
  wire              will_fire_stad_incoming_0 =
    _can_fire_sta_incoming_T & io_core_exe_0_req_bits_uop_ctrl_is_std
    & ~can_fire_load_incoming_0 & ~can_fire_load_incoming_0;	// lsu.scala:441:63, :444:63, :534:{35,63}, :535:35
  wire              _will_fire_sta_incoming_0_will_fire_T_2 =
    ~can_fire_load_incoming_0 & ~will_fire_stad_incoming_0;	// lsu.scala:441:63, :534:63, :538:{31,34}
  wire              _will_fire_sta_incoming_0_will_fire_T_6 =
    ~can_fire_load_incoming_0 & ~will_fire_stad_incoming_0;	// lsu.scala:441:63, :534:63, :539:{31,34}
  wire              will_fire_sta_incoming_0 =
    _can_fire_sta_incoming_T & ~io_core_exe_0_req_bits_uop_ctrl_is_std
    & _will_fire_sta_incoming_0_will_fire_T_2 & _will_fire_sta_incoming_0_will_fire_T_6
    & ~will_fire_stad_incoming_0;	// lsu.scala:444:63, :449:66, :534:63, :536:61, :537:35, :538:31, :539:31
  wire              _will_fire_sfence_0_will_fire_T_2 =
    _will_fire_sta_incoming_0_will_fire_T_2 & ~will_fire_sta_incoming_0;	// lsu.scala:536:61, :538:{31,34}
  wire              _will_fire_release_0_will_fire_T_6 =
    _will_fire_sta_incoming_0_will_fire_T_6 & ~will_fire_sta_incoming_0;	// lsu.scala:536:61, :539:{31,34}
  wire              _will_fire_std_incoming_0_will_fire_T_14 =
    ~will_fire_stad_incoming_0 & ~will_fire_sta_incoming_0;	// lsu.scala:534:63, :536:61, :541:{31,34}
  wire              will_fire_std_incoming_0 =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_ctrl_is_std
    & ~io_core_exe_0_req_bits_uop_ctrl_is_sta & _will_fire_std_incoming_0_will_fire_T_14;	// lsu.scala:453:66, :536:61, :541:31
  wire              _will_fire_sfence_0_will_fire_T_14 =
    _will_fire_std_incoming_0_will_fire_T_14 & ~will_fire_std_incoming_0;	// lsu.scala:536:61, :541:{31,34}
  wire              will_fire_sfence_0 =
    io_core_exe_0_req_valid & io_core_exe_0_req_bits_sfence_valid
    & _will_fire_sfence_0_will_fire_T_2 & _will_fire_sfence_0_will_fire_T_14;	// lsu.scala:536:61, :538:31, :541:31
  wire              _will_fire_hella_incoming_0_will_fire_T_2 =
    _will_fire_sfence_0_will_fire_T_2 & ~will_fire_sfence_0;	// lsu.scala:536:61, :538:{31,34}
  wire              will_fire_release_0 =
    io_dmem_release_valid & _will_fire_release_0_will_fire_T_6;	// lsu.scala:534:63, :539:31
  wire              _will_fire_load_retry_0_will_fire_T_6 =
    _will_fire_release_0_will_fire_T_6 & ~will_fire_release_0;	// lsu.scala:534:63, :539:{31,34}
  wire              will_fire_hella_incoming_0 =
    (|hella_state) & _GEN_1 & _will_fire_hella_incoming_0_will_fire_T_2
    & ~can_fire_load_incoming_0;	// lsu.scala:242:38, :441:63, :535:65, :536:35, :538:31, :593:24, :803:26
  wire              _will_fire_load_retry_0_will_fire_T_2 =
    _will_fire_hella_incoming_0_will_fire_T_2 & ~will_fire_hella_incoming_0;	// lsu.scala:535:65, :538:{31,34}
  wire              _will_fire_hella_wakeup_0_will_fire_T_10 =
    ~can_fire_load_incoming_0 & ~will_fire_hella_incoming_0;	// lsu.scala:441:63, :535:65, :540:{31,34}
  wire              will_fire_hella_wakeup_0 =
    _GEN & _GEN_0 & _will_fire_hella_wakeup_0_will_fire_T_10;	// lsu.scala:535:65, :540:31, :820:26, :1527:34, :1533:38, :1550:43, :1553:38, :1560:40, :1576:42
  wire              _will_fire_load_retry_0_will_fire_T_10 =
    _will_fire_hella_wakeup_0_will_fire_T_10 & ~will_fire_hella_wakeup_0;	// lsu.scala:535:65, :540:{31,34}
  wire              will_fire_load_retry_0 =
    _GEN_97[ldq_retry_idx] & _GEN_105[ldq_retry_idx] & _GEN_192[ldq_retry_idx]
    & ~_GEN_194[ldq_retry_idx] & ~_GEN_195[ldq_retry_idx] & can_fire_load_retry_REG
    & ~store_needs_order & ~_GEN_193[ldq_retry_idx]
    & _will_fire_load_retry_0_will_fire_T_2 & _will_fire_load_retry_0_will_fire_T_6
    & _will_fire_load_retry_0_will_fire_T_10;	// lsu.scala:264:49, :305:44, :415:30, :465:79, :468:33, :469:33, :470:40, :471:33, :473:33, :535:65, :538:31, :539:31, :540:31, :1495:3, :1496:64
  wire              _will_fire_sta_retry_0_will_fire_T_2 =
    _will_fire_load_retry_0_will_fire_T_2 & ~will_fire_load_retry_0;	// lsu.scala:535:65, :538:{31,34}
  wire              _will_fire_sta_retry_0_will_fire_T_6 =
    _will_fire_load_retry_0_will_fire_T_6 & ~will_fire_load_retry_0;	// lsu.scala:535:65, :539:{31,34}
  wire              _will_fire_load_wakeup_0_will_fire_T_10 =
    _will_fire_load_retry_0_will_fire_T_10 & ~will_fire_load_retry_0;	// lsu.scala:535:65, :540:{31,34}
  wire              will_fire_sta_retry_0 =
    _GEN_196 & _GEN_87[stq_retry_idx] & _GEN_90[stq_retry_idx] & can_fire_sta_retry_REG
    & _will_fire_sta_retry_0_will_fire_T_2 & _will_fire_sta_retry_0_will_fire_T_6
    & _will_fire_sfence_0_will_fire_T_14 & ~will_fire_sfence_0;	// lsu.scala:224:42, :422:30, :478:79, :482:41, :536:61, :538:31, :539:31, :541:{31,34}
  assign _will_fire_store_commit_0_T_2 =
    _will_fire_sta_retry_0_will_fire_T_2 & ~will_fire_sta_retry_0;	// lsu.scala:536:61, :538:{31,34}
  wire              will_fire_load_wakeup_0 =
    _GEN_97[ldq_wakeup_idx] & _GEN_105[ldq_wakeup_idx] & ~_GEN_206[ldq_wakeup_idx]
    & ~_GEN_203 & ~_GEN_205 & ~_GEN_193[ldq_wakeup_idx] & ~_GEN_194[ldq_wakeup_idx]
    & ~_GEN_195[ldq_wakeup_idx] & ~store_needs_order & ~block_load_wakeup
    & (~_GEN_204[ldq_wakeup_idx] | io_core_commit_load_at_rob_head
       & ldq_head == ldq_wakeup_idx & mem_ldq_wakeup_e_out_bits_st_dep_mask == 16'h0)
    & _will_fire_sta_retry_0_will_fire_T_6 & ~will_fire_sta_retry_0
    & _will_fire_load_wakeup_0_will_fire_T_10;	// lsu.scala:215:29, :259:32, :264:49, :305:44, :430:31, :465:79, :468:33, :469:33, :471:33, :502:88, :504:31, :505:31, :506:31, :507:31, :508:31, :509:31, :511:31, :513:{32,71}, :514:{84,103}, :515:112, :535:65, :536:61, :539:{31,34}, :540:31, :1199:80, :1210:43, :1211:25, :1495:3, :1496:64
  wire              will_fire_store_commit_0 =
    can_fire_store_commit_0 & _will_fire_load_wakeup_0_will_fire_T_10
    & ~will_fire_load_wakeup_0;	// lsu.scala:493:79, :535:65, :540:{31,34}
  wire              _exe_cmd_T = can_fire_load_incoming_0 | will_fire_stad_incoming_0;	// lsu.scala:441:63, :534:63, :567:63
  wire              _GEN_207 = _exe_cmd_T | will_fire_sta_incoming_0;	// lsu.scala:536:61, :567:{63,93}
  wire              _GEN_208 = ldq_wakeup_idx == 4'h0;	// lsu.scala:430:31, :570:49
  wire              _GEN_209 = ldq_wakeup_idx == 4'h1;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_210 = ldq_wakeup_idx == 4'h2;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_211 = ldq_wakeup_idx == 4'h3;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_212 = ldq_wakeup_idx == 4'h4;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_213 = ldq_wakeup_idx == 4'h5;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_214 = ldq_wakeup_idx == 4'h6;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_215 = ldq_wakeup_idx == 4'h7;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_216 = ldq_wakeup_idx == 4'h8;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_217 = ldq_wakeup_idx == 4'h9;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_218 = ldq_wakeup_idx == 4'hA;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_219 = ldq_wakeup_idx == 4'hB;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_220 = ldq_wakeup_idx == 4'hC;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_221 = ldq_wakeup_idx == 4'hD;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_222 = ldq_wakeup_idx == 4'hE;	// lsu.scala:305:44, :430:31, :570:49
  wire              _GEN_223 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h0;	// lsu.scala:572:52
  wire              _GEN_224 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h1;	// lsu.scala:305:44, :572:52
  wire              _GEN_225 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h2;	// lsu.scala:305:44, :572:52
  wire              _GEN_226 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h3;	// lsu.scala:305:44, :572:52
  wire              _GEN_227 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h4;	// lsu.scala:305:44, :572:52
  wire              _GEN_228 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h5;	// lsu.scala:305:44, :572:52
  wire              _GEN_229 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h6;	// lsu.scala:305:44, :572:52
  wire              _GEN_230 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h7;	// lsu.scala:305:44, :572:52
  wire              _GEN_231 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h8;	// lsu.scala:305:44, :572:52
  wire              _GEN_232 = io_core_exe_0_req_bits_uop_ldq_idx == 4'h9;	// lsu.scala:305:44, :572:52
  wire              _GEN_233 = io_core_exe_0_req_bits_uop_ldq_idx == 4'hA;	// lsu.scala:305:44, :572:52
  wire              _GEN_234 = io_core_exe_0_req_bits_uop_ldq_idx == 4'hB;	// lsu.scala:305:44, :572:52
  wire              _GEN_235 = io_core_exe_0_req_bits_uop_ldq_idx == 4'hC;	// lsu.scala:305:44, :572:52
  wire              _GEN_236 = io_core_exe_0_req_bits_uop_ldq_idx == 4'hD;	// lsu.scala:305:44, :572:52
  wire              _GEN_237 = io_core_exe_0_req_bits_uop_ldq_idx == 4'hE;	// lsu.scala:305:44, :572:52
  wire              _GEN_238 = ldq_retry_idx == 4'h0;	// lsu.scala:415:30, :574:49
  wire              _GEN_239 = will_fire_load_retry_0 & _GEN_238;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_240 = ldq_retry_idx == 4'h1;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_241 = will_fire_load_retry_0 & _GEN_240;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_242 = ldq_retry_idx == 4'h2;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_243 = will_fire_load_retry_0 & _GEN_242;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_244 = ldq_retry_idx == 4'h3;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_245 = will_fire_load_retry_0 & _GEN_244;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_246 = ldq_retry_idx == 4'h4;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_247 = will_fire_load_retry_0 & _GEN_246;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_248 = ldq_retry_idx == 4'h5;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_249 = will_fire_load_retry_0 & _GEN_248;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_250 = ldq_retry_idx == 4'h6;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_251 = will_fire_load_retry_0 & _GEN_250;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_252 = ldq_retry_idx == 4'h7;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_253 = will_fire_load_retry_0 & _GEN_252;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_254 = ldq_retry_idx == 4'h8;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_255 = will_fire_load_retry_0 & _GEN_254;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_256 = ldq_retry_idx == 4'h9;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_257 = will_fire_load_retry_0 & _GEN_256;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_258 = ldq_retry_idx == 4'hA;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_259 = will_fire_load_retry_0 & _GEN_258;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_260 = ldq_retry_idx == 4'hB;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_261 = will_fire_load_retry_0 & _GEN_260;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_262 = ldq_retry_idx == 4'hC;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_263 = will_fire_load_retry_0 & _GEN_262;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_264 = ldq_retry_idx == 4'hD;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_265 = will_fire_load_retry_0 & _GEN_264;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_266 = ldq_retry_idx == 4'hE;	// lsu.scala:305:44, :415:30, :574:49
  wire              _GEN_267 = will_fire_load_retry_0 & _GEN_266;	// lsu.scala:535:65, :573:43, :574:49
  wire              _GEN_268 = will_fire_load_retry_0 & (&ldq_retry_idx);	// lsu.scala:415:30, :535:65, :573:43, :574:49
  wire              _exe_tlb_uop_T_2 =
    _exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0;	// lsu.scala:536:61, :567:63, :599:53
  wire              _exe_tlb_uop_T_4_uses_ldq =
    will_fire_sta_retry_0 & _GEN_63[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79, :536:61, :602:24
  wire              _exe_tlb_uop_T_4_uses_stq =
    will_fire_sta_retry_0 & _GEN_64[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79, :536:61, :602:24
  wire              exe_tlb_uop_0_ctrl_is_load =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_ctrl_is_load
      : will_fire_load_retry_0
          ? _GEN_122[ldq_retry_idx]
          : will_fire_sta_retry_0 & _GEN_18[stq_retry_idx];	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire              exe_tlb_uop_0_ctrl_is_sta =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_ctrl_is_sta
      : will_fire_load_retry_0
          ? _GEN_123[ldq_retry_idx]
          : will_fire_sta_retry_0 & _GEN_19[stq_retry_idx];	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire [11:0]       exe_tlb_uop_0_br_mask =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_br_mask
      : will_fire_load_retry_0 ? _GEN_132 : will_fire_sta_retry_0 ? _GEN_197 : 12'h0;	// lsu.scala:465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire [4:0]        exe_tlb_uop_0_mem_cmd =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_mem_cmd
      : will_fire_load_retry_0
          ? _GEN_159[ldq_retry_idx]
          : will_fire_sta_retry_0 ? _GEN_54[stq_retry_idx] : 5'h0;	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire [1:0]        exe_tlb_uop_0_mem_size =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_mem_size
      : will_fire_load_retry_0
          ? mem_ldq_retry_e_out_bits_uop_mem_size
          : will_fire_sta_retry_0 ? mem_stq_retry_e_out_bits_uop_mem_size : 2'h0;	// lsu.scala:465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire              exe_tlb_uop_0_is_fence =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_is_fence
      : will_fire_load_retry_0
          ? _GEN_161[ldq_retry_idx]
          : will_fire_sta_retry_0 & _GEN_58[stq_retry_idx];	// lsu.scala:224:42, :415:30, :422:30, :465:79, :478:79, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24
  wire              _mem_xcpt_uops_WIRE_0_uses_ldq =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_uses_ldq
      : will_fire_load_retry_0 ? _GEN_165 : _exe_tlb_uop_T_4_uses_ldq;	// lsu.scala:465:79, :535:65, :597:24, :599:53, :601:24, :602:24
  wire              _mem_xcpt_uops_WIRE_0_uses_stq =
    _exe_tlb_uop_T_2
      ? io_core_exe_0_req_bits_uop_uses_stq
      : will_fire_load_retry_0 ? _GEN_167 : _exe_tlb_uop_T_4_uses_stq;	// lsu.scala:465:79, :535:65, :597:24, :599:53, :601:24, :602:24
  wire              _exe_tlb_vaddr_T_1 = _exe_cmd_T | will_fire_sta_incoming_0;	// lsu.scala:536:61, :567:63, :608:53
  wire [39:0]       _GEN_269 = {1'h0, io_core_exe_0_req_bits_sfence_bits_addr};	// lsu.scala:249:20, :610:24, :708:86
  wire [39:0]       exe_tlb_vaddr_0 =
    _exe_tlb_vaddr_T_1
      ? io_core_exe_0_req_bits_addr
      : will_fire_sfence_0
          ? _GEN_269
          : will_fire_load_retry_0
              ? _GEN_191
              : will_fire_sta_retry_0
                  ? _GEN_200
                  : will_fire_hella_incoming_0 ? hella_req_addr : 40'h0;	// lsu.scala:243:34, :465:79, :478:79, :535:65, :536:61, :607:24, :608:53, :610:24, :611:24, :612:24, :613:24
  wire              _stq_idx_T = will_fire_sta_incoming_0 | will_fire_stad_incoming_0;	// lsu.scala:534:63, :536:61, :660:56
  reg  [11:0]       mem_xcpt_uops_0_br_mask;	// lsu.scala:671:32
  reg  [5:0]        mem_xcpt_uops_0_rob_idx;	// lsu.scala:671:32
  reg  [3:0]        mem_xcpt_uops_0_ldq_idx;	// lsu.scala:671:32
  reg  [3:0]        mem_xcpt_uops_0_stq_idx;	// lsu.scala:671:32
  reg               mem_xcpt_uops_0_uses_ldq;	// lsu.scala:671:32
  reg               mem_xcpt_uops_0_uses_stq;	// lsu.scala:671:32
  reg  [3:0]        mem_xcpt_causes_0;	// lsu.scala:672:32
  reg  [39:0]       mem_xcpt_vaddrs_0;	// lsu.scala:679:32
  wire              exe_tlb_miss_0 =
    ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_miss;	// lsu.scala:249:20, :538:31, :576:25, :708:58
  wire [31:0]       exe_tlb_paddr_0 =
    {_dtlb_io_resp_0_paddr[31:12], exe_tlb_vaddr_0[11:0]};	// Cat.scala:30:58, lsu.scala:249:20, :607:24, :709:62, :710:57
  reg               REG;	// lsu.scala:718:21
  wire [39:0]       _GEN_270 =
    {8'h0, _dtlb_io_resp_0_paddr[31:12], exe_tlb_vaddr_0[11:0]};	// lsu.scala:249:20, :607:24, :709:62, :710:57, :768:30
  wire [3:0][63:0]  _GEN_271 =
    {{_GEN_93},
     {{2{_GEN_93[31:0]}}},
     {{2{{2{_GEN_93[15:0]}}}}},
     {{2{{2{{2{_GEN_93[7:0]}}}}}}}};	// AMOALU.scala:26:{13,19,66}, Cat.scala:30:58, lsu.scala:224:42
  wire              _GEN_272 = can_fire_load_incoming_0 | will_fire_load_retry_0;	// lsu.scala:220:29, :441:63, :535:65, :766:39, :773:43, :780:45
  assign _GEN_1 = hella_state == 3'h1;	// lsu.scala:242:38, :803:26
  wire              _GEN_273 = will_fire_store_commit_0 | will_fire_load_wakeup_0;	// lsu.scala:245:34, :535:65, :780:45, :794:44, :802:47
  assign _GEN_0 = hella_state == 3'h5;	// lsu.scala:242:38, :820:26, util.scala:351:72
  wire              dmem_req_0_valid =
    can_fire_load_incoming_0
      ? ~exe_tlb_miss_0 & _dtlb_io_resp_0_cacheable
      : will_fire_load_retry_0
          ? ~exe_tlb_miss_0 & _dtlb_io_resp_0_cacheable
          : _GEN_273
            | (will_fire_hella_incoming_0
                 ? ~io_hellacache_s1_kill & (~exe_tlb_miss_0 | hella_req_phys)
                 : will_fire_hella_wakeup_0);	// lsu.scala:243:34, :245:34, :249:20, :441:63, :535:65, :708:58, :766:39, :767:{30,33,50}, :773:43, :774:{30,33,50}, :780:45, :781:33, :794:44, :795:30, :802:47, :805:{39,42,65,69,86}, :819:5
  wire [39:0]       _GEN_274 = {8'h0, hella_paddr};	// lsu.scala:245:34, :768:30, :822:39
  wire              _GEN_275 = can_fire_load_incoming_0 | will_fire_load_retry_0;	// lsu.scala:441:63, :535:65, :766:39, :768:30, :773:43
  wire [3:0][63:0]  _GEN_276 =
    {{hella_data_data},
     {{2{hella_data_data[31:0]}}},
     {{2{{2{hella_data_data[15:0]}}}}},
     {{2{{2{{2{hella_data_data[7:0]}}}}}}}};	// AMOALU.scala:26:{13,19,66}, Cat.scala:30:58, lsu.scala:244:34
  wire              _GEN_277 = will_fire_hella_incoming_0 | will_fire_hella_wakeup_0;	// lsu.scala:535:65, :759:28, :802:47, :811:39, :819:5, :827:39
  wire              _GEN_278 = _stq_idx_T | will_fire_sta_retry_0;	// lsu.scala:536:61, :660:56, :848:67
  wire              _io_core_fp_stdata_ready_output =
    ~will_fire_std_incoming_0 & ~will_fire_stad_incoming_0;	// lsu.scala:534:63, :536:61, :866:{34,61,64}
  wire              fp_stdata_fire =
    _io_core_fp_stdata_ready_output & io_core_fp_stdata_valid;	// Decoupled.scala:40:37, lsu.scala:866:61
  wire              _stq_bits_data_bits_T =
    will_fire_std_incoming_0 | will_fire_stad_incoming_0;	// lsu.scala:534:63, :536:61, :868:37
  wire              _GEN_279 = _stq_bits_data_bits_T | fp_stdata_fire;	// Decoupled.scala:40:37, lsu.scala:868:{37,67}
  wire [3:0]        sidx =
    _stq_bits_data_bits_T
      ? io_core_exe_0_req_bits_uop_stq_idx
      : io_core_fp_stdata_bits_uop_stq_idx;	// lsu.scala:868:37, :870:21
  reg               fired_load_incoming_REG;	// lsu.scala:894:51
  reg               fired_stad_incoming_REG;	// lsu.scala:895:51
  reg               fired_sta_incoming_REG;	// lsu.scala:896:51
  reg               fired_std_incoming_REG;	// lsu.scala:897:51
  reg               fired_stdf_incoming;	// lsu.scala:898:37
  reg               fired_sfence_0;	// lsu.scala:899:37
  reg               fired_release_0;	// lsu.scala:900:37
  reg               fired_load_retry_REG;	// lsu.scala:901:51
  reg               fired_sta_retry_REG;	// lsu.scala:902:51
  reg               fired_load_wakeup_REG;	// lsu.scala:904:51
  reg  [11:0]       mem_incoming_uop_0_br_mask;	// lsu.scala:908:37
  reg  [5:0]        mem_incoming_uop_0_rob_idx;	// lsu.scala:908:37
  reg  [3:0]        mem_incoming_uop_0_ldq_idx;	// lsu.scala:908:37
  reg  [3:0]        mem_incoming_uop_0_stq_idx;	// lsu.scala:908:37
  reg  [6:0]        mem_incoming_uop_0_pdst;	// lsu.scala:908:37
  reg               mem_incoming_uop_0_fp_val;	// lsu.scala:908:37
  reg  [11:0]       mem_ldq_incoming_e_0_bits_uop_br_mask;	// lsu.scala:909:37
  reg  [3:0]        mem_ldq_incoming_e_0_bits_uop_stq_idx;	// lsu.scala:909:37
  reg  [1:0]        mem_ldq_incoming_e_0_bits_uop_mem_size;	// lsu.scala:909:37
  reg  [15:0]       mem_ldq_incoming_e_0_bits_st_dep_mask;	// lsu.scala:909:37
  reg               mem_stq_incoming_e_0_valid;	// lsu.scala:910:37
  reg  [11:0]       mem_stq_incoming_e_0_bits_uop_br_mask;	// lsu.scala:910:37
  reg  [5:0]        mem_stq_incoming_e_0_bits_uop_rob_idx;	// lsu.scala:910:37
  reg  [3:0]        mem_stq_incoming_e_0_bits_uop_stq_idx;	// lsu.scala:910:37
  reg  [1:0]        mem_stq_incoming_e_0_bits_uop_mem_size;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_uop_is_amo;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_addr_valid;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_addr_is_virtual;	// lsu.scala:910:37
  reg               mem_stq_incoming_e_0_bits_data_valid;	// lsu.scala:910:37
  reg  [11:0]       mem_ldq_wakeup_e_bits_uop_br_mask;	// lsu.scala:911:37
  reg  [3:0]        mem_ldq_wakeup_e_bits_uop_stq_idx;	// lsu.scala:911:37
  reg  [1:0]        mem_ldq_wakeup_e_bits_uop_mem_size;	// lsu.scala:911:37
  reg  [15:0]       mem_ldq_wakeup_e_bits_st_dep_mask;	// lsu.scala:911:37
  reg  [11:0]       mem_ldq_retry_e_bits_uop_br_mask;	// lsu.scala:912:37
  reg  [3:0]        mem_ldq_retry_e_bits_uop_stq_idx;	// lsu.scala:912:37
  reg  [1:0]        mem_ldq_retry_e_bits_uop_mem_size;	// lsu.scala:912:37
  reg  [15:0]       mem_ldq_retry_e_bits_st_dep_mask;	// lsu.scala:912:37
  reg               mem_stq_retry_e_valid;	// lsu.scala:913:37
  reg  [11:0]       mem_stq_retry_e_bits_uop_br_mask;	// lsu.scala:913:37
  reg  [5:0]        mem_stq_retry_e_bits_uop_rob_idx;	// lsu.scala:913:37
  reg  [3:0]        mem_stq_retry_e_bits_uop_stq_idx;	// lsu.scala:913:37
  reg  [1:0]        mem_stq_retry_e_bits_uop_mem_size;	// lsu.scala:913:37
  reg               mem_stq_retry_e_bits_uop_is_amo;	// lsu.scala:913:37
  reg               mem_stq_retry_e_bits_data_valid;	// lsu.scala:913:37
  wire [15:0]       lcam_st_dep_mask_0 =
    fired_load_incoming_REG
      ? mem_ldq_incoming_e_0_bits_st_dep_mask
      : fired_load_retry_REG
          ? mem_ldq_retry_e_bits_st_dep_mask
          : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_st_dep_mask : 16'h0;	// lsu.scala:259:32, :894:51, :901:51, :904:51, :909:37, :911:37, :912:37, :915:33, :916:33, :917:33
  wire              _lcam_stq_idx_T = fired_stad_incoming_REG | fired_sta_incoming_REG;	// lsu.scala:895:51, :896:51, :919:57
  reg  [11:0]       mem_stdf_uop_br_mask;	// lsu.scala:922:37
  reg  [5:0]        mem_stdf_uop_rob_idx;	// lsu.scala:922:37
  reg  [3:0]        mem_stdf_uop_stq_idx;	// lsu.scala:922:37
  reg               mem_tlb_miss_0;	// lsu.scala:925:41
  reg               mem_tlb_uncacheable_0;	// lsu.scala:926:41
  reg  [39:0]       mem_paddr_0;	// lsu.scala:927:41
  reg               clr_bsy_valid_0;	// lsu.scala:930:32
  reg  [5:0]        clr_bsy_rob_idx_0;	// lsu.scala:931:28
  reg  [11:0]       clr_bsy_brmask_0;	// lsu.scala:932:28
  reg               io_core_clr_bsy_0_valid_REG;	// lsu.scala:979:62
  reg               io_core_clr_bsy_0_valid_REG_1;	// lsu.scala:979:101
  reg               io_core_clr_bsy_0_valid_REG_2;	// lsu.scala:979:93
  reg               stdf_clr_bsy_valid;	// lsu.scala:983:37
  reg  [5:0]        stdf_clr_bsy_rob_idx;	// lsu.scala:984:33
  reg  [11:0]       stdf_clr_bsy_brmask;	// lsu.scala:985:33
  reg               io_core_clr_bsy_1_valid_REG;	// lsu.scala:1004:67
  reg               io_core_clr_bsy_1_valid_REG_1;	// lsu.scala:1004:106
  reg               io_core_clr_bsy_1_valid_REG_2;	// lsu.scala:1004:98
  wire              do_st_search_0 =
    (_lcam_stq_idx_T | fired_sta_retry_REG) & ~mem_tlb_miss_0;	// lsu.scala:902:51, :919:57, :925:41, :1014:{85,108,111}
  wire              _can_forward_T = fired_load_incoming_REG | fired_load_retry_REG;	// lsu.scala:894:51, :901:51, :1016:61
  wire              do_ld_search_0 =
    _can_forward_T & ~mem_tlb_miss_0 | fired_load_wakeup_REG;	// lsu.scala:904:51, :925:41, :1014:111, :1016:{61,85,106}
  wire              _lcam_addr_T_1 = _lcam_stq_idx_T | fired_sta_retry_REG;	// lsu.scala:902:51, :919:57, :1025:86
  reg  [31:0]       lcam_addr_REG;	// lsu.scala:1026:45
  reg  [31:0]       lcam_addr_REG_1;	// lsu.scala:1027:67
  wire [39:0]       _GEN_280 = {8'h0, lcam_addr_REG_1};	// lsu.scala:768:30, :1027:{41,67}
  wire [39:0]       _GEN_281 = {8'h0, lcam_addr_REG};	// lsu.scala:768:30, :1025:37, :1026:45
  wire [39:0]       lcam_addr_0 =
    _lcam_addr_T_1 ? _GEN_281 : fired_release_0 ? _GEN_280 : mem_paddr_0;	// lsu.scala:900:37, :927:41, :1025:{37,86}, :1027:41
  wire [14:0]       _lcam_mask_mask_T_2 = 15'h1 << lcam_addr_0[2:0];	// lsu.scala:1025:37, :1663:{48,55}
  wire [14:0]       _lcam_mask_mask_T_6 = 15'h3 << {12'h0, lcam_addr_0[2:1], 1'h0};	// lsu.scala:249:20, :708:86, :1025:37, :1664:{48,56}
  wire [3:0][7:0]   _GEN_282 =
    {{8'hFF},
     {lcam_addr_0[2] ? 8'hF0 : 8'hF},
     {_lcam_mask_mask_T_6[7:0]},
     {_lcam_mask_mask_T_2[7:0]}};	// Mux.scala:98:16, lsu.scala:1025:37, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire [7:0]        lcam_mask_0 =
    _GEN_282[do_st_search_0
               ? (_lcam_stq_idx_T
                    ? mem_stq_incoming_e_0_bits_uop_mem_size
                    : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_mem_size : 2'h0)
               : do_ld_search_0
                   ? (fired_load_incoming_REG
                        ? mem_ldq_incoming_e_0_bits_uop_mem_size
                        : fired_load_retry_REG
                            ? mem_ldq_retry_e_bits_uop_mem_size
                            : fired_load_wakeup_REG
                                ? mem_ldq_wakeup_e_bits_uop_mem_size
                                : 2'h0)
                   : 2'h0];	// Mux.scala:98:16, lsu.scala:894:51, :901:51, :902:51, :904:51, :909:37, :910:37, :911:37, :912:37, :913:37, :915:33, :916:33, :917:33, :919:{33,57}, :921:33, :1014:108, :1016:106, :1029:37, :1030:37, :1663:26, :1664:26, :1665:26
  reg  [3:0]        lcam_ldq_idx_REG;	// lsu.scala:1037:58
  reg  [3:0]        lcam_ldq_idx_REG_1;	// lsu.scala:1038:58
  wire [3:0]        lcam_ldq_idx_0 =
    fired_load_incoming_REG
      ? mem_incoming_uop_0_ldq_idx
      : fired_load_wakeup_REG
          ? lcam_ldq_idx_REG
          : fired_load_retry_REG ? lcam_ldq_idx_REG_1 : 4'h0;	// lsu.scala:894:51, :901:51, :904:51, :908:37, :1036:26, :1037:{26,58}, :1038:{26,58}
  reg  [3:0]        lcam_stq_idx_REG;	// lsu.scala:1042:58
  wire [3:0]        lcam_stq_idx_0 =
    _lcam_stq_idx_T
      ? mem_incoming_uop_0_stq_idx
      : fired_sta_retry_REG ? lcam_stq_idx_REG : 4'h0;	// lsu.scala:902:51, :908:37, :919:57, :1040:26, :1042:{26,58}
  reg               s1_executing_loads_0;	// lsu.scala:1056:35
  reg               s1_executing_loads_1;	// lsu.scala:1056:35
  reg               s1_executing_loads_2;	// lsu.scala:1056:35
  reg               s1_executing_loads_3;	// lsu.scala:1056:35
  reg               s1_executing_loads_4;	// lsu.scala:1056:35
  reg               s1_executing_loads_5;	// lsu.scala:1056:35
  reg               s1_executing_loads_6;	// lsu.scala:1056:35
  reg               s1_executing_loads_7;	// lsu.scala:1056:35
  reg               s1_executing_loads_8;	// lsu.scala:1056:35
  reg               s1_executing_loads_9;	// lsu.scala:1056:35
  reg               s1_executing_loads_10;	// lsu.scala:1056:35
  reg               s1_executing_loads_11;	// lsu.scala:1056:35
  reg               s1_executing_loads_12;	// lsu.scala:1056:35
  reg               s1_executing_loads_13;	// lsu.scala:1056:35
  reg               s1_executing_loads_14;	// lsu.scala:1056:35
  reg               s1_executing_loads_15;	// lsu.scala:1056:35
  reg               wb_forward_valid_0;	// lsu.scala:1064:36
  reg  [3:0]        wb_forward_ldq_idx_0;	// lsu.scala:1065:36
  reg  [39:0]       wb_forward_ld_addr_0;	// lsu.scala:1066:36
  reg  [3:0]        wb_forward_stq_idx_0;	// lsu.scala:1067:36
  wire [14:0]       _l_mask_mask_T_2 = 15'h1 << ldq_0_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_6 = 15'h3 << {12'h0, ldq_0_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_283 =
    {{8'hFF},
     {ldq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_6[7:0]},
     {_l_mask_mask_T_2[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_0 = wb_forward_valid_0 & ~(|wb_forward_ldq_idx_0);	// lsu.scala:1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_0 =
    lcam_addr_0[39:6] == ldq_0_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_0 =
    block_addr_matches_0 & lcam_addr_0[5:3] == ldq_0_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T = _GEN_283[ldq_0_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_284 =
    fired_release_0 & ldq_0_valid & ldq_0_bits_addr_valid & block_addr_matches_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_285 = ldq_0_bits_executed | ldq_0_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_286 = _GEN_285 | l_forwarders_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_287 = {12'h0, lcam_stq_idx_0};	// lsu.scala:1040:26, :1100:38
  wire [15:0]       _GEN_288 = ldq_0_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_289 =
    do_st_search_0 & ldq_0_valid & ldq_0_bits_addr_valid & _GEN_286
    & ~ldq_0_bits_addr_is_virtual & _GEN_288[0] & dword_addr_matches_0
    & (|_mask_overlap_T);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_290 =
    do_ld_search_0 & ldq_0_valid & ldq_0_bits_addr_valid & ~ldq_0_bits_addr_is_virtual
    & dword_addr_matches_0 & (|_mask_overlap_T);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older = lcam_ldq_idx_0 < ldq_head ^ (|ldq_head);	// lsu.scala:215:29, :1036:26, util.scala:363:{64,72,78}
  reg               older_nacked_REG;	// lsu.scala:1128:57
  wire              _GEN_291 = ~_GEN_285 | nacking_loads_0 | older_nacked_REG;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_292 = _GEN_284 | _GEN_289;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG;	// lsu.scala:1131:58
  wire              _GEN_293 = (|lcam_ldq_idx_0) & _GEN_291;	// lsu.scala:764:24, :1036:26, :1125:{38,47}, :1129:{56,73}, :1131:48
  wire [14:0]       _l_mask_mask_T_17 = 15'h1 << ldq_1_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_21 = 15'h3 << {12'h0, ldq_1_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_294 =
    {{8'hFF},
     {ldq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_21[7:0]},
     {_l_mask_mask_T_17[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_1_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h1;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_1_0 =
    lcam_addr_0[39:6] == ldq_1_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_1_0 =
    block_addr_matches_1_0 & lcam_addr_0[5:3] == ldq_1_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_2 = _GEN_294[ldq_1_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_295 =
    fired_release_0 & ldq_1_valid & ldq_1_bits_addr_valid & block_addr_matches_1_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_296 = ldq_1_bits_executed | ldq_1_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_297 = _GEN_296 | l_forwarders_1_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_298 = ldq_1_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_299 =
    do_st_search_0 & ldq_1_valid & ldq_1_bits_addr_valid & _GEN_297
    & ~ldq_1_bits_addr_is_virtual & _GEN_298[0] & dword_addr_matches_1_0
    & (|_mask_overlap_T_2);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_300 =
    do_ld_search_0 & ldq_1_valid & ldq_1_bits_addr_valid & ~ldq_1_bits_addr_is_virtual
    & dword_addr_matches_1_0 & (|_mask_overlap_T_2);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_1 =
    lcam_ldq_idx_0 == 4'h0 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[3:1]));	// lsu.scala:215:29, :1036:26, util.scala:351:72, :363:{52,64,72,78}
  wire              _GEN_301 = lcam_ldq_idx_0 != 4'h1;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_1;	// lsu.scala:1128:57
  wire              _GEN_302 = ~_GEN_296 | nacking_loads_1 | older_nacked_REG_1;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_303 = _GEN_295 | _GEN_299;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_1;	// lsu.scala:1131:58
  wire              _GEN_304 =
    _GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_32 = 15'h1 << ldq_2_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_36 = 15'h3 << {12'h0, ldq_2_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_305 =
    {{8'hFF},
     {ldq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_36[7:0]},
     {_l_mask_mask_T_32[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_2_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h2;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_2_0 =
    lcam_addr_0[39:6] == ldq_2_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_2_0 =
    block_addr_matches_2_0 & lcam_addr_0[5:3] == ldq_2_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_4 = _GEN_305[ldq_2_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_306 =
    fired_release_0 & ldq_2_valid & ldq_2_bits_addr_valid & block_addr_matches_2_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_307 = ldq_2_bits_executed | ldq_2_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_308 = _GEN_307 | l_forwarders_2_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_309 = ldq_2_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_310 =
    do_st_search_0 & ldq_2_valid & ldq_2_bits_addr_valid & _GEN_308
    & ~ldq_2_bits_addr_is_virtual & _GEN_309[0] & dword_addr_matches_2_0
    & (|_mask_overlap_T_4);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_311 =
    do_ld_search_0 & ldq_2_valid & ldq_2_bits_addr_valid & ~ldq_2_bits_addr_is_virtual
    & dword_addr_matches_2_0 & (|_mask_overlap_T_4);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_2 =
    lcam_ldq_idx_0 < 4'h2 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'h2;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_312 = lcam_ldq_idx_0 != 4'h2;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_2;	// lsu.scala:1128:57
  wire              _GEN_313 = ~_GEN_307 | nacking_loads_2 | older_nacked_REG_2;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_314 = _GEN_306 | _GEN_310;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_2;	// lsu.scala:1131:58
  wire              _GEN_315 =
    _GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_47 = 15'h1 << ldq_3_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_51 = 15'h3 << {12'h0, ldq_3_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_316 =
    {{8'hFF},
     {ldq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_51[7:0]},
     {_l_mask_mask_T_47[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_3_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h3;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_3_0 =
    lcam_addr_0[39:6] == ldq_3_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_3_0 =
    block_addr_matches_3_0 & lcam_addr_0[5:3] == ldq_3_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_6 = _GEN_316[ldq_3_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_317 =
    fired_release_0 & ldq_3_valid & ldq_3_bits_addr_valid & block_addr_matches_3_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_318 = ldq_3_bits_executed | ldq_3_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_319 = _GEN_318 | l_forwarders_3_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_320 = ldq_3_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_321 =
    do_st_search_0 & ldq_3_valid & ldq_3_bits_addr_valid & _GEN_319
    & ~ldq_3_bits_addr_is_virtual & _GEN_320[0] & dword_addr_matches_3_0
    & (|_mask_overlap_T_6);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_322 =
    do_ld_search_0 & ldq_3_valid & ldq_3_bits_addr_valid & ~ldq_3_bits_addr_is_virtual
    & dword_addr_matches_3_0 & (|_mask_overlap_T_6);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_3 =
    lcam_ldq_idx_0 < 4'h3 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[3:2]));	// lsu.scala:215:29, :305:44, :1036:26, util.scala:351:72, :363:{52,64,72,78}
  wire              _GEN_323 = lcam_ldq_idx_0 != 4'h3;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_3;	// lsu.scala:1128:57
  wire              _GEN_324 = ~_GEN_318 | nacking_loads_3 | older_nacked_REG_3;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_325 = _GEN_317 | _GEN_321;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_3;	// lsu.scala:1131:58
  wire              _GEN_326 =
    _GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_62 = 15'h1 << ldq_4_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_66 = 15'h3 << {12'h0, ldq_4_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_327 =
    {{8'hFF},
     {ldq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_66[7:0]},
     {_l_mask_mask_T_62[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_4_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h4;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_4_0 =
    lcam_addr_0[39:6] == ldq_4_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_4_0 =
    block_addr_matches_4_0 & lcam_addr_0[5:3] == ldq_4_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_8 = _GEN_327[ldq_4_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_328 =
    fired_release_0 & ldq_4_valid & ldq_4_bits_addr_valid & block_addr_matches_4_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_329 = ldq_4_bits_executed | ldq_4_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_330 = _GEN_329 | l_forwarders_4_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_331 = ldq_4_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_332 =
    do_st_search_0 & ldq_4_valid & ldq_4_bits_addr_valid & _GEN_330
    & ~ldq_4_bits_addr_is_virtual & _GEN_331[0] & dword_addr_matches_4_0
    & (|_mask_overlap_T_8);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_333 =
    do_ld_search_0 & ldq_4_valid & ldq_4_bits_addr_valid & ~ldq_4_bits_addr_is_virtual
    & dword_addr_matches_4_0 & (|_mask_overlap_T_8);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_4 =
    lcam_ldq_idx_0 < 4'h4 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'h4;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_334 = lcam_ldq_idx_0 != 4'h4;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_4;	// lsu.scala:1128:57
  wire              _GEN_335 = ~_GEN_329 | nacking_loads_4 | older_nacked_REG_4;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_336 = _GEN_328 | _GEN_332;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_4;	// lsu.scala:1131:58
  wire              _GEN_337 =
    _GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_77 = 15'h1 << ldq_5_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_81 = 15'h3 << {12'h0, ldq_5_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_338 =
    {{8'hFF},
     {ldq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_81[7:0]},
     {_l_mask_mask_T_77[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_5_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h5;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_5_0 =
    lcam_addr_0[39:6] == ldq_5_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_5_0 =
    block_addr_matches_5_0 & lcam_addr_0[5:3] == ldq_5_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_10 = _GEN_338[ldq_5_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_339 =
    fired_release_0 & ldq_5_valid & ldq_5_bits_addr_valid & block_addr_matches_5_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_340 = ldq_5_bits_executed | ldq_5_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_341 = _GEN_340 | l_forwarders_5_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_342 = ldq_5_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_343 =
    do_st_search_0 & ldq_5_valid & ldq_5_bits_addr_valid & _GEN_341
    & ~ldq_5_bits_addr_is_virtual & _GEN_342[0] & dword_addr_matches_5_0
    & (|_mask_overlap_T_10);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_344 =
    do_ld_search_0 & ldq_5_valid & ldq_5_bits_addr_valid & ~ldq_5_bits_addr_is_virtual
    & dword_addr_matches_5_0 & (|_mask_overlap_T_10);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_5 =
    lcam_ldq_idx_0 < 4'h5 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'h5;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_345 = lcam_ldq_idx_0 != 4'h5;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_5;	// lsu.scala:1128:57
  wire              _GEN_346 = ~_GEN_340 | nacking_loads_5 | older_nacked_REG_5;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_347 = _GEN_339 | _GEN_343;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_5;	// lsu.scala:1131:58
  wire              _GEN_348 =
    _GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_92 = 15'h1 << ldq_6_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_96 = 15'h3 << {12'h0, ldq_6_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_349 =
    {{8'hFF},
     {ldq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_96[7:0]},
     {_l_mask_mask_T_92[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_6_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h6;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_6_0 =
    lcam_addr_0[39:6] == ldq_6_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_6_0 =
    block_addr_matches_6_0 & lcam_addr_0[5:3] == ldq_6_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_12 = _GEN_349[ldq_6_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_350 =
    fired_release_0 & ldq_6_valid & ldq_6_bits_addr_valid & block_addr_matches_6_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_351 = ldq_6_bits_executed | ldq_6_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_352 = _GEN_351 | l_forwarders_6_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_353 = ldq_6_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_354 =
    do_st_search_0 & ldq_6_valid & ldq_6_bits_addr_valid & _GEN_352
    & ~ldq_6_bits_addr_is_virtual & _GEN_353[0] & dword_addr_matches_6_0
    & (|_mask_overlap_T_12);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_355 =
    do_ld_search_0 & ldq_6_valid & ldq_6_bits_addr_valid & ~ldq_6_bits_addr_is_virtual
    & dword_addr_matches_6_0 & (|_mask_overlap_T_12);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_6 =
    lcam_ldq_idx_0 < 4'h6 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'h6;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_356 = lcam_ldq_idx_0 != 4'h6;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_6;	// lsu.scala:1128:57
  wire              _GEN_357 = ~_GEN_351 | nacking_loads_6 | older_nacked_REG_6;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_358 = _GEN_350 | _GEN_354;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_6;	// lsu.scala:1131:58
  wire              _GEN_359 =
    _GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_107 = 15'h1 << ldq_7_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_111 =
    15'h3 << {12'h0, ldq_7_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_360 =
    {{8'hFF},
     {ldq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_111[7:0]},
     {_l_mask_mask_T_107[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_7_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h7;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_7_0 =
    lcam_addr_0[39:6] == ldq_7_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_7_0 =
    block_addr_matches_7_0 & lcam_addr_0[5:3] == ldq_7_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_14 = _GEN_360[ldq_7_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_361 =
    fired_release_0 & ldq_7_valid & ldq_7_bits_addr_valid & block_addr_matches_7_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_362 = ldq_7_bits_executed | ldq_7_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_363 = _GEN_362 | l_forwarders_7_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_364 = ldq_7_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_365 =
    do_st_search_0 & ldq_7_valid & ldq_7_bits_addr_valid & _GEN_363
    & ~ldq_7_bits_addr_is_virtual & _GEN_364[0] & dword_addr_matches_7_0
    & (|_mask_overlap_T_14);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_366 =
    do_ld_search_0 & ldq_7_valid & ldq_7_bits_addr_valid & ~ldq_7_bits_addr_is_virtual
    & dword_addr_matches_7_0 & (|_mask_overlap_T_14);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_7 =
    lcam_ldq_idx_0 < 4'h7 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head[3];	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_367 = lcam_ldq_idx_0 != 4'h7;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_7;	// lsu.scala:1128:57
  wire              _GEN_368 = ~_GEN_362 | nacking_loads_7 | older_nacked_REG_7;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_369 = _GEN_361 | _GEN_365;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_7;	// lsu.scala:1131:58
  wire              _GEN_370 =
    _GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_122 = 15'h1 << ldq_8_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_126 =
    15'h3 << {12'h0, ldq_8_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_371 =
    {{8'hFF},
     {ldq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_126[7:0]},
     {_l_mask_mask_T_122[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_8_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h8;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_8_0 =
    lcam_addr_0[39:6] == ldq_8_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_8_0 =
    block_addr_matches_8_0 & lcam_addr_0[5:3] == ldq_8_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_16 = _GEN_371[ldq_8_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_372 =
    fired_release_0 & ldq_8_valid & ldq_8_bits_addr_valid & block_addr_matches_8_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_373 = ldq_8_bits_executed | ldq_8_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_374 = _GEN_373 | l_forwarders_8_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_375 = ldq_8_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_376 =
    do_st_search_0 & ldq_8_valid & ldq_8_bits_addr_valid & _GEN_374
    & ~ldq_8_bits_addr_is_virtual & _GEN_375[0] & dword_addr_matches_8_0
    & (|_mask_overlap_T_16);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_377 =
    do_ld_search_0 & ldq_8_valid & ldq_8_bits_addr_valid & ~ldq_8_bits_addr_is_virtual
    & dword_addr_matches_8_0 & (|_mask_overlap_T_16);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_8 =
    lcam_ldq_idx_0[3] ^ lcam_ldq_idx_0 >= ldq_head ^ ldq_head > 4'h8;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_378 = lcam_ldq_idx_0 != 4'h8;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_8;	// lsu.scala:1128:57
  wire              _GEN_379 = ~_GEN_373 | nacking_loads_8 | older_nacked_REG_8;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_380 = _GEN_372 | _GEN_376;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_8;	// lsu.scala:1131:58
  wire              _GEN_381 =
    _GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_137 = 15'h1 << ldq_9_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_141 =
    15'h3 << {12'h0, ldq_9_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_382 =
    {{8'hFF},
     {ldq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_141[7:0]},
     {_l_mask_mask_T_137[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_9_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'h9;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_9_0 =
    lcam_addr_0[39:6] == ldq_9_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_9_0 =
    block_addr_matches_9_0 & lcam_addr_0[5:3] == ldq_9_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_18 = _GEN_382[ldq_9_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_383 =
    fired_release_0 & ldq_9_valid & ldq_9_bits_addr_valid & block_addr_matches_9_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_384 = ldq_9_bits_executed | ldq_9_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_385 = _GEN_384 | l_forwarders_9_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_386 = ldq_9_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_387 =
    do_st_search_0 & ldq_9_valid & ldq_9_bits_addr_valid & _GEN_385
    & ~ldq_9_bits_addr_is_virtual & _GEN_386[0] & dword_addr_matches_9_0
    & (|_mask_overlap_T_18);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_388 =
    do_ld_search_0 & ldq_9_valid & ldq_9_bits_addr_valid & ~ldq_9_bits_addr_is_virtual
    & dword_addr_matches_9_0 & (|_mask_overlap_T_18);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_9 =
    lcam_ldq_idx_0 < 4'h9 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'h9;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_389 = lcam_ldq_idx_0 != 4'h9;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_9;	// lsu.scala:1128:57
  wire              _GEN_390 = ~_GEN_384 | nacking_loads_9 | older_nacked_REG_9;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_391 = _GEN_383 | _GEN_387;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_9;	// lsu.scala:1131:58
  wire              _GEN_392 =
    _GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_152 = 15'h1 << ldq_10_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_156 =
    15'h3 << {12'h0, ldq_10_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_393 =
    {{8'hFF},
     {ldq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_156[7:0]},
     {_l_mask_mask_T_152[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_10_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'hA;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_10_0 =
    lcam_addr_0[39:6] == ldq_10_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_10_0 =
    block_addr_matches_10_0 & lcam_addr_0[5:3] == ldq_10_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_20 = _GEN_393[ldq_10_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_394 =
    fired_release_0 & ldq_10_valid & ldq_10_bits_addr_valid & block_addr_matches_10_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_395 = ldq_10_bits_executed | ldq_10_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_396 = _GEN_395 | l_forwarders_10_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_397 = ldq_10_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_398 =
    do_st_search_0 & ldq_10_valid & ldq_10_bits_addr_valid & _GEN_396
    & ~ldq_10_bits_addr_is_virtual & _GEN_397[0] & dword_addr_matches_10_0
    & (|_mask_overlap_T_20);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_399 =
    do_ld_search_0 & ldq_10_valid & ldq_10_bits_addr_valid & ~ldq_10_bits_addr_is_virtual
    & dword_addr_matches_10_0 & (|_mask_overlap_T_20);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_10 =
    lcam_ldq_idx_0 < 4'hA ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'hA;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_400 = lcam_ldq_idx_0 != 4'hA;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_10;	// lsu.scala:1128:57
  wire              _GEN_401 = ~_GEN_395 | nacking_loads_10 | older_nacked_REG_10;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_402 = _GEN_394 | _GEN_398;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_10;	// lsu.scala:1131:58
  wire              _GEN_403 =
    _GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_167 = 15'h1 << ldq_11_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_171 =
    15'h3 << {12'h0, ldq_11_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_404 =
    {{8'hFF},
     {ldq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_171[7:0]},
     {_l_mask_mask_T_167[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_11_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'hB;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_11_0 =
    lcam_addr_0[39:6] == ldq_11_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_11_0 =
    block_addr_matches_11_0 & lcam_addr_0[5:3] == ldq_11_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_22 = _GEN_404[ldq_11_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_405 =
    fired_release_0 & ldq_11_valid & ldq_11_bits_addr_valid & block_addr_matches_11_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_406 = ldq_11_bits_executed | ldq_11_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_407 = _GEN_406 | l_forwarders_11_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_408 = ldq_11_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_409 =
    do_st_search_0 & ldq_11_valid & ldq_11_bits_addr_valid & _GEN_407
    & ~ldq_11_bits_addr_is_virtual & _GEN_408[0] & dword_addr_matches_11_0
    & (|_mask_overlap_T_22);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_410 =
    do_ld_search_0 & ldq_11_valid & ldq_11_bits_addr_valid & ~ldq_11_bits_addr_is_virtual
    & dword_addr_matches_11_0 & (|_mask_overlap_T_22);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_11 =
    lcam_ldq_idx_0 < 4'hB ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'hB;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_411 = lcam_ldq_idx_0 != 4'hB;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_11;	// lsu.scala:1128:57
  wire              _GEN_412 = ~_GEN_406 | nacking_loads_11 | older_nacked_REG_11;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_413 = _GEN_405 | _GEN_409;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_11;	// lsu.scala:1131:58
  wire              _GEN_414 =
    _GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_182 = 15'h1 << ldq_12_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_186 =
    15'h3 << {12'h0, ldq_12_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_415 =
    {{8'hFF},
     {ldq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_186[7:0]},
     {_l_mask_mask_T_182[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_12_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'hC;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_12_0 =
    lcam_addr_0[39:6] == ldq_12_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_12_0 =
    block_addr_matches_12_0 & lcam_addr_0[5:3] == ldq_12_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_24 = _GEN_415[ldq_12_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_416 =
    fired_release_0 & ldq_12_valid & ldq_12_bits_addr_valid & block_addr_matches_12_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_417 = ldq_12_bits_executed | ldq_12_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_418 = _GEN_417 | l_forwarders_12_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_419 = ldq_12_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_420 =
    do_st_search_0 & ldq_12_valid & ldq_12_bits_addr_valid & _GEN_418
    & ~ldq_12_bits_addr_is_virtual & _GEN_419[0] & dword_addr_matches_12_0
    & (|_mask_overlap_T_24);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_421 =
    do_ld_search_0 & ldq_12_valid & ldq_12_bits_addr_valid & ~ldq_12_bits_addr_is_virtual
    & dword_addr_matches_12_0 & (|_mask_overlap_T_24);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_12 =
    lcam_ldq_idx_0[3:2] != 2'h3 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'hC;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_422 = lcam_ldq_idx_0 != 4'hC;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_12;	// lsu.scala:1128:57
  wire              _GEN_423 = ~_GEN_417 | nacking_loads_12 | older_nacked_REG_12;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_424 = _GEN_416 | _GEN_420;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_12;	// lsu.scala:1131:58
  wire              _GEN_425 =
    _GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_197 = 15'h1 << ldq_13_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_201 =
    15'h3 << {12'h0, ldq_13_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_426 =
    {{8'hFF},
     {ldq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_201[7:0]},
     {_l_mask_mask_T_197[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_13_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'hD;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_13_0 =
    lcam_addr_0[39:6] == ldq_13_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_13_0 =
    block_addr_matches_13_0 & lcam_addr_0[5:3] == ldq_13_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_26 = _GEN_426[ldq_13_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_427 =
    fired_release_0 & ldq_13_valid & ldq_13_bits_addr_valid & block_addr_matches_13_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_428 = ldq_13_bits_executed | ldq_13_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_429 = _GEN_428 | l_forwarders_13_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_430 = ldq_13_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_431 =
    do_st_search_0 & ldq_13_valid & ldq_13_bits_addr_valid & _GEN_429
    & ~ldq_13_bits_addr_is_virtual & _GEN_430[0] & dword_addr_matches_13_0
    & (|_mask_overlap_T_26);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_432 =
    do_ld_search_0 & ldq_13_valid & ldq_13_bits_addr_valid & ~ldq_13_bits_addr_is_virtual
    & dword_addr_matches_13_0 & (|_mask_overlap_T_26);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_13 =
    lcam_ldq_idx_0 < 4'hD ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 4'hD;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,64,72,78}
  wire              _GEN_433 = lcam_ldq_idx_0 != 4'hD;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_13;	// lsu.scala:1128:57
  wire              _GEN_434 = ~_GEN_428 | nacking_loads_13 | older_nacked_REG_13;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_435 = _GEN_427 | _GEN_431;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_13;	// lsu.scala:1131:58
  wire              _GEN_436 =
    _GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_212 = 15'h1 << ldq_14_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_216 =
    15'h3 << {12'h0, ldq_14_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_437 =
    {{8'hFF},
     {ldq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_216[7:0]},
     {_l_mask_mask_T_212[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_14_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 4'hE;	// lsu.scala:305:44, :1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_14_0 =
    lcam_addr_0[39:6] == ldq_14_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_14_0 =
    block_addr_matches_14_0 & lcam_addr_0[5:3] == ldq_14_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_28 = _GEN_437[ldq_14_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_438 =
    fired_release_0 & ldq_14_valid & ldq_14_bits_addr_valid & block_addr_matches_14_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_439 = ldq_14_bits_executed | ldq_14_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_440 = _GEN_439 | l_forwarders_14_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_441 = ldq_14_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_442 =
    do_st_search_0 & ldq_14_valid & ldq_14_bits_addr_valid & _GEN_440
    & ~ldq_14_bits_addr_is_virtual & _GEN_441[0] & dword_addr_matches_14_0
    & (|_mask_overlap_T_28);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_443 =
    do_ld_search_0 & ldq_14_valid & ldq_14_bits_addr_valid & ~ldq_14_bits_addr_is_virtual
    & dword_addr_matches_14_0 & (|_mask_overlap_T_28);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_14 =
    lcam_ldq_idx_0[3:1] != 3'h7 ^ lcam_ldq_idx_0 < ldq_head ^ (&ldq_head);	// lsu.scala:215:29, :1036:26, util.scala:351:72, :363:{52,64,72,78}
  wire              _GEN_444 = lcam_ldq_idx_0 != 4'hE;	// lsu.scala:305:44, :1036:26, :1125:38
  reg               older_nacked_REG_14;	// lsu.scala:1128:57
  wire              _GEN_445 = ~_GEN_439 | nacking_loads_14 | older_nacked_REG_14;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_446 = _GEN_438 | _GEN_442;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_14;	// lsu.scala:1131:58
  wire              _GEN_447 =
    _GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445);	// lsu.scala:1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1131:48, util.scala:363:72
  wire [14:0]       _l_mask_mask_T_227 = 15'h1 << ldq_15_bits_addr_bits[2:0];	// lsu.scala:210:16, :1663:{48,55}
  wire [14:0]       _l_mask_mask_T_231 =
    15'h3 << {12'h0, ldq_15_bits_addr_bits[2:1], 1'h0};	// lsu.scala:210:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_448 =
    {{8'hFF},
     {ldq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_l_mask_mask_T_231[7:0]},
     {_l_mask_mask_T_227[7:0]}};	// Mux.scala:98:16, lsu.scala:210:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              l_forwarders_15_0 = wb_forward_valid_0 & (&wb_forward_ldq_idx_0);	// lsu.scala:1064:36, :1065:36, :1075:{63,88}
  wire              block_addr_matches_15_0 =
    lcam_addr_0[39:6] == ldq_15_bits_addr_bits[39:6];	// lsu.scala:210:16, :1025:37, :1080:{57,73,84}
  wire              dword_addr_matches_15_0 =
    block_addr_matches_15_0 & lcam_addr_0[5:3] == ldq_15_bits_addr_bits[5:3];	// lsu.scala:210:16, :1025:37, :1080:73, :1081:{66,81,100,110}
  wire [7:0]        _mask_overlap_T_30 = _GEN_448[ldq_15_bits_uop_mem_size] & lcam_mask_0;	// Mux.scala:98:16, lsu.scala:210:16, :1082:46, :1663:26, :1664:26, :1665:26
  wire              _GEN_449 =
    fired_release_0 & ldq_15_valid & ldq_15_bits_addr_valid & block_addr_matches_15_0;	// lsu.scala:210:16, :900:37, :1080:73, :1090:34
  wire              _GEN_450 = ldq_15_bits_executed | ldq_15_bits_succeeded;	// lsu.scala:210:16, :1098:37
  wire              _GEN_451 = _GEN_450 | l_forwarders_15_0;	// lsu.scala:1075:63, :1098:{37,57}
  wire [15:0]       _GEN_452 = ldq_15_bits_st_dep_mask >> _GEN_287;	// lsu.scala:210:16, :1100:38
  wire              _GEN_453 =
    do_st_search_0 & ldq_15_valid & ldq_15_bits_addr_valid & _GEN_451
    & ~ldq_15_bits_addr_is_virtual & _GEN_452[0] & dword_addr_matches_15_0
    & (|_mask_overlap_T_30);	// lsu.scala:210:16, :433:52, :1014:108, :1081:66, :1082:46, :1083:62, :1098:57, :1100:38, :1101:131
  wire              _GEN_454 =
    do_ld_search_0 & ldq_15_valid & ldq_15_bits_addr_valid & ~ldq_15_bits_addr_is_virtual
    & dword_addr_matches_15_0 & (|_mask_overlap_T_30);	// lsu.scala:210:16, :433:52, :1016:106, :1081:66, :1082:46, :1083:62, :1115:47
  wire              searcher_is_older_15 =
    lcam_ldq_idx_0 != 4'hF ^ lcam_ldq_idx_0 < ldq_head;	// lsu.scala:215:29, :305:44, :1036:26, util.scala:363:{52,58,64}
  reg               older_nacked_REG_15;	// lsu.scala:1128:57
  wire              _GEN_455 = ~_GEN_450 | nacking_loads_15 | older_nacked_REG_15;	// lsu.scala:1098:37, :1128:57, :1129:{17,56}, :1284:5, :1287:7
  wire              _GEN_456 = _GEN_449 | _GEN_453;	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1116:37
  reg               io_dmem_s1_kill_0_REG_15;	// lsu.scala:1131:58
  wire              _GEN_457 =
    _GEN_456 | ~_GEN_454 | searcher_is_older_15 | ~(~(&lcam_ldq_idx_0) & _GEN_455);	// lsu.scala:1036:26, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, :1131:48, util.scala:363:58
  wire              _GEN_458 =
    _GEN_457
      ? (_GEN_447
           ? (_GEN_436
                ? (_GEN_425
                     ? (_GEN_414
                          ? (_GEN_403
                               ? (_GEN_392
                                    ? (_GEN_381
                                         ? (_GEN_370
                                              ? (_GEN_359
                                                   ? (_GEN_348
                                                        ? (_GEN_337
                                                             ? (_GEN_326
                                                                  ? (_GEN_315
                                                                       ? (_GEN_304
                                                                            ? ~_GEN_292
                                                                              & _GEN_290
                                                                              & ~searcher_is_older
                                                                              & _GEN_293
                                                                              & io_dmem_s1_kill_0_REG
                                                                            : io_dmem_s1_kill_0_REG_1)
                                                                       : io_dmem_s1_kill_0_REG_2)
                                                                  : io_dmem_s1_kill_0_REG_3)
                                                             : io_dmem_s1_kill_0_REG_4)
                                                        : io_dmem_s1_kill_0_REG_5)
                                                   : io_dmem_s1_kill_0_REG_6)
                                              : io_dmem_s1_kill_0_REG_7)
                                         : io_dmem_s1_kill_0_REG_8)
                                    : io_dmem_s1_kill_0_REG_9)
                               : io_dmem_s1_kill_0_REG_10)
                          : io_dmem_s1_kill_0_REG_11)
                     : io_dmem_s1_kill_0_REG_12)
                : io_dmem_s1_kill_0_REG_13)
           : io_dmem_s1_kill_0_REG_14)
      : io_dmem_s1_kill_0_REG_15;	// lsu.scala:764:24, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:47, :1129:73, :1131:{48,58}, util.scala:363:72
  wire              can_forward_0 =
    _GEN_457 & _GEN_447 & _GEN_436 & _GEN_425 & _GEN_414 & _GEN_403 & _GEN_392 & _GEN_381
    & _GEN_370 & _GEN_359 & _GEN_348 & _GEN_337 & _GEN_326 & _GEN_315 & _GEN_304
    & (_GEN_292 | ~_GEN_290 | searcher_is_older | ~_GEN_293)
    & (_can_forward_T ? ~mem_tlb_uncacheable_0 : ~_GEN_204[lcam_ldq_idx_0]);	// lsu.scala:502:88, :764:24, :926:41, :1016:61, :1036:26, :1045:{8,56}, :1046:7, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:47, :1129:73, :1131:48, :1132:48, util.scala:363:72
  wire              dword_addr_matches_16_0 =
    stq_0_bits_addr_valid & ~stq_0_bits_addr_is_virtual
    & stq_0_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_2 = 15'h1 << stq_0_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_6 =
    15'h3 << {12'h0, stq_0_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_459 =
    {{8'hFF},
     {stq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_6[7:0]},
     {_write_mask_mask_T_2[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_460 = do_ld_search_0 & stq_0_valid & lcam_st_dep_mask_0[0];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_461 = lcam_mask_0 & _GEN_459[stq_0_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_462 =
    _GEN_461 == lcam_mask_0 & ~stq_0_bits_uop_is_fence & dword_addr_matches_16_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_16;	// lsu.scala:1153:56
  wire              _GEN_463 = (|_GEN_461) & dword_addr_matches_16_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_17;	// lsu.scala:1159:56
  wire              _GEN_464 = stq_0_bits_uop_is_fence | stq_0_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_0 = _GEN_460 & (_GEN_462 | _GEN_463 | _GEN_464);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_18;	// lsu.scala:1165:56
  wire              _GEN_465 =
    _GEN_460
      ? (_GEN_462
           ? io_dmem_s1_kill_0_REG_16
           : _GEN_463
               ? io_dmem_s1_kill_0_REG_17
               : _GEN_464 ? io_dmem_s1_kill_0_REG_18 : _GEN_458)
      : _GEN_458;	// lsu.scala:1091:36, :1102:37, :1116:37, :1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_17_0 =
    stq_1_bits_addr_valid & ~stq_1_bits_addr_is_virtual
    & stq_1_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_17 = 15'h1 << stq_1_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_21 =
    15'h3 << {12'h0, stq_1_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_466 =
    {{8'hFF},
     {stq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_21[7:0]},
     {_write_mask_mask_T_17[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_467 = do_ld_search_0 & stq_1_valid & lcam_st_dep_mask_0[1];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_468 = lcam_mask_0 & _GEN_466[stq_1_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_469 =
    _GEN_468 == lcam_mask_0 & ~stq_1_bits_uop_is_fence & dword_addr_matches_17_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_19;	// lsu.scala:1153:56
  wire              _GEN_470 = (|_GEN_468) & dword_addr_matches_17_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_20;	// lsu.scala:1159:56
  wire              _GEN_471 = stq_1_bits_uop_is_fence | stq_1_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_1 = _GEN_467 & (_GEN_469 | _GEN_470 | _GEN_471);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_21;	// lsu.scala:1165:56
  wire              _GEN_472 =
    _GEN_467
      ? (_GEN_469
           ? io_dmem_s1_kill_0_REG_19
           : _GEN_470
               ? io_dmem_s1_kill_0_REG_20
               : _GEN_471 ? io_dmem_s1_kill_0_REG_21 : _GEN_465)
      : _GEN_465;	// lsu.scala:1091:36, :1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_18_0 =
    stq_2_bits_addr_valid & ~stq_2_bits_addr_is_virtual
    & stq_2_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_32 = 15'h1 << stq_2_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_36 =
    15'h3 << {12'h0, stq_2_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_473 =
    {{8'hFF},
     {stq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_36[7:0]},
     {_write_mask_mask_T_32[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_474 = do_ld_search_0 & stq_2_valid & lcam_st_dep_mask_0[2];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_475 = lcam_mask_0 & _GEN_473[stq_2_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_476 =
    _GEN_475 == lcam_mask_0 & ~stq_2_bits_uop_is_fence & dword_addr_matches_18_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_22;	// lsu.scala:1153:56
  wire              _GEN_477 = (|_GEN_475) & dword_addr_matches_18_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_23;	// lsu.scala:1159:56
  wire              _GEN_478 = stq_2_bits_uop_is_fence | stq_2_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_2 = _GEN_474 & (_GEN_476 | _GEN_477 | _GEN_478);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_24;	// lsu.scala:1165:56
  wire              _GEN_479 =
    _GEN_474
      ? (_GEN_476
           ? io_dmem_s1_kill_0_REG_22
           : _GEN_477
               ? io_dmem_s1_kill_0_REG_23
               : _GEN_478 ? io_dmem_s1_kill_0_REG_24 : _GEN_472)
      : _GEN_472;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_19_0 =
    stq_3_bits_addr_valid & ~stq_3_bits_addr_is_virtual
    & stq_3_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_47 = 15'h1 << stq_3_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_51 =
    15'h3 << {12'h0, stq_3_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_480 =
    {{8'hFF},
     {stq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_51[7:0]},
     {_write_mask_mask_T_47[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_481 = do_ld_search_0 & stq_3_valid & lcam_st_dep_mask_0[3];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_482 = lcam_mask_0 & _GEN_480[stq_3_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_483 =
    _GEN_482 == lcam_mask_0 & ~stq_3_bits_uop_is_fence & dword_addr_matches_19_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_25;	// lsu.scala:1153:56
  wire              _GEN_484 = (|_GEN_482) & dword_addr_matches_19_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_26;	// lsu.scala:1159:56
  wire              _GEN_485 = stq_3_bits_uop_is_fence | stq_3_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_3 = _GEN_481 & (_GEN_483 | _GEN_484 | _GEN_485);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_27;	// lsu.scala:1165:56
  wire              _GEN_486 =
    _GEN_481
      ? (_GEN_483
           ? io_dmem_s1_kill_0_REG_25
           : _GEN_484
               ? io_dmem_s1_kill_0_REG_26
               : _GEN_485 ? io_dmem_s1_kill_0_REG_27 : _GEN_479)
      : _GEN_479;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_20_0 =
    stq_4_bits_addr_valid & ~stq_4_bits_addr_is_virtual
    & stq_4_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_62 = 15'h1 << stq_4_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_66 =
    15'h3 << {12'h0, stq_4_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_487 =
    {{8'hFF},
     {stq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_66[7:0]},
     {_write_mask_mask_T_62[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_488 = do_ld_search_0 & stq_4_valid & lcam_st_dep_mask_0[4];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_489 = lcam_mask_0 & _GEN_487[stq_4_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_490 =
    _GEN_489 == lcam_mask_0 & ~stq_4_bits_uop_is_fence & dword_addr_matches_20_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_28;	// lsu.scala:1153:56
  wire              _GEN_491 = (|_GEN_489) & dword_addr_matches_20_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_29;	// lsu.scala:1159:56
  wire              _GEN_492 = stq_4_bits_uop_is_fence | stq_4_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_4 = _GEN_488 & (_GEN_490 | _GEN_491 | _GEN_492);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_30;	// lsu.scala:1165:56
  wire              _GEN_493 =
    _GEN_488
      ? (_GEN_490
           ? io_dmem_s1_kill_0_REG_28
           : _GEN_491
               ? io_dmem_s1_kill_0_REG_29
               : _GEN_492 ? io_dmem_s1_kill_0_REG_30 : _GEN_486)
      : _GEN_486;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_21_0 =
    stq_5_bits_addr_valid & ~stq_5_bits_addr_is_virtual
    & stq_5_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_77 = 15'h1 << stq_5_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_81 =
    15'h3 << {12'h0, stq_5_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_494 =
    {{8'hFF},
     {stq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_81[7:0]},
     {_write_mask_mask_T_77[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_495 = do_ld_search_0 & stq_5_valid & lcam_st_dep_mask_0[5];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_496 = lcam_mask_0 & _GEN_494[stq_5_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_497 =
    _GEN_496 == lcam_mask_0 & ~stq_5_bits_uop_is_fence & dword_addr_matches_21_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_31;	// lsu.scala:1153:56
  wire              _GEN_498 = (|_GEN_496) & dword_addr_matches_21_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_32;	// lsu.scala:1159:56
  wire              _GEN_499 = stq_5_bits_uop_is_fence | stq_5_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_5 = _GEN_495 & (_GEN_497 | _GEN_498 | _GEN_499);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_33;	// lsu.scala:1165:56
  wire              _GEN_500 =
    _GEN_495
      ? (_GEN_497
           ? io_dmem_s1_kill_0_REG_31
           : _GEN_498
               ? io_dmem_s1_kill_0_REG_32
               : _GEN_499 ? io_dmem_s1_kill_0_REG_33 : _GEN_493)
      : _GEN_493;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_22_0 =
    stq_6_bits_addr_valid & ~stq_6_bits_addr_is_virtual
    & stq_6_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_92 = 15'h1 << stq_6_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_96 =
    15'h3 << {12'h0, stq_6_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_501 =
    {{8'hFF},
     {stq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_96[7:0]},
     {_write_mask_mask_T_92[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_502 = do_ld_search_0 & stq_6_valid & lcam_st_dep_mask_0[6];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_503 = lcam_mask_0 & _GEN_501[stq_6_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_504 =
    _GEN_503 == lcam_mask_0 & ~stq_6_bits_uop_is_fence & dword_addr_matches_22_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_34;	// lsu.scala:1153:56
  wire              _GEN_505 = (|_GEN_503) & dword_addr_matches_22_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_35;	// lsu.scala:1159:56
  wire              _GEN_506 = stq_6_bits_uop_is_fence | stq_6_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_6 = _GEN_502 & (_GEN_504 | _GEN_505 | _GEN_506);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_36;	// lsu.scala:1165:56
  wire              _GEN_507 =
    _GEN_502
      ? (_GEN_504
           ? io_dmem_s1_kill_0_REG_34
           : _GEN_505
               ? io_dmem_s1_kill_0_REG_35
               : _GEN_506 ? io_dmem_s1_kill_0_REG_36 : _GEN_500)
      : _GEN_500;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_23_0 =
    stq_7_bits_addr_valid & ~stq_7_bits_addr_is_virtual
    & stq_7_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_107 = 15'h1 << stq_7_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_111 =
    15'h3 << {12'h0, stq_7_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_508 =
    {{8'hFF},
     {stq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_111[7:0]},
     {_write_mask_mask_T_107[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_509 = do_ld_search_0 & stq_7_valid & lcam_st_dep_mask_0[7];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_510 = lcam_mask_0 & _GEN_508[stq_7_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_511 =
    _GEN_510 == lcam_mask_0 & ~stq_7_bits_uop_is_fence & dword_addr_matches_23_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_37;	// lsu.scala:1153:56
  wire              _GEN_512 = (|_GEN_510) & dword_addr_matches_23_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_38;	// lsu.scala:1159:56
  wire              _GEN_513 = stq_7_bits_uop_is_fence | stq_7_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_7 = _GEN_509 & (_GEN_511 | _GEN_512 | _GEN_513);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_39;	// lsu.scala:1165:56
  wire              _GEN_514 =
    _GEN_509
      ? (_GEN_511
           ? io_dmem_s1_kill_0_REG_37
           : _GEN_512
               ? io_dmem_s1_kill_0_REG_38
               : _GEN_513 ? io_dmem_s1_kill_0_REG_39 : _GEN_507)
      : _GEN_507;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_24_0 =
    stq_8_bits_addr_valid & ~stq_8_bits_addr_is_virtual
    & stq_8_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_122 = 15'h1 << stq_8_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_126 =
    15'h3 << {12'h0, stq_8_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_515 =
    {{8'hFF},
     {stq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_126[7:0]},
     {_write_mask_mask_T_122[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_516 = do_ld_search_0 & stq_8_valid & lcam_st_dep_mask_0[8];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_517 = lcam_mask_0 & _GEN_515[stq_8_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_518 =
    _GEN_517 == lcam_mask_0 & ~stq_8_bits_uop_is_fence & dword_addr_matches_24_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_40;	// lsu.scala:1153:56
  wire              _GEN_519 = (|_GEN_517) & dword_addr_matches_24_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_41;	// lsu.scala:1159:56
  wire              _GEN_520 = stq_8_bits_uop_is_fence | stq_8_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_8 = _GEN_516 & (_GEN_518 | _GEN_519 | _GEN_520);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_42;	// lsu.scala:1165:56
  wire              _GEN_521 =
    _GEN_516
      ? (_GEN_518
           ? io_dmem_s1_kill_0_REG_40
           : _GEN_519
               ? io_dmem_s1_kill_0_REG_41
               : _GEN_520 ? io_dmem_s1_kill_0_REG_42 : _GEN_514)
      : _GEN_514;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_25_0 =
    stq_9_bits_addr_valid & ~stq_9_bits_addr_is_virtual
    & stq_9_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_137 = 15'h1 << stq_9_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_141 =
    15'h3 << {12'h0, stq_9_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_522 =
    {{8'hFF},
     {stq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_141[7:0]},
     {_write_mask_mask_T_137[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_523 = do_ld_search_0 & stq_9_valid & lcam_st_dep_mask_0[9];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_524 = lcam_mask_0 & _GEN_522[stq_9_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_525 =
    _GEN_524 == lcam_mask_0 & ~stq_9_bits_uop_is_fence & dword_addr_matches_25_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_43;	// lsu.scala:1153:56
  wire              _GEN_526 = (|_GEN_524) & dword_addr_matches_25_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_44;	// lsu.scala:1159:56
  wire              _GEN_527 = stq_9_bits_uop_is_fence | stq_9_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_9 = _GEN_523 & (_GEN_525 | _GEN_526 | _GEN_527);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_45;	// lsu.scala:1165:56
  wire              _GEN_528 =
    _GEN_523
      ? (_GEN_525
           ? io_dmem_s1_kill_0_REG_43
           : _GEN_526
               ? io_dmem_s1_kill_0_REG_44
               : _GEN_527 ? io_dmem_s1_kill_0_REG_45 : _GEN_521)
      : _GEN_521;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_26_0 =
    stq_10_bits_addr_valid & ~stq_10_bits_addr_is_virtual
    & stq_10_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_152 = 15'h1 << stq_10_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_156 =
    15'h3 << {12'h0, stq_10_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_529 =
    {{8'hFF},
     {stq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_156[7:0]},
     {_write_mask_mask_T_152[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_530 = do_ld_search_0 & stq_10_valid & lcam_st_dep_mask_0[10];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_531 = lcam_mask_0 & _GEN_529[stq_10_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_532 =
    _GEN_531 == lcam_mask_0 & ~stq_10_bits_uop_is_fence & dword_addr_matches_26_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_46;	// lsu.scala:1153:56
  wire              _GEN_533 = (|_GEN_531) & dword_addr_matches_26_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_47;	// lsu.scala:1159:56
  wire              _GEN_534 = stq_10_bits_uop_is_fence | stq_10_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_10 = _GEN_530 & (_GEN_532 | _GEN_533 | _GEN_534);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_48;	// lsu.scala:1165:56
  wire              _GEN_535 =
    _GEN_530
      ? (_GEN_532
           ? io_dmem_s1_kill_0_REG_46
           : _GEN_533
               ? io_dmem_s1_kill_0_REG_47
               : _GEN_534 ? io_dmem_s1_kill_0_REG_48 : _GEN_528)
      : _GEN_528;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_27_0 =
    stq_11_bits_addr_valid & ~stq_11_bits_addr_is_virtual
    & stq_11_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_167 = 15'h1 << stq_11_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_171 =
    15'h3 << {12'h0, stq_11_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_536 =
    {{8'hFF},
     {stq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_171[7:0]},
     {_write_mask_mask_T_167[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_537 = do_ld_search_0 & stq_11_valid & lcam_st_dep_mask_0[11];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_538 = lcam_mask_0 & _GEN_536[stq_11_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_539 =
    _GEN_538 == lcam_mask_0 & ~stq_11_bits_uop_is_fence & dword_addr_matches_27_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_49;	// lsu.scala:1153:56
  wire              _GEN_540 = (|_GEN_538) & dword_addr_matches_27_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_50;	// lsu.scala:1159:56
  wire              _GEN_541 = stq_11_bits_uop_is_fence | stq_11_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_11 = _GEN_537 & (_GEN_539 | _GEN_540 | _GEN_541);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_51;	// lsu.scala:1165:56
  wire              _GEN_542 =
    _GEN_537
      ? (_GEN_539
           ? io_dmem_s1_kill_0_REG_49
           : _GEN_540
               ? io_dmem_s1_kill_0_REG_50
               : _GEN_541 ? io_dmem_s1_kill_0_REG_51 : _GEN_535)
      : _GEN_535;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_28_0 =
    stq_12_bits_addr_valid & ~stq_12_bits_addr_is_virtual
    & stq_12_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_182 = 15'h1 << stq_12_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_186 =
    15'h3 << {12'h0, stq_12_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_543 =
    {{8'hFF},
     {stq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_186[7:0]},
     {_write_mask_mask_T_182[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_544 = do_ld_search_0 & stq_12_valid & lcam_st_dep_mask_0[12];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_545 = lcam_mask_0 & _GEN_543[stq_12_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_546 =
    _GEN_545 == lcam_mask_0 & ~stq_12_bits_uop_is_fence & dword_addr_matches_28_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_52;	// lsu.scala:1153:56
  wire              _GEN_547 = (|_GEN_545) & dword_addr_matches_28_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_53;	// lsu.scala:1159:56
  wire              _GEN_548 = stq_12_bits_uop_is_fence | stq_12_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_12 = _GEN_544 & (_GEN_546 | _GEN_547 | _GEN_548);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_54;	// lsu.scala:1165:56
  wire              _GEN_549 =
    _GEN_544
      ? (_GEN_546
           ? io_dmem_s1_kill_0_REG_52
           : _GEN_547
               ? io_dmem_s1_kill_0_REG_53
               : _GEN_548 ? io_dmem_s1_kill_0_REG_54 : _GEN_542)
      : _GEN_542;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_29_0 =
    stq_13_bits_addr_valid & ~stq_13_bits_addr_is_virtual
    & stq_13_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_197 = 15'h1 << stq_13_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_201 =
    15'h3 << {12'h0, stq_13_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_550 =
    {{8'hFF},
     {stq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_201[7:0]},
     {_write_mask_mask_T_197[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_551 = do_ld_search_0 & stq_13_valid & lcam_st_dep_mask_0[13];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_552 = lcam_mask_0 & _GEN_550[stq_13_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_553 =
    _GEN_552 == lcam_mask_0 & ~stq_13_bits_uop_is_fence & dword_addr_matches_29_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_55;	// lsu.scala:1153:56
  wire              _GEN_554 = (|_GEN_552) & dword_addr_matches_29_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_56;	// lsu.scala:1159:56
  wire              _GEN_555 = stq_13_bits_uop_is_fence | stq_13_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_13 = _GEN_551 & (_GEN_553 | _GEN_554 | _GEN_555);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_57;	// lsu.scala:1165:56
  wire              _GEN_556 =
    _GEN_551
      ? (_GEN_553
           ? io_dmem_s1_kill_0_REG_55
           : _GEN_554
               ? io_dmem_s1_kill_0_REG_56
               : _GEN_555 ? io_dmem_s1_kill_0_REG_57 : _GEN_549)
      : _GEN_549;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_30_0 =
    stq_14_bits_addr_valid & ~stq_14_bits_addr_is_virtual
    & stq_14_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_212 = 15'h1 << stq_14_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_216 =
    15'h3 << {12'h0, stq_14_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_557 =
    {{8'hFF},
     {stq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_216[7:0]},
     {_write_mask_mask_T_212[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_558 = do_ld_search_0 & stq_14_valid & lcam_st_dep_mask_0[14];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_559 = lcam_mask_0 & _GEN_557[stq_14_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_560 =
    _GEN_559 == lcam_mask_0 & ~stq_14_bits_uop_is_fence & dword_addr_matches_30_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_58;	// lsu.scala:1153:56
  wire              _GEN_561 = (|_GEN_559) & dword_addr_matches_30_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_59;	// lsu.scala:1159:56
  wire              _GEN_562 = stq_14_bits_uop_is_fence | stq_14_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_14 = _GEN_558 & (_GEN_560 | _GEN_561 | _GEN_562);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_60;	// lsu.scala:1165:56
  wire              _GEN_563 =
    _GEN_558
      ? (_GEN_560
           ? io_dmem_s1_kill_0_REG_58
           : _GEN_561
               ? io_dmem_s1_kill_0_REG_59
               : _GEN_562 ? io_dmem_s1_kill_0_REG_60 : _GEN_556)
      : _GEN_556;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  wire              dword_addr_matches_31_0 =
    stq_15_bits_addr_valid & ~stq_15_bits_addr_is_virtual
    & stq_15_bits_addr_bits[31:3] == lcam_addr_0[31:3];	// lsu.scala:211:16, :1025:37, :1144:{31,60}, :1145:{38,58,74}
  wire [14:0]       _write_mask_mask_T_227 = 15'h1 << stq_15_bits_addr_bits[2:0];	// lsu.scala:211:16, :1663:{48,55}
  wire [14:0]       _write_mask_mask_T_231 =
    15'h3 << {12'h0, stq_15_bits_addr_bits[2:1], 1'h0};	// lsu.scala:211:16, :249:20, :708:86, :1664:{48,56}
  wire [3:0][7:0]   _GEN_564 =
    {{8'hFF},
     {stq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF},
     {_write_mask_mask_T_231[7:0]},
     {_write_mask_mask_T_227[7:0]}};	// Mux.scala:98:16, lsu.scala:211:16, :1663:{26,48}, :1664:{26,48}, :1665:{26,41,46}
  wire              _GEN_565 = do_ld_search_0 & stq_15_valid & lcam_st_dep_mask_0[15];	// lsu.scala:211:16, :915:33, :1016:106, :1148:{45,67}
  wire [7:0]        _GEN_566 = lcam_mask_0 & _GEN_564[stq_15_bits_uop_mem_size];	// Mux.scala:98:16, lsu.scala:211:16, :1149:30, :1663:26, :1664:26, :1665:26
  wire              _GEN_567 =
    _GEN_566 == lcam_mask_0 & ~stq_15_bits_uop_is_fence & dword_addr_matches_31_0
    & can_forward_0;	// Mux.scala:98:16, lsu.scala:211:16, :1091:36, :1102:37, :1116:37, :1144:60, :1149:{30,44,65,106}
  reg               io_dmem_s1_kill_0_REG_61;	// lsu.scala:1153:56
  wire              _GEN_568 = (|_GEN_566) & dword_addr_matches_31_0;	// lsu.scala:1144:60, :1149:30, :1156:{51,60}
  reg               io_dmem_s1_kill_0_REG_62;	// lsu.scala:1159:56
  wire              _GEN_569 = stq_15_bits_uop_is_fence | stq_15_bits_uop_is_amo;	// lsu.scala:211:16, :1162:37
  wire              ldst_addr_matches_0_15 = _GEN_565 & (_GEN_567 | _GEN_568 | _GEN_569);	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1151:46, :1156:60, :1157:9, :1158:46, :1162:37, :1163:9
  reg               io_dmem_s1_kill_0_REG_63;	// lsu.scala:1165:56
  reg               REG_1;	// lsu.scala:1189:64
  reg               REG_2;	// lsu.scala:1199:18
  reg  [3:0]        store_blocked_counter;	// lsu.scala:1204:36
  assign block_load_wakeup = (&store_blocked_counter) | REG_2;	// lsu.scala:1199:{18,80}, :1204:36, :1210:{33,43}, :1211:25
  reg               r_xcpt_valid;	// lsu.scala:1235:29
  reg  [11:0]       r_xcpt_uop_br_mask;	// lsu.scala:1236:25
  reg  [5:0]        r_xcpt_uop_rob_idx;	// lsu.scala:1236:25
  reg  [4:0]        r_xcpt_cause;	// lsu.scala:1236:25
  reg  [39:0]       r_xcpt_badvaddr;	// lsu.scala:1236:25
  wire              _io_core_spec_ld_wakeup_0_valid_output =
    fired_load_incoming_REG & ~mem_incoming_uop_0_fp_val & (|mem_incoming_uop_0_pdst);	// lsu.scala:894:51, :908:37, :1260:{40,69}, :1261:65
  wire              _GEN_570 = io_dmem_nack_0_valid & io_dmem_nack_0_bits_is_hella;	// lsu.scala:1287:7
  wire              _GEN_571 = hella_state == 3'h4;	// lsu.scala:242:38, :1288:28, util.scala:351:72
  wire              _GEN_572 = hella_state == 3'h6;	// lsu.scala:242:38, :1288:54, util.scala:351:72
  wire              _GEN_573 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h0;	// lsu.scala:1293:62
  wire              _GEN_574 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h1;	// lsu.scala:305:44, :1293:62
  wire              _GEN_575 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h2;	// lsu.scala:305:44, :1293:62
  wire              _GEN_576 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h3;	// lsu.scala:305:44, :1293:62
  wire              _GEN_577 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h4;	// lsu.scala:305:44, :1293:62
  wire              _GEN_578 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h5;	// lsu.scala:305:44, :1293:62
  wire              _GEN_579 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h6;	// lsu.scala:305:44, :1293:62
  wire              _GEN_580 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h7;	// lsu.scala:305:44, :1293:62
  wire              _GEN_581 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h8;	// lsu.scala:305:44, :1293:62
  wire              _GEN_582 = io_dmem_nack_0_bits_uop_ldq_idx == 4'h9;	// lsu.scala:305:44, :1293:62
  wire              _GEN_583 = io_dmem_nack_0_bits_uop_ldq_idx == 4'hA;	// lsu.scala:305:44, :1293:62
  wire              _GEN_584 = io_dmem_nack_0_bits_uop_ldq_idx == 4'hB;	// lsu.scala:305:44, :1293:62
  wire              _GEN_585 = io_dmem_nack_0_bits_uop_ldq_idx == 4'hC;	// lsu.scala:305:44, :1293:62
  wire              _GEN_586 = io_dmem_nack_0_bits_uop_ldq_idx == 4'hD;	// lsu.scala:305:44, :1293:62
  wire              _GEN_587 = io_dmem_nack_0_bits_uop_ldq_idx == 4'hE;	// lsu.scala:305:44, :1293:62
  assign nacking_loads_0 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_573;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_1 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_574;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_2 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_575;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_3 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_576;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_4 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_577;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_5 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_578;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_6 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_579;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_7 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_580;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_8 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_581;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_9 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_582;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_10 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_583;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_11 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_584;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_12 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_585;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_13 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_586;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_14 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_587;	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  assign nacking_loads_15 =
    io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella
    & io_dmem_nack_0_bits_uop_uses_ldq & (&io_dmem_nack_0_bits_uop_ldq_idx);	// lsu.scala:1284:5, :1287:7, :1291:7, :1293:62
  wire              _GEN_588 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq;	// lsu.scala:1308:7
  wire              send_iresp = _GEN_177[io_dmem_resp_0_bits_uop_ldq_idx] == 2'h0;	// lsu.scala:465:79, :1311:58
  wire              send_fresp = _GEN_177[io_dmem_resp_0_bits_uop_ldq_idx] == 2'h1;	// lsu.scala:465:79, :1311:58, :1312:58
  wire              _GEN_589 =
    io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_is_amo;	// lsu.scala:1328:7, :1331:48
  wire              dmem_resp_fired_0 =
    io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq | _GEN_589);	// lsu.scala:1306:5, :1308:7, :1322:28, :1328:7, :1331:48
  wire              _GEN_590 = dmem_resp_fired_0 & wb_forward_valid_0;	// lsu.scala:1064:36, :1306:5, :1308:7, :1343:30
  wire              _GEN_591 = ~dmem_resp_fired_0 & wb_forward_valid_0;	// lsu.scala:1064:36, :1306:5, :1308:7, :1347:{18,38}
  wire [11:0]       _GEN_592 = _GEN_102[wb_forward_ldq_idx_0];	// lsu.scala:264:49, :1065:36, util.scala:118:51
  wire [5:0]        _GEN_593 = _GEN_140[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire [6:0]        _GEN_594 = _GEN_145[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire [1:0]        _GEN_595 = _GEN_104[wb_forward_ldq_idx_0];	// lsu.scala:264:49, :1065:36, util.scala:118:51
  wire              _GEN_596 = _GEN_160[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire              _GEN_597 = _GEN_163[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire              _GEN_598 = _GEN_166[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire [1:0]        _GEN_599 = _GEN_177[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, util.scala:118:51
  wire              live = (io_core_brupdate_b1_mispredict_mask & _GEN_592) == 12'h0;	// util.scala:118:{51,59}
  wire              _GEN_600 = _GEN_91[wb_forward_stq_idx_0];	// AMOALU.scala:10:17, lsu.scala:224:42, :1067:36
  wire [63:0]       _GEN_601 = _GEN_92[wb_forward_stq_idx_0];	// AMOALU.scala:10:17, lsu.scala:224:42, :1067:36
  wire [3:0][63:0]  _GEN_602 =
    {{_GEN_601},
     {{2{_GEN_601[31:0]}}},
     {{2{{2{_GEN_601[15:0]}}}}},
     {{2{{2{{2{_GEN_601[7:0]}}}}}}}};	// AMOALU.scala:10:17, :26:{13,19,66}, Cat.scala:30:58
  wire [63:0]       _GEN_603 = _GEN_602[_GEN_55[wb_forward_stq_idx_0]];	// AMOALU.scala:10:17, :26:{13,19}, lsu.scala:224:42, :1067:36
  wire              _GEN_604 = _GEN_590 | ~_GEN_591;	// lsu.scala:1306:5, :1343:30, :1344:5, :1347:38, :1348:5
  wire              _io_core_exe_0_iresp_valid_output =
    _GEN_604
      ? io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq ? send_iresp : _GEN_589)
      : _GEN_599 == 2'h0 & _GEN_600 & live;	// AMOALU.scala:10:17, lsu.scala:1275:32, :1306:5, :1308:7, :1311:58, :1316:40, :1328:7, :1331:48, :1344:5, :1348:5, :1362:{60,86}, util.scala:118:{51,59}
  wire              _io_core_exe_0_fresp_valid_output =
    _GEN_604 ? _GEN_588 & send_fresp : _GEN_599 == 2'h1 & _GEN_600 & live;	// AMOALU.scala:10:17, lsu.scala:1276:32, :1306:5, :1308:7, :1312:58, :1318:40, :1344:5, :1348:5, :1363:{60,86}, util.scala:118:{51,59}
  wire [31:0]       io_core_exe_0_iresp_bits_data_lo =
    wb_forward_ld_addr_0[2] ? _GEN_603[63:32] : _GEN_603[31:0];	// AMOALU.scala:26:13, :39:{24,29,37,55}, lsu.scala:1066:36
  wire              _ldq_bits_debug_wb_data_T_1 = _GEN_595 == 2'h2;	// AMOALU.scala:42:26, util.scala:118:51, :351:72
  wire [15:0]       io_core_exe_0_iresp_bits_data_lo_1 =
    wb_forward_ld_addr_0[1]
      ? io_core_exe_0_iresp_bits_data_lo[31:16]
      : io_core_exe_0_iresp_bits_data_lo[15:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  wire              _ldq_bits_debug_wb_data_T_9 = _GEN_595 == 2'h1;	// AMOALU.scala:42:26, lsu.scala:1312:58, util.scala:118:51
  wire [7:0]        io_core_exe_0_iresp_bits_data_lo_2 =
    wb_forward_ld_addr_0[0]
      ? io_core_exe_0_iresp_bits_data_lo_1[15:8]
      : io_core_exe_0_iresp_bits_data_lo_1[7:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  wire              _ldq_bits_debug_wb_data_T_17 = _GEN_595 == 2'h0;	// AMOALU.scala:42:26, util.scala:118:51
  wire [31:0]       io_core_exe_0_fresp_bits_data_lo =
    wb_forward_ld_addr_0[2] ? _GEN_603[63:32] : _GEN_603[31:0];	// AMOALU.scala:26:13, :39:{24,29,37,55}, lsu.scala:1066:36
  wire [15:0]       io_core_exe_0_fresp_bits_data_lo_1 =
    wb_forward_ld_addr_0[1]
      ? io_core_exe_0_fresp_bits_data_lo[31:16]
      : io_core_exe_0_fresp_bits_data_lo[15:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  wire [7:0]        io_core_exe_0_fresp_bits_data_lo_2 =
    wb_forward_ld_addr_0[0]
      ? io_core_exe_0_fresp_bits_data_lo_1[15:8]
      : io_core_exe_0_fresp_bits_data_lo_1[7:0];	// AMOALU.scala:39:{24,29,37,55}, lsu.scala:1066:36
  reg               io_core_ld_miss_REG;	// lsu.scala:1380:37
  reg               spec_ld_succeed_REG;	// lsu.scala:1382:13
  reg  [3:0]        spec_ld_succeed_REG_1;	// lsu.scala:1384:56
  wire [11:0]       _GEN_605 =
    io_core_brupdate_b1_mispredict_mask & stq_0_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_606 =
    io_core_brupdate_b1_mispredict_mask & stq_1_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_607 =
    io_core_brupdate_b1_mispredict_mask & stq_2_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_608 =
    io_core_brupdate_b1_mispredict_mask & stq_3_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_609 =
    io_core_brupdate_b1_mispredict_mask & stq_4_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_610 =
    io_core_brupdate_b1_mispredict_mask & stq_5_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_611 =
    io_core_brupdate_b1_mispredict_mask & stq_6_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_612 =
    io_core_brupdate_b1_mispredict_mask & stq_7_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_613 =
    io_core_brupdate_b1_mispredict_mask & stq_8_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_614 =
    io_core_brupdate_b1_mispredict_mask & stq_9_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_615 =
    io_core_brupdate_b1_mispredict_mask & stq_10_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_616 =
    io_core_brupdate_b1_mispredict_mask & stq_11_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_617 =
    io_core_brupdate_b1_mispredict_mask & stq_12_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_618 =
    io_core_brupdate_b1_mispredict_mask & stq_13_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_619 =
    io_core_brupdate_b1_mispredict_mask & stq_14_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire [11:0]       _GEN_620 =
    io_core_brupdate_b1_mispredict_mask & stq_15_bits_uop_br_mask;	// lsu.scala:211:16, util.scala:118:51
  wire              commit_store =
    io_core_commit_valids_0 & io_core_commit_uops_0_uses_stq;	// lsu.scala:1451:49
  wire              commit_load =
    io_core_commit_valids_0 & io_core_commit_uops_0_uses_ldq;	// lsu.scala:1452:49
  wire [3:0]        idx = commit_store ? stq_commit_head : ldq_head;	// lsu.scala:215:29, :219:29, :1451:49, :1453:18
  wire [3:0]        _GEN_621 = stq_commit_head + 4'h1;	// lsu.scala:219:29, :305:44, util.scala:203:14
  wire [3:0]        _GEN_622 = commit_store ? _GEN_621 : stq_commit_head;	// lsu.scala:219:29, :1451:49, :1482:31, util.scala:203:14
  wire [3:0]        _GEN_623 = ldq_head + 4'h1;	// lsu.scala:215:29, :305:44, util.scala:203:14
  wire [3:0]        _GEN_624 = commit_load ? _GEN_623 : ldq_head;	// lsu.scala:215:29, :1452:49, :1486:31, util.scala:203:14
  wire              commit_store_1 =
    io_core_commit_valids_1 & io_core_commit_uops_1_uses_stq;	// lsu.scala:1451:49
  wire              commit_load_1 =
    io_core_commit_valids_1 & io_core_commit_uops_1_uses_ldq;	// lsu.scala:1452:49
  wire [3:0]        idx_1 = commit_store_1 ? _GEN_622 : _GEN_624;	// lsu.scala:1451:49, :1453:18, :1482:31, :1486:31
  `ifndef SYNTHESIS	// lsu.scala:224:10
    always @(posedge clock) begin	// lsu.scala:224:10
      automatic logic        _GEN_625 = ~dis_ld_val & dis_st_val;	// lsu.scala:301:85, :302:85, :304:5, :321:5
      automatic logic        _GEN_626 = ~dis_ld_val_1 & dis_st_val_1;	// lsu.scala:301:85, :302:85, :304:5, :321:5
      automatic logic        _GEN_627 =
        ~can_fire_load_incoming_0 & ~will_fire_load_retry_0 & ~will_fire_store_commit_0;	// lsu.scala:441:63, :535:65, :584:6, :766:39, :773:43, :780:45
      automatic logic        _GEN_628 = _GEN_627 & ~will_fire_load_wakeup_0;	// lsu.scala:535:65, :780:45, :794:44
      automatic logic        _GEN_629 =
        io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella;	// lsu.scala:1287:7
      automatic logic        _GEN_630 = ~io_dmem_resp_0_bits_is_hella | reset;	// lsu.scala:1309:{15,16}
      automatic logic        _GEN_631 = ~commit_store & commit_load;	// lsu.scala:1451:49, :1452:49, :1455:5, :1457:31
      automatic logic [15:0] _GEN_632;	// lsu.scala:1458:14
      automatic logic        _GEN_633 = ~commit_store_1 & commit_load_1;	// lsu.scala:1451:49, :1452:49, :1455:5, :1457:31
      _GEN_632 =
        {{ldq_15_bits_forward_std_val},
         {ldq_14_bits_forward_std_val},
         {ldq_13_bits_forward_std_val},
         {ldq_12_bits_forward_std_val},
         {ldq_11_bits_forward_std_val},
         {ldq_10_bits_forward_std_val},
         {ldq_9_bits_forward_std_val},
         {ldq_8_bits_forward_std_val},
         {ldq_7_bits_forward_std_val},
         {ldq_6_bits_forward_std_val},
         {ldq_5_bits_forward_std_val},
         {ldq_4_bits_forward_std_val},
         {ldq_3_bits_forward_std_val},
         {ldq_2_bits_forward_std_val},
         {ldq_1_bits_forward_std_val},
         {ldq_0_bits_forward_std_val}};	// lsu.scala:210:16, :1458:14
      if (~(io_core_brupdate_b2_mispredict | _GEN_3 | stq_head == stq_execute_head
            | stq_tail == stq_execute_head | reset)) begin	// lsu.scala:217:29, :218:29, :220:29, :224:{10,42}, :226:20, :227:20
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:224:10
          $error("Assertion failed: stq_execute_head got off track.\n    at lsu.scala:224 assert (io.core.brupdate.b2.mispredict ||\n");	// lsu.scala:224:10
        if (`STOP_COND_)	// lsu.scala:224:10
          $fatal;	// lsu.scala:224:10
      end
      if (dis_ld_val & ~(ldq_tail == io_core_dis_uops_0_bits_ldq_idx | reset)) begin	// lsu.scala:216:29, :301:85, :317:{14,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:317:14
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:317 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");	// lsu.scala:317:14
        if (`STOP_COND_)	// lsu.scala:317:14
          $fatal;	// lsu.scala:317:14
      end
      if (dis_ld_val & ~(~_GEN_97[ldq_tail] | reset)) begin	// lsu.scala:216:29, :301:85, :305:44, :318:{14,15}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:318:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:318 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");	// lsu.scala:318:14
        if (`STOP_COND_)	// lsu.scala:318:14
          $fatal;	// lsu.scala:318:14
      end
      if (_GEN_625 & ~(stq_tail == io_core_dis_uops_0_bits_stq_idx | reset)) begin	// lsu.scala:218:29, :321:5, :329:{14,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:329:14
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:329 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");	// lsu.scala:329:14
        if (`STOP_COND_)	// lsu.scala:329:14
          $fatal;	// lsu.scala:329:14
      end
      if (_GEN_625 & ~(~_GEN_2[stq_tail] | reset)) begin	// lsu.scala:218:29, :224:42, :321:5, :322:39, :330:{14,15}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:330:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:330 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");	// lsu.scala:330:14
        if (`STOP_COND_)	// lsu.scala:330:14
          $fatal;	// lsu.scala:330:14
      end
      if (~(~(dis_ld_val & dis_st_val) | reset)) begin	// lsu.scala:301:85, :302:85, :341:{11,12,25}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:341:11
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:341 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");	// lsu.scala:341:11
        if (`STOP_COND_)	// lsu.scala:341:11
          $fatal;	// lsu.scala:341:11
      end
      if (dis_ld_val_1 & ~(_GEN_98 == io_core_dis_uops_1_bits_ldq_idx | reset)) begin	// lsu.scala:301:85, :317:{14,26}, :333:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:317:14
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:317 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");	// lsu.scala:317:14
        if (`STOP_COND_)	// lsu.scala:317:14
          $fatal;	// lsu.scala:317:14
      end
      if (dis_ld_val_1 & ~(~_GEN_97[_GEN_98] | reset)) begin	// lsu.scala:301:85, :305:44, :318:{14,15}, :333:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:318:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:318 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");	// lsu.scala:318:14
        if (`STOP_COND_)	// lsu.scala:318:14
          $fatal;	// lsu.scala:318:14
      end
      if (_GEN_626 & ~(_GEN_99 == io_core_dis_uops_1_bits_stq_idx | reset)) begin	// lsu.scala:321:5, :329:{14,26}, :338:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:329:14
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:329 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");	// lsu.scala:329:14
        if (`STOP_COND_)	// lsu.scala:329:14
          $fatal;	// lsu.scala:329:14
      end
      if (_GEN_626 & ~(~_GEN_2[_GEN_99] | reset)) begin	// lsu.scala:224:42, :321:5, :322:39, :330:{14,15}, :338:21
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:330:14
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:330 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");	// lsu.scala:330:14
        if (`STOP_COND_)	// lsu.scala:330:14
          $fatal;	// lsu.scala:330:14
      end
      if (~(~(dis_ld_val_1 & dis_st_val_1) | reset)) begin	// lsu.scala:301:85, :302:85, :341:{11,12,25}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:341:11
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:341 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");	// lsu.scala:341:11
        if (`STOP_COND_)	// lsu.scala:341:11
          $fatal;	// lsu.scala:341:11
      end
      if (~(~(io_core_exe_0_req_valid
              & ~(_GEN_207 | will_fire_std_incoming_0 | will_fire_sfence_0))
            | reset)) begin	// lsu.scala:536:61, :567:{11,12,31,34,93,151}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:567:11
          $error("Assertion failed\n    at lsu.scala:567 assert(!(exe_req(w).valid && !(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) || will_fire_std_incoming(w) || will_fire_sfence(w))))\n");	// lsu.scala:567:11
        if (`STOP_COND_)	// lsu.scala:567:11
          $fatal;	// lsu.scala:567:11
      end
      if (~(~((|hella_state) & hella_req_cmd == 5'h14) | reset)) begin	// Mux.scala:47:69, lsu.scala:242:38, :243:34, :593:{9,10,24,36,53}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:593:9
          $error("Assertion failed: SFENCE through hella interface not supported\n    at lsu.scala:593 assert(!(hella_state =/= h_ready && hella_req.cmd === rocket.M_SFENCE),\n");	// lsu.scala:593:9
        if (`STOP_COND_)	// lsu.scala:593:9
          $fatal;	// lsu.scala:593:9
      end
      if (~(~(~_will_fire_store_commit_0_T_2 & exe_tlb_uop_0_is_fence) | reset)) begin	// lsu.scala:538:31, :576:25, :597:24, :682:{12,13,36}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:682:12
          $error("Assertion failed: Fence is pretending to talk to the TLB\n    at lsu.scala:682 assert (!(dtlb.io.req(w).valid && exe_tlb_uop(w).is_fence), \"Fence is pretending to talk to the TLB\")\n");	// lsu.scala:682:12
        if (`STOP_COND_)	// lsu.scala:682:12
          $fatal;	// lsu.scala:682:12
      end
      if (~(~((can_fire_load_incoming_0 | will_fire_sta_incoming_0
               | will_fire_stad_incoming_0) & io_core_exe_0_req_bits_mxcpt_valid
              & ~_will_fire_store_commit_0_T_2
              & ~(exe_tlb_uop_0_ctrl_is_load | exe_tlb_uop_0_ctrl_is_sta)) | reset)) begin	// lsu.scala:441:63, :534:63, :536:61, :538:31, :576:25, :597:24, :683:{12,13,72}, :684:59, :685:{5,35}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:683:12
          $error("Assertion failed: A uop that's not a load or store-address is throwing a memory exception.\n    at lsu.scala:683 assert (!((will_fire_load_incoming(w) || will_fire_sta_incoming(w) || will_fire_stad_incoming(w)) &&\n");	// lsu.scala:683:12
        if (`STOP_COND_)	// lsu.scala:683:12
          $fatal;	// lsu.scala:683:12
      end
      if (~(exe_tlb_paddr_0 == _dtlb_io_resp_0_paddr | io_core_exe_0_req_bits_sfence_valid
            | reset)) begin	// Cat.scala:30:58, lsu.scala:249:20, :714:{12,30}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:714:12
          $error("Assertion failed: [lsu] paddrs should match.\n    at lsu.scala:714 assert (exe_tlb_paddr(w) === dtlb.io.resp(w).paddr || exe_req(w).bits.sfence.valid, \"[lsu] paddrs should match.\")\n");	// lsu.scala:714:12
        if (`STOP_COND_)	// lsu.scala:714:12
          $fatal;	// lsu.scala:714:12
      end
      if (mem_xcpt_valids_0 & ~(REG | reset)) begin	// lsu.scala:667:32, :718:{13,21}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:718:13
          $error("Assertion failed\n    at lsu.scala:718 assert(RegNext(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) ||\n");	// lsu.scala:718:13
        if (`STOP_COND_)	// lsu.scala:718:13
          $fatal;	// lsu.scala:718:13
      end
      if (mem_xcpt_valids_0
          & ~(mem_xcpt_uops_0_uses_ldq ^ mem_xcpt_uops_0_uses_stq | reset)) begin	// lsu.scala:667:32, :671:32, :721:{13,40}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:721:13
          $error("Assertion failed\n    at lsu.scala:721 assert(mem_xcpt_uops(w).uses_ldq ^ mem_xcpt_uops(w).uses_stq)\n");	// lsu.scala:721:13
        if (`STOP_COND_)	// lsu.scala:721:13
          $fatal;	// lsu.scala:721:13
      end
      if (can_fire_load_incoming_0
          & ~(~_GEN_106[io_core_exe_0_req_bits_uop_ldq_idx] | reset)) begin	// lsu.scala:264:49, :441:63, :772:{13,14}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:772:13
          $error("Assertion failed\n    at lsu.scala:772 assert(!ldq_incoming_e(w).bits.executed)\n");	// lsu.scala:772:13
        if (`STOP_COND_)	// lsu.scala:772:13
          $fatal;	// lsu.scala:772:13
      end
      if (~can_fire_load_incoming_0 & will_fire_load_retry_0
          & ~(~_GEN_106[ldq_retry_idx] | reset)) begin	// lsu.scala:264:49, :415:30, :441:63, :465:79, :535:65, :766:39, :779:{13,14}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:779:13
          $error("Assertion failed\n    at lsu.scala:779 assert(!ldq_retry_e.bits.executed)\n");	// lsu.scala:779:13
        if (`STOP_COND_)	// lsu.scala:779:13
          $fatal;	// lsu.scala:779:13
      end
      if (_GEN_627 & will_fire_load_wakeup_0 & ~(~_GEN_205 & ~_GEN_203 | reset)) begin	// lsu.scala:502:88, :505:31, :506:31, :535:65, :780:45, :801:{13,42}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:801:13
          $error("Assertion failed\n    at lsu.scala:801 assert(!ldq_wakeup_e.bits.executed && !ldq_wakeup_e.bits.addr_is_virtual)\n");	// lsu.scala:801:13
        if (`STOP_COND_)	// lsu.scala:801:13
          $fatal;	// lsu.scala:801:13
      end
      if (_GEN_628 & will_fire_hella_incoming_0 & ~(_GEN_1 | reset)) begin	// lsu.scala:535:65, :794:44, :803:{13,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:803:13
          $error("Assertion failed\n    at lsu.scala:803 assert(hella_state === h_s1)\n");	// lsu.scala:803:13
        if (`STOP_COND_)	// lsu.scala:803:13
          $fatal;	// lsu.scala:803:13
      end
      if (_GEN_628 & ~will_fire_hella_incoming_0 & will_fire_hella_wakeup_0
          & ~(_GEN_0 | reset)) begin	// lsu.scala:535:65, :794:44, :802:47, :820:{13,26}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:820:13
          $error("Assertion failed\n    at lsu.scala:820 assert(hella_state === h_replay)\n");	// lsu.scala:820:13
        if (`STOP_COND_)	// lsu.scala:820:13
          $fatal;	// lsu.scala:820:13
      end
      if (_GEN_272
          & ~(~(can_fire_load_incoming_0 & _GEN_105[io_core_exe_0_req_bits_uop_ldq_idx])
              | reset)) begin	// lsu.scala:220:29, :264:49, :441:63, :766:39, :773:43, :780:45, :844:{13,14,43}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:844:13
          $error("Assertion failed: [lsu] Incoming load is overwriting a valid address\n    at lsu.scala:844 assert(!(will_fire_load_incoming(w) && ldq_incoming_e(w).bits.addr.valid),\n");	// lsu.scala:844:13
        if (`STOP_COND_)	// lsu.scala:844:13
          $fatal;	// lsu.scala:844:13
      end
      if (_GEN_278
          & ~(~(will_fire_sta_incoming_0 & _GEN_87[io_core_exe_0_req_bits_uop_stq_idx])
              | reset)) begin	// lsu.scala:224:42, :264:49, :536:61, :848:67, :858:{13,14,42}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:858:13
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid address\n    at lsu.scala:858 assert(!(will_fire_sta_incoming(w) && stq_incoming_e(w).bits.addr.valid),\n");	// lsu.scala:858:13
        if (`STOP_COND_)	// lsu.scala:858:13
          $fatal;	// lsu.scala:858:13
      end
      if (_GEN_279 & ~(~_GEN_91[sidx] | reset)) begin	// lsu.scala:224:42, :868:67, :870:21, :873:33, :877:{13,14}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:877:13
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid data entry\n    at lsu.scala:877 assert(!(stq(sidx).bits.data.valid),\n");	// lsu.scala:877:13
        if (`STOP_COND_)	// lsu.scala:877:13
          $fatal;	// lsu.scala:877:13
      end
      if (_GEN_570 & ~(_GEN_571 | _GEN_572 | reset)) begin	// lsu.scala:1287:7, :1288:{15,28,54}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1288:15
          $error("Assertion failed\n    at lsu.scala:1288 assert(hella_state === h_wait || hella_state === h_dead)\n");	// lsu.scala:1288:15
        if (`STOP_COND_)	// lsu.scala:1288:15
          $fatal;	// lsu.scala:1288:15
      end
      if (_GEN_629 & io_dmem_nack_0_bits_uop_uses_ldq
          & ~(_GEN_106[io_dmem_nack_0_bits_uop_ldq_idx] | reset)) begin	// lsu.scala:264:49, :1287:7, :1292:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1292:15
          $error("Assertion failed\n    at lsu.scala:1292 assert(ldq(io.dmem.nack(w).bits.uop.ldq_idx).bits.executed)\n");	// lsu.scala:1292:15
        if (`STOP_COND_)	// lsu.scala:1292:15
          $fatal;	// lsu.scala:1292:15
      end
      if (_GEN_629 & ~io_dmem_nack_0_bits_uop_uses_ldq
          & ~(io_dmem_nack_0_bits_uop_uses_stq | reset)) begin	// lsu.scala:1287:7, :1291:7, :1298:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1298:15
          $error("Assertion failed\n    at lsu.scala:1298 assert(io.dmem.nack(w).bits.uop.uses_stq)\n");	// lsu.scala:1298:15
        if (`STOP_COND_)	// lsu.scala:1298:15
          $fatal;	// lsu.scala:1298:15
      end
      if (_GEN_588 & ~_GEN_630) begin	// lsu.scala:1308:7, :1309:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1309:15
          $error("Assertion failed\n    at lsu.scala:1309 assert(!io.dmem.resp(w).bits.is_hella)\n");	// lsu.scala:1309:15
        if (`STOP_COND_)	// lsu.scala:1309:15
          $fatal;	// lsu.scala:1309:15
      end
      if (_GEN_588 & ~(send_iresp ^ send_fresp | reset)) begin	// lsu.scala:1308:7, :1311:58, :1312:58, :1321:{15,27}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1321:15
          $error("Assertion failed\n    at lsu.scala:1321 assert(send_iresp ^ send_fresp)\n");	// lsu.scala:1321:15
        if (`STOP_COND_)	// lsu.scala:1321:15
          $fatal;	// lsu.scala:1321:15
      end
      if (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
          & io_dmem_resp_0_bits_uop_uses_stq & ~_GEN_630) begin	// lsu.scala:1308:7, :1309:15, :1329:15
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1329:15
          $error("Assertion failed\n    at lsu.scala:1329 assert(!io.dmem.resp(w).bits.is_hella)\n");	// lsu.scala:1329:15
        if (`STOP_COND_)	// lsu.scala:1329:15
          $fatal;	// lsu.scala:1329:15
      end
      if (~(~((|_GEN_605) & stq_0_valid & stq_0_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_606) & stq_1_valid & stq_1_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_607) & stq_2_valid & stq_2_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_608) & stq_3_valid & stq_3_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_609) & stq_4_valid & stq_4_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_610) & stq_5_valid & stq_5_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_611) & stq_6_valid & stq_6_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_612) & stq_7_valid & stq_7_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_613) & stq_8_valid & stq_8_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_614) & stq_9_valid & stq_9_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_615) & stq_10_valid & stq_10_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_616) & stq_11_valid & stq_11_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_617) & stq_12_valid & stq_12_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_618) & stq_13_valid & stq_13_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_619) & stq_14_valid & stq_14_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (~(~((|_GEN_620) & stq_15_valid & stq_15_bits_committed) | reset)) begin	// lsu.scala:211:16, :1416:{12,13,83}, util.scala:118:{51,59}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1416:12
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1416 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");	// lsu.scala:1416:12
        if (`STOP_COND_)	// lsu.scala:1416:12
          $fatal;	// lsu.scala:1416:12
      end
      if (_GEN_631 & ~(_GEN_97[idx] | reset)) begin	// lsu.scala:305:44, :1453:18, :1457:31, :1458:14
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1458:14
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1458 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");	// lsu.scala:1458:14
        if (`STOP_COND_)	// lsu.scala:1458:14
          $fatal;	// lsu.scala:1458:14
      end
      if (_GEN_631 & ~((_GEN_106[idx] | _GEN_632[idx]) & _GEN_206[idx] | reset)) begin	// lsu.scala:264:49, :502:88, :1453:18, :1457:31, :1458:14, :1459:{14,39,73}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1459:14
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1459 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");	// lsu.scala:1459:14
        if (`STOP_COND_)	// lsu.scala:1459:14
          $fatal;	// lsu.scala:1459:14
      end
      if (_GEN_633 & ~(_GEN_97[idx_1] | reset)) begin	// lsu.scala:305:44, :1453:18, :1457:31, :1458:14
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1458:14
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1458 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");	// lsu.scala:1458:14
        if (`STOP_COND_)	// lsu.scala:1458:14
          $fatal;	// lsu.scala:1458:14
      end
      if (_GEN_633
          & ~((_GEN_106[idx_1] | _GEN_632[idx_1]) & _GEN_206[idx_1] | reset)) begin	// lsu.scala:264:49, :502:88, :1453:18, :1457:31, :1458:14, :1459:{14,39,73}
        if (`ASSERT_VERBOSE_COND_)	// lsu.scala:1459:14
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1459 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");	// lsu.scala:1459:14
        if (`STOP_COND_)	// lsu.scala:1459:14
          $fatal;	// lsu.scala:1459:14
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire              _GEN_634 = _GEN_58[stq_head];	// lsu.scala:217:29, :224:42, :1494:29
  wire [15:0]       _GEN_635 =
    {{stq_15_bits_succeeded},
     {stq_14_bits_succeeded},
     {stq_13_bits_succeeded},
     {stq_12_bits_succeeded},
     {stq_11_bits_succeeded},
     {stq_10_bits_succeeded},
     {stq_9_bits_succeeded},
     {stq_8_bits_succeeded},
     {stq_7_bits_succeeded},
     {stq_6_bits_succeeded},
     {stq_5_bits_succeeded},
     {stq_4_bits_succeeded},
     {stq_3_bits_succeeded},
     {stq_2_bits_succeeded},
     {stq_1_bits_succeeded},
     {stq_0_bits_succeeded}};	// lsu.scala:211:16, :1494:29
  wire              _GEN_636 = _GEN_2[stq_head] & _GEN_94[stq_head];	// lsu.scala:217:29, :224:42, :1494:29
  wire              _GEN_637 = _GEN_634 & ~io_dmem_ordered;	// lsu.scala:1494:29, :1496:{43,46}
  assign store_needs_order = _GEN_636 & _GEN_637;	// lsu.scala:1494:29, :1495:3, :1496:{43,64}
  wire              clear_store =
    _GEN_636 & (_GEN_634 ? io_dmem_ordered : _GEN_635[stq_head]);	// lsu.scala:217:29, :1494:29, :1495:3, :1500:{17,23}
  wire              _GEN_638 = hella_state == 3'h3;	// lsu.scala:242:38, :1548:19, :1550:28
  wire              _GEN_639 = ~(|hella_state) | _GEN_1;	// lsu.scala:242:38, :593:24, :803:26, :1524:27, :1527:{21,34}, :1533:38, :1550:43
  wire              _GEN_640 = hella_state == 3'h2;	// lsu.scala:242:38, :1546:19, :1553:28
  wire              _GEN_641 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_is_hella;	// lsu.scala:1562:35
  assign _GEN = ~(~(|hella_state) | _GEN_1 | _GEN_638 | _GEN_640 | _GEN_571);	// lsu.scala:242:38, :593:24, :803:26, :1288:28, :1527:{21,34}, :1533:38, :1550:{28,43}, :1553:{28,38}, :1560:40, :1576:42
  always @(posedge clock) begin
    automatic logic [15:0] _ldq_15_bits_st_dep_mask_T;	// lsu.scala:260:71
    automatic logic [15:0] _GEN_642;	// lsu.scala:260:33
    automatic logic [15:0] next_live_store_mask;	// lsu.scala:260:33
    automatic logic        _GEN_643;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_644;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_645;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_646;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_647;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_648;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_649;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_650;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_651;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_652;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_653;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_654;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_655;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_656;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_657;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_658;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_659;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_660;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_661;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_662;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_663;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_664;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_665;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_666;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_667;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_668;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_669;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_670;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_671;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_672;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_673;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_674;	// lsu.scala:211:16, :321:5, :322:39
    automatic logic        _GEN_675;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_676;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_677;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_678;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_679;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_680;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_681;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_682;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_683;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_684;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_685;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_686;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_687;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_688;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_689;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic        _GEN_690;	// lsu.scala:211:16, :304:5, :321:5
    automatic logic [15:0] _GEN_691;	// lsu.scala:336:31
    automatic logic        _GEN_692 = _GEN_98 == 4'h0;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_693;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_694;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_695 = _GEN_98 == 4'h1;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_696;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_697;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_698 = _GEN_98 == 4'h2;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_699;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_700;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_701 = _GEN_98 == 4'h3;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_702;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_703;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_704 = _GEN_98 == 4'h4;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_705;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_706;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_707 = _GEN_98 == 4'h5;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_708;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_709;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_710 = _GEN_98 == 4'h6;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_711;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_712;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_713 = _GEN_98 == 4'h7;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_714;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_715;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_716 = _GEN_98 == 4'h8;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_717;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_718;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_719 = _GEN_98 == 4'h9;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_720;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_721;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_722 = _GEN_98 == 4'hA;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_723;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_724;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_725 = _GEN_98 == 4'hB;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_726;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_727;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_728 = _GEN_98 == 4'hC;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_729;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_730;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_731 = _GEN_98 == 4'hD;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_732;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_733;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_734 = _GEN_98 == 4'hE;	// lsu.scala:305:44, :333:21
    automatic logic        _GEN_735;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_736;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_737;	// lsu.scala:210:16, :304:5, :305:44
    automatic logic        _GEN_738;	// lsu.scala:304:5, :305:44
    automatic logic        _GEN_739;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_740;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_741;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_742;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_743;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_744;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_745;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_746;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_747;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_748;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_749;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_750;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_751;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_752;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_753;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_754;	// lsu.scala:304:5, :306:44
    automatic logic        _GEN_755;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_756;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_757;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_758;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_759;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_760;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_761;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_762;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_763;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_764;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_765;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_766;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_767;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_768;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_769;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_770;	// lsu.scala:210:16, :304:5, :306:44
    automatic logic        _GEN_771;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_772;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_773;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_774;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_775;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_776;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_777;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_778;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_779;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_780;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_781;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_782;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_783;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_784;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_785;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_786;	// lsu.scala:304:5, :313:44
    automatic logic        _GEN_787;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_788;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_789;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_790;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_791;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_792;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_793;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_794;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_795;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_796;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_797;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_798;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_799;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_800;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_801;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_802;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_803;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_804;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_805;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_806;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_807;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_808;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_809;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_810;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_811;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_812;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_813;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_814;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_815;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_816;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_817;	// lsu.scala:304:5, :321:5, :322:39
    automatic logic        _GEN_818;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_819;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_820;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_821;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_822;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_823;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_824;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_825;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_826;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_827;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_828;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_829;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_830;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_831;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_832;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_833;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_834;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_835;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_836;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_837;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_838;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_839;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_840;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_841;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_842;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_843;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_844;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_845;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_846;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_847;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_848;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_849;	// lsu.scala:304:5, :321:5
    automatic logic        _GEN_850;	// lsu.scala:304:5, :321:5
    automatic logic        ldq_retry_idx_block;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_2;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_1;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_5;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_2;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_8;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_3;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_11;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_4;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_14;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_5;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_17;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_6;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_20;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_7;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_23;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_8;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_26;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_9;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_29;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_10;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_32;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_11;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_35;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_12;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_38;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_13;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_41;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_14;	// lsu.scala:417:36
    automatic logic        _ldq_retry_idx_T_44;	// lsu.scala:418:39
    automatic logic        ldq_retry_idx_block_15;	// lsu.scala:417:36
    automatic logic        _temp_bits_T;	// util.scala:351:72
    automatic logic        _temp_bits_T_2;	// util.scala:351:72
    automatic logic        _temp_bits_T_4;	// util.scala:351:72
    automatic logic        _temp_bits_T_6;	// util.scala:351:72
    automatic logic        _temp_bits_T_8;	// util.scala:351:72
    automatic logic        _temp_bits_T_10;	// util.scala:351:72
    automatic logic        _temp_bits_T_12;	// util.scala:351:72
    automatic logic        _temp_bits_T_16;	// util.scala:351:72
    automatic logic        _temp_bits_T_18;	// util.scala:351:72
    automatic logic        _temp_bits_T_20;	// util.scala:351:72
    automatic logic        _temp_bits_T_22;	// util.scala:351:72
    automatic logic        _temp_bits_T_24;	// util.scala:351:72
    automatic logic        _temp_bits_T_26;	// util.scala:351:72
    automatic logic        _temp_bits_T_28;	// util.scala:351:72
    automatic logic        _stq_retry_idx_T;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_1;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_2;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_3;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_4;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_5;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_6;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_7;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_8;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_9;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_10;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_11;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_12;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_13;	// lsu.scala:424:18
    automatic logic        _stq_retry_idx_T_14;	// lsu.scala:424:18
    automatic logic        _ldq_wakeup_idx_T_7;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_15;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_23;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_31;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_39;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_47;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_55;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_63;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_71;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_79;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_87;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_95;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_103;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_111;	// lsu.scala:433:71
    automatic logic        _ldq_wakeup_idx_T_119;	// lsu.scala:433:71
    automatic logic        ma_ld_0 =
      can_fire_load_incoming_0 & io_core_exe_0_req_bits_mxcpt_valid;	// lsu.scala:441:63, :659:56
    automatic logic        ma_st_0;	// lsu.scala:660:87
    automatic logic        pf_ld_0;	// lsu.scala:661:75
    automatic logic        pf_st_0;	// lsu.scala:662:75
    automatic logic        ae_ld_0;	// lsu.scala:663:75
    automatic logic        dmem_req_fire_0;	// lsu.scala:752:55
    automatic logic [3:0]  ldq_idx;	// lsu.scala:837:24
    automatic logic        _GEN_851;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_852;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_853;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_854;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_855;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_856;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_857;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_858;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_859;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_860;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_861;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_862;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_863;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_864;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_865;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_866;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_867;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_868;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_869;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_870;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_871;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_872;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_873;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_874;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_875;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_876;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_877;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_878;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_879;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_880;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_881;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _GEN_882;	// lsu.scala:304:5, :836:5, :838:45
    automatic logic        _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:842:71
    automatic logic [3:0]  stq_idx;	// lsu.scala:850:24
    automatic logic        _GEN_883;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_884;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_885;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_886;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_887;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_888;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_889;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_890;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_891;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_892;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_893;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_894;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_895;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_896;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_897;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_898;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_899;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_900;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_901;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_902;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_903;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_904;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_905;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_906;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_907;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_908;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_909;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_910;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_911;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_912;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_913;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_914;	// lsu.scala:304:5, :849:5, :853:36
    automatic logic        _GEN_915 = _GEN_279 & sidx == 4'h0;	// lsu.scala:304:5, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_916;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_917 = _GEN_279 & sidx == 4'h1;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_918;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_919 = _GEN_279 & sidx == 4'h2;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_920;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_921 = _GEN_279 & sidx == 4'h3;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_922;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_923 = _GEN_279 & sidx == 4'h4;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_924;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_925 = _GEN_279 & sidx == 4'h5;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_926;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_927 = _GEN_279 & sidx == 4'h6;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_928;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_929 = _GEN_279 & sidx == 4'h7;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_930;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_931 = _GEN_279 & sidx == 4'h8;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_932;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_933 = _GEN_279 & sidx == 4'h9;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_934;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_935 = _GEN_279 & sidx == 4'hA;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_936;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_937 = _GEN_279 & sidx == 4'hB;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_938;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_939 = _GEN_279 & sidx == 4'hC;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_940;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_941 = _GEN_279 & sidx == 4'hD;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_942;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_943 = _GEN_279 & sidx == 4'hE;	// lsu.scala:304:5, :305:44, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_944;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _GEN_945 = _GEN_279 & (&sidx);	// lsu.scala:304:5, :868:67, :869:5, :870:21, :873:33
    automatic logic        _GEN_946;	// lsu.scala:304:5, :869:5, :873:33
    automatic logic        _fired_std_incoming_T =
      (io_core_brupdate_b1_mispredict_mask & io_core_exe_0_req_bits_uop_br_mask) == 12'h0;	// util.scala:118:{51,59}
    automatic logic [11:0] _mem_stq_retry_e_out_valid_T =
      io_core_brupdate_b1_mispredict_mask & _GEN_197;	// lsu.scala:478:79, util.scala:118:51
    automatic logic [3:0]  l_forward_stq_idx;	// lsu.scala:1077:32
    automatic logic        _GEN_947;	// lsu.scala:1106:39
    automatic logic        _GEN_948;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_16;	// lsu.scala:1091:36, :1102:37
    automatic logic        _GEN_949 = lcam_ldq_idx_0 == 4'h1;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_950 = lcam_ldq_idx_0 == 4'h2;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_951 = lcam_ldq_idx_0 == 4'h3;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_952 = lcam_ldq_idx_0 == 4'h4;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_953 = lcam_ldq_idx_0 == 4'h5;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_954 = lcam_ldq_idx_0 == 4'h6;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_955 = lcam_ldq_idx_0 == 4'h7;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_956 = lcam_ldq_idx_0 == 4'h8;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_957 = lcam_ldq_idx_0 == 4'h9;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_958 = lcam_ldq_idx_0 == 4'hA;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_959 = lcam_ldq_idx_0 == 4'hB;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_960 = lcam_ldq_idx_0 == 4'hC;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_961 = lcam_ldq_idx_0 == 4'hD;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic        _GEN_962 = lcam_ldq_idx_0 == 4'hE;	// lsu.scala:305:44, :1036:26, :1130:48
    automatic logic [3:0]  l_forward_stq_idx_1;	// lsu.scala:1077:32
    automatic logic        _GEN_963;	// lsu.scala:1106:39
    automatic logic        _GEN_964;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_17;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_2;	// lsu.scala:1077:32
    automatic logic        _GEN_965;	// lsu.scala:1106:39
    automatic logic        _GEN_966;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_18;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_3;	// lsu.scala:1077:32
    automatic logic        _GEN_967;	// lsu.scala:1106:39
    automatic logic        _GEN_968;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_19;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_4;	// lsu.scala:1077:32
    automatic logic        _GEN_969;	// lsu.scala:1106:39
    automatic logic        _GEN_970;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_20;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_5;	// lsu.scala:1077:32
    automatic logic        _GEN_971;	// lsu.scala:1106:39
    automatic logic        _GEN_972;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_21;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_6;	// lsu.scala:1077:32
    automatic logic        _GEN_973;	// lsu.scala:1106:39
    automatic logic        _GEN_974;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_22;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_7;	// lsu.scala:1077:32
    automatic logic        _GEN_975;	// lsu.scala:1106:39
    automatic logic        _GEN_976;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_23;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_8;	// lsu.scala:1077:32
    automatic logic        _GEN_977;	// lsu.scala:1106:39
    automatic logic        _GEN_978;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_24;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_9;	// lsu.scala:1077:32
    automatic logic        _GEN_979;	// lsu.scala:1106:39
    automatic logic        _GEN_980;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_25;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_10;	// lsu.scala:1077:32
    automatic logic        _GEN_981;	// lsu.scala:1106:39
    automatic logic        _GEN_982;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_26;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_11;	// lsu.scala:1077:32
    automatic logic        _GEN_983;	// lsu.scala:1106:39
    automatic logic        _GEN_984;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_27;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_12;	// lsu.scala:1077:32
    automatic logic        _GEN_985;	// lsu.scala:1106:39
    automatic logic        _GEN_986;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_28;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_13;	// lsu.scala:1077:32
    automatic logic        _GEN_987;	// lsu.scala:1106:39
    automatic logic        _GEN_988;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_29;	// lsu.scala:1091:36, :1102:37
    automatic logic [3:0]  l_forward_stq_idx_14;	// lsu.scala:1077:32
    automatic logic        _GEN_989;	// lsu.scala:1106:39
    automatic logic        _GEN_990;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_30;	// lsu.scala:1091:36, :1102:37
    automatic logic        _GEN_991;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic [3:0]  l_forward_stq_idx_15;	// lsu.scala:1077:32
    automatic logic        _GEN_992;	// lsu.scala:1106:39
    automatic logic        _GEN_993;	// lsu.scala:1120:40
    automatic logic        _temp_bits_WIRE_1_31;	// lsu.scala:1091:36, :1102:37
    automatic logic        _GEN_994;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_995;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_996;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_997;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_998;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_999;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1000;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1001;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1002;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1003;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1004;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1005;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1006;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1007;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1008;	// lsu.scala:1091:36, :1102:37, :1116:37
    automatic logic        _GEN_1009 = _GEN_462 | _GEN_463;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1010;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1011;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1012;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1013;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1014;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1015;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1016;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1017;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1018;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1019;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1020;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1021;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1022;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1023;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1024;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1025;	// lsu.scala:1091:36, :1148:72, :1150:9
    automatic logic        _GEN_1026 = _GEN_469 | _GEN_470;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1027;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1028;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1029;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1030;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1031;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1032;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1033;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1034;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1035;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1036;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1037;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1038;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1039;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1040;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1041;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1042;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1043 = _GEN_476 | _GEN_477;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1044;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1045;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1046;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1047;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1048;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1049;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1050;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1051;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1052;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1053;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1054;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1055;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1056;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1057;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1058;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1059;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1060 = _GEN_483 | _GEN_484;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1061;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1062;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1063;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1064;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1065;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1066;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1067;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1068;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1069;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1070;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1071;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1072;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1073;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1074;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1075;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1076;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1077 = _GEN_490 | _GEN_491;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1078;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1079;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1080;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1081;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1082;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1083;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1084;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1085;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1086;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1087;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1088;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1089;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1090;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1091;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1092;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1093;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1094 = _GEN_497 | _GEN_498;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1095;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1096;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1097;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1098;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1099;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1100;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1101;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1102;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1103;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1104;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1105;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1106;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1107;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1108;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1109;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1110;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1111 = _GEN_504 | _GEN_505;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1112;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1113;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1114;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1115;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1116;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1117;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1118;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1119;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1120;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1121;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1122;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1123;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1124;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1125;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1126;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1127;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1128 = _GEN_511 | _GEN_512;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1129;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1130;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1131;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1132;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1133;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1134;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1135;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1136;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1137;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1138;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1139;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1140;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1141;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1142;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1143;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1144;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1145 = _GEN_518 | _GEN_519;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1146;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1147;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1148;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1149;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1150;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1151;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1152;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1153;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1154;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1155;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1156;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1157;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1158;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1159;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1160;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1161;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1162 = _GEN_525 | _GEN_526;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1163;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1164;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1165;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1166;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1167;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1168;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1169;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1170;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1171;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1172;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1173;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1174;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1175;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1176;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1177;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1178;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1179 = _GEN_532 | _GEN_533;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1180;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1181;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1182;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1183;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1184;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1185;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1186;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1187;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1188;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1189;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1190;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1191;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1192;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1193;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1194;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1195;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1196 = _GEN_539 | _GEN_540;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1197;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1198;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1199;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1200;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1201;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1202;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1203;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1204;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1205;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1206;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1207;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1208;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1209;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1210;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1211;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1212;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1213 = _GEN_546 | _GEN_547;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1214;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1215;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1216;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1217;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1218;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1219;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1220;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1221;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1222;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1223;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1224;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1225;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1226;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1227;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1228;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1229;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1230 = _GEN_553 | _GEN_554;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1231;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1232;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1233;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1234;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1235;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1236;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1237;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1238;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1239;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1240;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1241;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1242;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1243;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1244;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1245;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1246;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1247 = _GEN_560 | _GEN_561;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic        _GEN_1248;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1249;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1250;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1251;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1252;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1253;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1254;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1255;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1256;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1257;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1258;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1259;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1260;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1261;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1262;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1263;	// lsu.scala:1148:72, :1150:9
    automatic logic        _GEN_1264 = _GEN_567 | _GEN_568;	// lsu.scala:1149:106, :1150:9, :1154:46, :1156:60, :1157:9
    automatic logic [15:0] _GEN_1265 =
      {{_GEN_565 & _GEN_567},
       {_GEN_558 & _GEN_560},
       {_GEN_551 & _GEN_553},
       {_GEN_544 & _GEN_546},
       {_GEN_537 & _GEN_539},
       {_GEN_530 & _GEN_532},
       {_GEN_523 & _GEN_525},
       {_GEN_516 & _GEN_518},
       {_GEN_509 & _GEN_511},
       {_GEN_502 & _GEN_504},
       {_GEN_495 & _GEN_497},
       {_GEN_488 & _GEN_490},
       {_GEN_481 & _GEN_483},
       {_GEN_474 & _GEN_476},
       {_GEN_467 & _GEN_469},
       {_GEN_460 & _GEN_462}};	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1187:86
    automatic logic        mem_forward_valid_0;	// lsu.scala:1189:53
    automatic logic [4:0]  _l_idx_T_53;	// Mux.scala:47:69
    automatic logic [3:0]  l_idx;	// Mux.scala:47:69
    automatic logic        ld_xcpt_valid;	// lsu.scala:1238:44
    automatic logic        use_mem_xcpt;	// lsu.scala:1241:115
    automatic logic [11:0] xcpt_uop_br_mask;	// lsu.scala:1243:21
    automatic logic        _ldq_bits_succeeded_T =
      _io_core_exe_0_iresp_valid_output | _io_core_exe_0_fresp_valid_output;	// lsu.scala:1306:5, :1324:72, :1344:5, :1348:5
    automatic logic        _GEN_1266 = _GEN_600 & live;	// AMOALU.scala:10:17, lsu.scala:1369:24, util.scala:118:59
    automatic logic        _GEN_1267;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1268;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1269;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1270;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1271;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1272;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1273;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1274;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1275;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1276;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1277;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1278;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1279;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1280;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1281;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1282;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1283;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1284;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1285;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1286;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1287;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1288;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1289;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1290;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1291;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1292;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1293;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1294;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1295;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1296;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1297;	// lsu.scala:1306:5, :1348:5, :1369:33, :1370:35
    automatic logic        _GEN_1298;	// lsu.scala:1306:5, :1344:5, :1348:5
    automatic logic        _GEN_1299;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1300;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1301;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1302;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1303;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1304;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1305;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1306;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1307;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1308;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1309;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1310;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1311;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1312;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1313;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1314;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32
    automatic logic        _GEN_1315;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1316;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1317;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1318;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1319;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1320;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1321;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1322;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1323;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1324;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1325;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1326;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1327;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1328;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1329;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1330;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32
    automatic logic        _GEN_1331 = idx == 4'h0;	// lsu.scala:1453:18, :1456:31
    automatic logic        _GEN_1332 = commit_store & _GEN_1331;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1333 = idx == 4'h1;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1334 = commit_store & _GEN_1333;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1335 = idx == 4'h2;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1336 = commit_store & _GEN_1335;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1337 = idx == 4'h3;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1338 = commit_store & _GEN_1337;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1339 = idx == 4'h4;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1340 = commit_store & _GEN_1339;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1341 = idx == 4'h5;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1342 = commit_store & _GEN_1341;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1343 = idx == 4'h6;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1344 = commit_store & _GEN_1343;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1345 = idx == 4'h7;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1346 = commit_store & _GEN_1345;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1347 = idx == 4'h8;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1348 = commit_store & _GEN_1347;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1349 = idx == 4'h9;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1350 = commit_store & _GEN_1349;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1351 = idx == 4'hA;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1352 = commit_store & _GEN_1351;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1353 = idx == 4'hB;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1354 = commit_store & _GEN_1353;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1355 = idx == 4'hC;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1356 = commit_store & _GEN_1355;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1357 = idx == 4'hD;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1358 = commit_store & _GEN_1357;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1359 = idx == 4'hE;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1360 = commit_store & _GEN_1359;	// lsu.scala:304:5, :1451:49, :1455:5, :1456:31
    automatic logic        _GEN_1361 = commit_store & (&idx);	// lsu.scala:304:5, :1451:49, :1453:18, :1455:5, :1456:31
    automatic logic        _GEN_1362;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1363 = commit_store | ~commit_load;	// lsu.scala:1424:5, :1451:49, :1452:49, :1455:5, :1457:31
    automatic logic        _GEN_1364;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1365;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1366;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1367;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1368;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1369;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1370;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1371;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1372;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1373;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1374;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1375;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1376;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1377;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1378;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1462:38
    automatic logic        _GEN_1379 = commit_store | ~(commit_load & _GEN_1331);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1380 = commit_store | ~(commit_load & _GEN_1333);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1381 = commit_store | ~(commit_load & _GEN_1335);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1382 = commit_store | ~(commit_load & _GEN_1337);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1383 = commit_store | ~(commit_load & _GEN_1339);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1384 = commit_store | ~(commit_load & _GEN_1341);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1385 = commit_store | ~(commit_load & _GEN_1343);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1386 = commit_store | ~(commit_load & _GEN_1345);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1387 = commit_store | ~(commit_load & _GEN_1347);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1388 = commit_store | ~(commit_load & _GEN_1349);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1389 = commit_store | ~(commit_load & _GEN_1351);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1390 = commit_store | ~(commit_load & _GEN_1353);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1391 = commit_store | ~(commit_load & _GEN_1355);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1392 = commit_store | ~(commit_load & _GEN_1357);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1393 = commit_store | ~(commit_load & _GEN_1359);	// lsu.scala:1284:5, :1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1394 = commit_store | ~(commit_load & (&idx));	// lsu.scala:1284:5, :1451:49, :1452:49, :1453:18, :1455:5, :1456:31, :1457:31, :1464:38
    automatic logic        _GEN_1395 = idx_1 == 4'h0;	// lsu.scala:1453:18, :1456:31
    automatic logic        _GEN_1396 = idx_1 == 4'h1;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1397 = idx_1 == 4'h2;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1398 = idx_1 == 4'h3;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1399 = idx_1 == 4'h4;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1400 = idx_1 == 4'h5;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1401 = idx_1 == 4'h6;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1402 = idx_1 == 4'h7;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1403 = idx_1 == 4'h8;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1404 = idx_1 == 4'h9;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1405 = idx_1 == 4'hA;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1406 = idx_1 == 4'hB;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1407 = idx_1 == 4'hC;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1408 = idx_1 == 4'hD;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1409 = idx_1 == 4'hE;	// lsu.scala:305:44, :1453:18, :1456:31
    automatic logic        _GEN_1410 = commit_store_1 | ~(commit_load_1 & _GEN_1395);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1411 = commit_store_1 | ~(commit_load_1 & _GEN_1396);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1412 = commit_store_1 | ~(commit_load_1 & _GEN_1397);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1413 = commit_store_1 | ~(commit_load_1 & _GEN_1398);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1414 = commit_store_1 | ~(commit_load_1 & _GEN_1399);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1415 = commit_store_1 | ~(commit_load_1 & _GEN_1400);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1416 = commit_store_1 | ~(commit_load_1 & _GEN_1401);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1417 = commit_store_1 | ~(commit_load_1 & _GEN_1402);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1418 = commit_store_1 | ~(commit_load_1 & _GEN_1403);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1419 = commit_store_1 | ~(commit_load_1 & _GEN_1404);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1420 = commit_store_1 | ~(commit_load_1 & _GEN_1405);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1421 = commit_store_1 | ~(commit_load_1 & _GEN_1406);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1422 = commit_store_1 | ~(commit_load_1 & _GEN_1407);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1423 = commit_store_1 | ~(commit_load_1 & _GEN_1408);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1424 = commit_store_1 | ~(commit_load_1 & _GEN_1409);	// lsu.scala:1451:49, :1452:49, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1425 = commit_store_1 | ~(commit_load_1 & (&idx_1));	// lsu.scala:1451:49, :1452:49, :1453:18, :1455:5, :1456:31, :1457:31, :1462:38
    automatic logic        _GEN_1426;	// lsu.scala:1506:35
    automatic logic        _GEN_1427;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1428;	// lsu.scala:1506:35
    automatic logic        _GEN_1429;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1430;	// lsu.scala:1506:35
    automatic logic        _GEN_1431;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1432;	// lsu.scala:1506:35
    automatic logic        _GEN_1433;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1434;	// lsu.scala:1506:35
    automatic logic        _GEN_1435;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1436;	// lsu.scala:1506:35
    automatic logic        _GEN_1437;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1438;	// lsu.scala:1506:35
    automatic logic        _GEN_1439;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1440;	// lsu.scala:1506:35
    automatic logic        _GEN_1441;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1442;	// lsu.scala:1506:35
    automatic logic        _GEN_1443;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1444;	// lsu.scala:1506:35
    automatic logic        _GEN_1445;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1446;	// lsu.scala:1506:35
    automatic logic        _GEN_1447;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1448;	// lsu.scala:1506:35
    automatic logic        _GEN_1449;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1450;	// lsu.scala:1506:35
    automatic logic        _GEN_1451;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1452;	// lsu.scala:1506:35
    automatic logic        _GEN_1453;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1454;	// lsu.scala:1506:35
    automatic logic        _GEN_1455;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1456;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    automatic logic        _GEN_1457;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1458;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1459;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1460;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1461;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1462;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1463;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1464;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1465;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1466;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1467;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1468;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1469;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1470;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1471;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1472;	// lsu.scala:1306:5, :1505:3, :1509:35
    automatic logic        _GEN_1473;	// Decoupled.scala:40:37
    automatic logic        _GEN_1474;	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
    automatic logic        _GEN_1475;	// lsu.scala:244:34, :1527:34, :1533:38
    automatic logic        _GEN_1476;	// lsu.scala:1596:22
    automatic logic        _GEN_1477;	// lsu.scala:1505:3, :1597:3, :1602:5, :1603:16
    automatic logic        _GEN_1478;	// lsu.scala:1622:38
    automatic logic        _GEN_1479;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1480;	// lsu.scala:1622:38
    automatic logic        _GEN_1481;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1482;	// lsu.scala:1622:38
    automatic logic        _GEN_1483;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1484;	// lsu.scala:1622:38
    automatic logic        _GEN_1485;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1486;	// lsu.scala:1622:38
    automatic logic        _GEN_1487;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1488;	// lsu.scala:1622:38
    automatic logic        _GEN_1489;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1490;	// lsu.scala:1622:38
    automatic logic        _GEN_1491;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1492;	// lsu.scala:1622:38
    automatic logic        _GEN_1493;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1494;	// lsu.scala:1622:38
    automatic logic        _GEN_1495;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1496;	// lsu.scala:1622:38
    automatic logic        _GEN_1497;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1498;	// lsu.scala:1622:38
    automatic logic        _GEN_1499;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1500;	// lsu.scala:1622:38
    automatic logic        _GEN_1501;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1502;	// lsu.scala:1622:38
    automatic logic        _GEN_1503;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1504;	// lsu.scala:1622:38
    automatic logic        _GEN_1505;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1506;	// lsu.scala:1622:38
    automatic logic        _GEN_1507;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic        _GEN_1508;	// lsu.scala:1622:38
    automatic logic        _GEN_1509;	// lsu.scala:1505:3, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    automatic logic [4:0]  _ldq_retry_idx_idx_T_10;	// Mux.scala:47:69
    automatic logic [4:0]  _stq_retry_idx_idx_T_10;	// Mux.scala:47:69
    automatic logic [4:0]  _ldq_wakeup_idx_idx_T_10;	// Mux.scala:47:69
    _ldq_15_bits_st_dep_mask_T = 16'h1 << stq_head;	// lsu.scala:217:29, :260:71
    _GEN_642 = {16{~clear_store}};	// lsu.scala:260:33, :1495:3, :1500:17
    next_live_store_mask = (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & live_store_mask;	// lsu.scala:259:32, :260:{33,65,71}
    _GEN_643 = dis_ld_val & ldq_tail == 4'h0;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_644 = dis_ld_val & ldq_tail == 4'h1;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_645 = dis_ld_val & ldq_tail == 4'h2;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_646 = dis_ld_val & ldq_tail == 4'h3;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_647 = dis_ld_val & ldq_tail == 4'h4;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_648 = dis_ld_val & ldq_tail == 4'h5;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_649 = dis_ld_val & ldq_tail == 4'h6;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_650 = dis_ld_val & ldq_tail == 4'h7;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_651 = dis_ld_val & ldq_tail == 4'h8;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_652 = dis_ld_val & ldq_tail == 4'h9;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_653 = dis_ld_val & ldq_tail == 4'hA;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_654 = dis_ld_val & ldq_tail == 4'hB;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_655 = dis_ld_val & ldq_tail == 4'hC;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_656 = dis_ld_val & ldq_tail == 4'hD;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_657 = dis_ld_val & ldq_tail == 4'hE;	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_658 = dis_ld_val & (&ldq_tail);	// lsu.scala:210:16, :216:29, :301:85, :304:5, :305:44
    _GEN_659 = dis_st_val & stq_tail == 4'h0;	// lsu.scala:211:16, :218:29, :302:85, :321:5, :322:39
    _GEN_660 = dis_st_val & stq_tail == 4'h1;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_661 = dis_st_val & stq_tail == 4'h2;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_662 = dis_st_val & stq_tail == 4'h3;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_663 = dis_st_val & stq_tail == 4'h4;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_664 = dis_st_val & stq_tail == 4'h5;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_665 = dis_st_val & stq_tail == 4'h6;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_666 = dis_st_val & stq_tail == 4'h7;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_667 = dis_st_val & stq_tail == 4'h8;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_668 = dis_st_val & stq_tail == 4'h9;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_669 = dis_st_val & stq_tail == 4'hA;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_670 = dis_st_val & stq_tail == 4'hB;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_671 = dis_st_val & stq_tail == 4'hC;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_672 = dis_st_val & stq_tail == 4'hD;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_673 = dis_st_val & stq_tail == 4'hE;	// lsu.scala:211:16, :218:29, :302:85, :305:44, :321:5, :322:39
    _GEN_674 = dis_st_val & (&stq_tail);	// lsu.scala:211:16, :218:29, :302:85, :321:5, :322:39
    _GEN_675 = dis_ld_val | ~_GEN_659;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_676 = dis_ld_val | ~_GEN_660;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_677 = dis_ld_val | ~_GEN_661;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_678 = dis_ld_val | ~_GEN_662;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_679 = dis_ld_val | ~_GEN_663;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_680 = dis_ld_val | ~_GEN_664;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_681 = dis_ld_val | ~_GEN_665;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_682 = dis_ld_val | ~_GEN_666;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_683 = dis_ld_val | ~_GEN_667;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_684 = dis_ld_val | ~_GEN_668;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_685 = dis_ld_val | ~_GEN_669;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_686 = dis_ld_val | ~_GEN_670;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_687 = dis_ld_val | ~_GEN_671;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_688 = dis_ld_val | ~_GEN_672;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_689 = dis_ld_val | ~_GEN_673;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_690 = dis_ld_val | ~_GEN_674;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_691 = {16{dis_st_val}} & 16'h1 << stq_tail | next_live_store_mask;	// lsu.scala:218:29, :260:{33,71}, :302:85, :336:{31,72}
    _GEN_693 = _GEN_692 | _GEN_643;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_694 = dis_ld_val_1 ? _GEN_693 | ldq_0_valid : _GEN_643 | ldq_0_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_696 = _GEN_695 | _GEN_644;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_697 = dis_ld_val_1 ? _GEN_696 | ldq_1_valid : _GEN_644 | ldq_1_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_699 = _GEN_698 | _GEN_645;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_700 = dis_ld_val_1 ? _GEN_699 | ldq_2_valid : _GEN_645 | ldq_2_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_702 = _GEN_701 | _GEN_646;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_703 = dis_ld_val_1 ? _GEN_702 | ldq_3_valid : _GEN_646 | ldq_3_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_705 = _GEN_704 | _GEN_647;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_706 = dis_ld_val_1 ? _GEN_705 | ldq_4_valid : _GEN_647 | ldq_4_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_708 = _GEN_707 | _GEN_648;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_709 = dis_ld_val_1 ? _GEN_708 | ldq_5_valid : _GEN_648 | ldq_5_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_711 = _GEN_710 | _GEN_649;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_712 = dis_ld_val_1 ? _GEN_711 | ldq_6_valid : _GEN_649 | ldq_6_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_714 = _GEN_713 | _GEN_650;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_715 = dis_ld_val_1 ? _GEN_714 | ldq_7_valid : _GEN_650 | ldq_7_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_717 = _GEN_716 | _GEN_651;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_718 = dis_ld_val_1 ? _GEN_717 | ldq_8_valid : _GEN_651 | ldq_8_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_720 = _GEN_719 | _GEN_652;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_721 = dis_ld_val_1 ? _GEN_720 | ldq_9_valid : _GEN_652 | ldq_9_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_723 = _GEN_722 | _GEN_653;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_724 = dis_ld_val_1 ? _GEN_723 | ldq_10_valid : _GEN_653 | ldq_10_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_726 = _GEN_725 | _GEN_654;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_727 = dis_ld_val_1 ? _GEN_726 | ldq_11_valid : _GEN_654 | ldq_11_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_729 = _GEN_728 | _GEN_655;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_730 = dis_ld_val_1 ? _GEN_729 | ldq_12_valid : _GEN_655 | ldq_12_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_732 = _GEN_731 | _GEN_656;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_733 = dis_ld_val_1 ? _GEN_732 | ldq_13_valid : _GEN_656 | ldq_13_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_735 = _GEN_734 | _GEN_657;	// lsu.scala:210:16, :304:5, :305:44
    _GEN_736 = dis_ld_val_1 ? _GEN_735 | ldq_14_valid : _GEN_657 | ldq_14_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_737 = (&_GEN_98) | _GEN_658;	// lsu.scala:210:16, :304:5, :305:44, :333:21
    _GEN_738 = dis_ld_val_1 ? _GEN_737 | ldq_15_valid : _GEN_658 | ldq_15_valid;	// lsu.scala:210:16, :301:85, :304:5, :305:44
    _GEN_739 = dis_ld_val_1 & _GEN_692;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_740 = dis_ld_val_1 & _GEN_695;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_741 = dis_ld_val_1 & _GEN_698;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_742 = dis_ld_val_1 & _GEN_701;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_743 = dis_ld_val_1 & _GEN_704;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_744 = dis_ld_val_1 & _GEN_707;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_745 = dis_ld_val_1 & _GEN_710;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_746 = dis_ld_val_1 & _GEN_713;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_747 = dis_ld_val_1 & _GEN_716;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_748 = dis_ld_val_1 & _GEN_719;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_749 = dis_ld_val_1 & _GEN_722;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_750 = dis_ld_val_1 & _GEN_725;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_751 = dis_ld_val_1 & _GEN_728;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_752 = dis_ld_val_1 & _GEN_731;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_753 = dis_ld_val_1 & _GEN_734;	// lsu.scala:301:85, :304:5, :305:44, :306:44
    _GEN_754 = dis_ld_val_1 & (&_GEN_98);	// lsu.scala:301:85, :304:5, :305:44, :306:44, :333:21
    _GEN_755 = _GEN_739 | _GEN_643;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_756 = _GEN_740 | _GEN_644;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_757 = _GEN_741 | _GEN_645;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_758 = _GEN_742 | _GEN_646;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_759 = _GEN_743 | _GEN_647;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_760 = _GEN_744 | _GEN_648;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_761 = _GEN_745 | _GEN_649;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_762 = _GEN_746 | _GEN_650;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_763 = _GEN_747 | _GEN_651;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_764 = _GEN_748 | _GEN_652;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_765 = _GEN_749 | _GEN_653;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_766 = _GEN_750 | _GEN_654;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_767 = _GEN_751 | _GEN_655;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_768 = _GEN_752 | _GEN_656;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_769 = _GEN_753 | _GEN_657;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_770 = _GEN_754 | _GEN_658;	// lsu.scala:210:16, :304:5, :305:44, :306:44
    _GEN_771 =
      dis_ld_val_1
        ? ~_GEN_693 & ldq_0_bits_order_fail
        : ~_GEN_643 & ldq_0_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_772 =
      dis_ld_val_1
        ? ~_GEN_696 & ldq_1_bits_order_fail
        : ~_GEN_644 & ldq_1_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_773 =
      dis_ld_val_1
        ? ~_GEN_699 & ldq_2_bits_order_fail
        : ~_GEN_645 & ldq_2_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_774 =
      dis_ld_val_1
        ? ~_GEN_702 & ldq_3_bits_order_fail
        : ~_GEN_646 & ldq_3_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_775 =
      dis_ld_val_1
        ? ~_GEN_705 & ldq_4_bits_order_fail
        : ~_GEN_647 & ldq_4_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_776 =
      dis_ld_val_1
        ? ~_GEN_708 & ldq_5_bits_order_fail
        : ~_GEN_648 & ldq_5_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_777 =
      dis_ld_val_1
        ? ~_GEN_711 & ldq_6_bits_order_fail
        : ~_GEN_649 & ldq_6_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_778 =
      dis_ld_val_1
        ? ~_GEN_714 & ldq_7_bits_order_fail
        : ~_GEN_650 & ldq_7_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_779 =
      dis_ld_val_1
        ? ~_GEN_717 & ldq_8_bits_order_fail
        : ~_GEN_651 & ldq_8_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_780 =
      dis_ld_val_1
        ? ~_GEN_720 & ldq_9_bits_order_fail
        : ~_GEN_652 & ldq_9_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_781 =
      dis_ld_val_1
        ? ~_GEN_723 & ldq_10_bits_order_fail
        : ~_GEN_653 & ldq_10_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_782 =
      dis_ld_val_1
        ? ~_GEN_726 & ldq_11_bits_order_fail
        : ~_GEN_654 & ldq_11_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_783 =
      dis_ld_val_1
        ? ~_GEN_729 & ldq_12_bits_order_fail
        : ~_GEN_655 & ldq_12_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_784 =
      dis_ld_val_1
        ? ~_GEN_732 & ldq_13_bits_order_fail
        : ~_GEN_656 & ldq_13_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_785 =
      dis_ld_val_1
        ? ~_GEN_735 & ldq_14_bits_order_fail
        : ~_GEN_657 & ldq_14_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_786 =
      dis_ld_val_1
        ? ~_GEN_737 & ldq_15_bits_order_fail
        : ~_GEN_658 & ldq_15_bits_order_fail;	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :313:44
    _GEN_787 = dis_st_val_1 & _GEN_99 == 4'h0;	// lsu.scala:302:85, :304:5, :321:5, :322:39, :338:21
    _GEN_788 = ~dis_ld_val_1 & _GEN_787 | ~dis_ld_val & _GEN_659 | stq_0_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_789 = dis_st_val_1 & _GEN_99 == 4'h1;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_790 = ~dis_ld_val_1 & _GEN_789 | ~dis_ld_val & _GEN_660 | stq_1_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_791 = dis_st_val_1 & _GEN_99 == 4'h2;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_792 = ~dis_ld_val_1 & _GEN_791 | ~dis_ld_val & _GEN_661 | stq_2_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_793 = dis_st_val_1 & _GEN_99 == 4'h3;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_794 = ~dis_ld_val_1 & _GEN_793 | ~dis_ld_val & _GEN_662 | stq_3_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_795 = dis_st_val_1 & _GEN_99 == 4'h4;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_796 = ~dis_ld_val_1 & _GEN_795 | ~dis_ld_val & _GEN_663 | stq_4_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_797 = dis_st_val_1 & _GEN_99 == 4'h5;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_798 = ~dis_ld_val_1 & _GEN_797 | ~dis_ld_val & _GEN_664 | stq_5_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_799 = dis_st_val_1 & _GEN_99 == 4'h6;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_800 = ~dis_ld_val_1 & _GEN_799 | ~dis_ld_val & _GEN_665 | stq_6_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_801 = dis_st_val_1 & _GEN_99 == 4'h7;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_802 = ~dis_ld_val_1 & _GEN_801 | ~dis_ld_val & _GEN_666 | stq_7_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_803 = dis_st_val_1 & _GEN_99 == 4'h8;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_804 = ~dis_ld_val_1 & _GEN_803 | ~dis_ld_val & _GEN_667 | stq_8_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_805 = dis_st_val_1 & _GEN_99 == 4'h9;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_806 = ~dis_ld_val_1 & _GEN_805 | ~dis_ld_val & _GEN_668 | stq_9_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_807 = dis_st_val_1 & _GEN_99 == 4'hA;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_808 = ~dis_ld_val_1 & _GEN_807 | ~dis_ld_val & _GEN_669 | stq_10_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_809 = dis_st_val_1 & _GEN_99 == 4'hB;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_810 = ~dis_ld_val_1 & _GEN_809 | ~dis_ld_val & _GEN_670 | stq_11_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_811 = dis_st_val_1 & _GEN_99 == 4'hC;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_812 = ~dis_ld_val_1 & _GEN_811 | ~dis_ld_val & _GEN_671 | stq_12_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_813 = dis_st_val_1 & _GEN_99 == 4'hD;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_814 = ~dis_ld_val_1 & _GEN_813 | ~dis_ld_val & _GEN_672 | stq_13_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_815 = dis_st_val_1 & _GEN_99 == 4'hE;	// lsu.scala:302:85, :304:5, :305:44, :321:5, :322:39, :338:21
    _GEN_816 = ~dis_ld_val_1 & _GEN_815 | ~dis_ld_val & _GEN_673 | stq_14_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_817 = dis_st_val_1 & (&_GEN_99);	// lsu.scala:302:85, :304:5, :321:5, :322:39, :338:21
    _GEN_818 = ~dis_ld_val_1 & _GEN_817 | ~dis_ld_val & _GEN_674 | stq_15_valid;	// lsu.scala:211:16, :301:85, :304:5, :321:5, :322:39
    _GEN_819 = dis_ld_val_1 | ~_GEN_787;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_820 = dis_ld_val_1 | ~_GEN_789;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_821 = dis_ld_val_1 | ~_GEN_791;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_822 = dis_ld_val_1 | ~_GEN_793;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_823 = dis_ld_val_1 | ~_GEN_795;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_824 = dis_ld_val_1 | ~_GEN_797;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_825 = dis_ld_val_1 | ~_GEN_799;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_826 = dis_ld_val_1 | ~_GEN_801;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_827 = dis_ld_val_1 | ~_GEN_803;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_828 = dis_ld_val_1 | ~_GEN_805;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_829 = dis_ld_val_1 | ~_GEN_807;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_830 = dis_ld_val_1 | ~_GEN_809;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_831 = dis_ld_val_1 | ~_GEN_811;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_832 = dis_ld_val_1 | ~_GEN_813;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_833 = dis_ld_val_1 | ~_GEN_815;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_834 = dis_ld_val_1 | ~_GEN_817;	// lsu.scala:301:85, :304:5, :321:5, :322:39
    _GEN_835 = _GEN_819 & _GEN_675 & stq_0_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_836 = _GEN_820 & _GEN_676 & stq_1_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_837 = _GEN_821 & _GEN_677 & stq_2_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_838 = _GEN_822 & _GEN_678 & stq_3_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_839 = _GEN_823 & _GEN_679 & stq_4_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_840 = _GEN_824 & _GEN_680 & stq_5_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_841 = _GEN_825 & _GEN_681 & stq_6_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_842 = _GEN_826 & _GEN_682 & stq_7_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_843 = _GEN_827 & _GEN_683 & stq_8_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_844 = _GEN_828 & _GEN_684 & stq_9_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_845 = _GEN_829 & _GEN_685 & stq_10_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_846 = _GEN_830 & _GEN_686 & stq_11_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_847 = _GEN_831 & _GEN_687 & stq_12_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_848 = _GEN_832 & _GEN_688 & stq_13_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_849 = _GEN_833 & _GEN_689 & stq_14_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    _GEN_850 = _GEN_834 & _GEN_690 & stq_15_bits_committed;	// lsu.scala:211:16, :304:5, :321:5
    ldq_retry_idx_block =
      (will_fire_load_wakeup_0
         ? _GEN_208
         : can_fire_load_incoming_0 ? _GEN_223 : _GEN_239) | p1_block_load_mask_0;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_2 =
      ldq_0_bits_addr_valid & ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_1 =
      (will_fire_load_wakeup_0
         ? _GEN_209
         : can_fire_load_incoming_0 ? _GEN_224 : _GEN_241) | p1_block_load_mask_1;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_5 =
      ldq_1_bits_addr_valid & ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_2 =
      (will_fire_load_wakeup_0
         ? _GEN_210
         : can_fire_load_incoming_0 ? _GEN_225 : _GEN_243) | p1_block_load_mask_2;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_8 =
      ldq_2_bits_addr_valid & ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_3 =
      (will_fire_load_wakeup_0
         ? _GEN_211
         : can_fire_load_incoming_0 ? _GEN_226 : _GEN_245) | p1_block_load_mask_3;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_11 =
      ldq_3_bits_addr_valid & ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_4 =
      (will_fire_load_wakeup_0
         ? _GEN_212
         : can_fire_load_incoming_0 ? _GEN_227 : _GEN_247) | p1_block_load_mask_4;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_14 =
      ldq_4_bits_addr_valid & ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_5 =
      (will_fire_load_wakeup_0
         ? _GEN_213
         : can_fire_load_incoming_0 ? _GEN_228 : _GEN_249) | p1_block_load_mask_5;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_17 =
      ldq_5_bits_addr_valid & ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_6 =
      (will_fire_load_wakeup_0
         ? _GEN_214
         : can_fire_load_incoming_0 ? _GEN_229 : _GEN_251) | p1_block_load_mask_6;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_20 =
      ldq_6_bits_addr_valid & ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_7 =
      (will_fire_load_wakeup_0
         ? _GEN_215
         : can_fire_load_incoming_0 ? _GEN_230 : _GEN_253) | p1_block_load_mask_7;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_23 =
      ldq_7_bits_addr_valid & ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_8 =
      (will_fire_load_wakeup_0
         ? _GEN_216
         : can_fire_load_incoming_0 ? _GEN_231 : _GEN_255) | p1_block_load_mask_8;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_26 =
      ldq_8_bits_addr_valid & ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_9 =
      (will_fire_load_wakeup_0
         ? _GEN_217
         : can_fire_load_incoming_0 ? _GEN_232 : _GEN_257) | p1_block_load_mask_9;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_29 =
      ldq_9_bits_addr_valid & ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_10 =
      (will_fire_load_wakeup_0
         ? _GEN_218
         : can_fire_load_incoming_0 ? _GEN_233 : _GEN_259) | p1_block_load_mask_10;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_32 =
      ldq_10_bits_addr_valid & ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_11 =
      (will_fire_load_wakeup_0
         ? _GEN_219
         : can_fire_load_incoming_0 ? _GEN_234 : _GEN_261) | p1_block_load_mask_11;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_35 =
      ldq_11_bits_addr_valid & ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_12 =
      (will_fire_load_wakeup_0
         ? _GEN_220
         : can_fire_load_incoming_0 ? _GEN_235 : _GEN_263) | p1_block_load_mask_12;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_38 =
      ldq_12_bits_addr_valid & ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_13 =
      (will_fire_load_wakeup_0
         ? _GEN_221
         : can_fire_load_incoming_0 ? _GEN_236 : _GEN_265) | p1_block_load_mask_13;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_41 =
      ldq_13_bits_addr_valid & ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_14 =
      (will_fire_load_wakeup_0
         ? _GEN_222
         : can_fire_load_incoming_0 ? _GEN_237 : _GEN_267) | p1_block_load_mask_14;	// lsu.scala:398:35, :417:36, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _ldq_retry_idx_T_44 =
      ldq_14_bits_addr_valid & ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;	// lsu.scala:210:16, :417:36, :418:{39,42}
    ldq_retry_idx_block_15 =
      (will_fire_load_wakeup_0
         ? (&ldq_wakeup_idx)
         : can_fire_load_incoming_0 ? (&io_core_exe_0_req_bits_uop_ldq_idx) : _GEN_268)
      | p1_block_load_mask_15;	// lsu.scala:398:35, :417:36, :430:31, :441:63, :535:65, :569:37, :570:49, :571:46, :572:52, :573:43, :574:49
    _temp_bits_T = ldq_head == 4'h0;	// lsu.scala:215:29, util.scala:351:72
    _temp_bits_T_2 = ldq_head < 4'h2;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_4 = ldq_head < 4'h3;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_6 = ldq_head < 4'h4;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_8 = ldq_head < 4'h5;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_10 = ldq_head < 4'h6;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_12 = ldq_head < 4'h7;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_16 = ldq_head < 4'h9;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_18 = ldq_head < 4'hA;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_20 = ldq_head < 4'hB;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_22 = ldq_head[3:2] != 2'h3;	// lsu.scala:215:29, util.scala:351:72
    _temp_bits_T_24 = ldq_head < 4'hD;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _temp_bits_T_26 = ldq_head[3:1] != 3'h7;	// lsu.scala:215:29, util.scala:351:72
    _temp_bits_T_28 = ldq_head != 4'hF;	// lsu.scala:215:29, :305:44, util.scala:351:72
    _stq_retry_idx_T = stq_0_bits_addr_valid & stq_0_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_1 = stq_1_bits_addr_valid & stq_1_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_2 = stq_2_bits_addr_valid & stq_2_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_3 = stq_3_bits_addr_valid & stq_3_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_4 = stq_4_bits_addr_valid & stq_4_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_5 = stq_5_bits_addr_valid & stq_5_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_6 = stq_6_bits_addr_valid & stq_6_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_7 = stq_7_bits_addr_valid & stq_7_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_8 = stq_8_bits_addr_valid & stq_8_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_9 = stq_9_bits_addr_valid & stq_9_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_10 = stq_10_bits_addr_valid & stq_10_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_11 = stq_11_bits_addr_valid & stq_11_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_12 = stq_12_bits_addr_valid & stq_12_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_13 = stq_13_bits_addr_valid & stq_13_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _stq_retry_idx_T_14 = stq_14_bits_addr_valid & stq_14_bits_addr_is_virtual;	// lsu.scala:211:16, :424:18
    _ldq_wakeup_idx_T_7 =
      ldq_0_bits_addr_valid & ~ldq_0_bits_executed & ~ldq_0_bits_succeeded
      & ~ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_15 =
      ldq_1_bits_addr_valid & ~ldq_1_bits_executed & ~ldq_1_bits_succeeded
      & ~ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_23 =
      ldq_2_bits_addr_valid & ~ldq_2_bits_executed & ~ldq_2_bits_succeeded
      & ~ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_31 =
      ldq_3_bits_addr_valid & ~ldq_3_bits_executed & ~ldq_3_bits_succeeded
      & ~ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_39 =
      ldq_4_bits_addr_valid & ~ldq_4_bits_executed & ~ldq_4_bits_succeeded
      & ~ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_47 =
      ldq_5_bits_addr_valid & ~ldq_5_bits_executed & ~ldq_5_bits_succeeded
      & ~ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_55 =
      ldq_6_bits_addr_valid & ~ldq_6_bits_executed & ~ldq_6_bits_succeeded
      & ~ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_63 =
      ldq_7_bits_addr_valid & ~ldq_7_bits_executed & ~ldq_7_bits_succeeded
      & ~ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_71 =
      ldq_8_bits_addr_valid & ~ldq_8_bits_executed & ~ldq_8_bits_succeeded
      & ~ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_79 =
      ldq_9_bits_addr_valid & ~ldq_9_bits_executed & ~ldq_9_bits_succeeded
      & ~ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_87 =
      ldq_10_bits_addr_valid & ~ldq_10_bits_executed & ~ldq_10_bits_succeeded
      & ~ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_95 =
      ldq_11_bits_addr_valid & ~ldq_11_bits_executed & ~ldq_11_bits_succeeded
      & ~ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_103 =
      ldq_12_bits_addr_valid & ~ldq_12_bits_executed & ~ldq_12_bits_succeeded
      & ~ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_111 =
      ldq_13_bits_addr_valid & ~ldq_13_bits_executed & ~ldq_13_bits_succeeded
      & ~ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    _ldq_wakeup_idx_T_119 =
      ldq_14_bits_addr_valid & ~ldq_14_bits_executed & ~ldq_14_bits_succeeded
      & ~ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;	// lsu.scala:210:16, :417:36, :433:{21,36,52,71,74}
    ma_st_0 = _stq_idx_T & io_core_exe_0_req_bits_mxcpt_valid;	// lsu.scala:660:{56,87}
    pf_ld_0 =
      ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_ld
      & _mem_xcpt_uops_WIRE_0_uses_ldq;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :661:75
    pf_st_0 =
      ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_st
      & _mem_xcpt_uops_WIRE_0_uses_stq;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :662:75
    ae_ld_0 =
      ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_ae_ld
      & _mem_xcpt_uops_WIRE_0_uses_ldq;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :663:75
    dmem_req_fire_0 = dmem_req_0_valid & io_dmem_req_ready;	// lsu.scala:752:55, :766:39, :767:30, :773:43
    ldq_idx =
      can_fire_load_incoming_0 ? io_core_exe_0_req_bits_uop_ldq_idx : ldq_retry_idx;	// lsu.scala:415:30, :441:63, :837:24
    _GEN_851 = _GEN_272 & ldq_idx == 4'h0;	// lsu.scala:220:29, :304:5, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_852 =
      _GEN_851
      | (dis_ld_val_1
           ? ~_GEN_693 & ldq_0_bits_addr_valid
           : ~_GEN_643 & ldq_0_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_853 = _GEN_272 & ldq_idx == 4'h1;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_854 =
      _GEN_853
      | (dis_ld_val_1
           ? ~_GEN_696 & ldq_1_bits_addr_valid
           : ~_GEN_644 & ldq_1_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_855 = _GEN_272 & ldq_idx == 4'h2;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_856 =
      _GEN_855
      | (dis_ld_val_1
           ? ~_GEN_699 & ldq_2_bits_addr_valid
           : ~_GEN_645 & ldq_2_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_857 = _GEN_272 & ldq_idx == 4'h3;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_858 =
      _GEN_857
      | (dis_ld_val_1
           ? ~_GEN_702 & ldq_3_bits_addr_valid
           : ~_GEN_646 & ldq_3_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_859 = _GEN_272 & ldq_idx == 4'h4;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_860 =
      _GEN_859
      | (dis_ld_val_1
           ? ~_GEN_705 & ldq_4_bits_addr_valid
           : ~_GEN_647 & ldq_4_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_861 = _GEN_272 & ldq_idx == 4'h5;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_862 =
      _GEN_861
      | (dis_ld_val_1
           ? ~_GEN_708 & ldq_5_bits_addr_valid
           : ~_GEN_648 & ldq_5_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_863 = _GEN_272 & ldq_idx == 4'h6;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_864 =
      _GEN_863
      | (dis_ld_val_1
           ? ~_GEN_711 & ldq_6_bits_addr_valid
           : ~_GEN_649 & ldq_6_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_865 = _GEN_272 & ldq_idx == 4'h7;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_866 =
      _GEN_865
      | (dis_ld_val_1
           ? ~_GEN_714 & ldq_7_bits_addr_valid
           : ~_GEN_650 & ldq_7_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_867 = _GEN_272 & ldq_idx == 4'h8;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_868 =
      _GEN_867
      | (dis_ld_val_1
           ? ~_GEN_717 & ldq_8_bits_addr_valid
           : ~_GEN_651 & ldq_8_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_869 = _GEN_272 & ldq_idx == 4'h9;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_870 =
      _GEN_869
      | (dis_ld_val_1
           ? ~_GEN_720 & ldq_9_bits_addr_valid
           : ~_GEN_652 & ldq_9_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_871 = _GEN_272 & ldq_idx == 4'hA;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_872 =
      _GEN_871
      | (dis_ld_val_1
           ? ~_GEN_723 & ldq_10_bits_addr_valid
           : ~_GEN_653 & ldq_10_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_873 = _GEN_272 & ldq_idx == 4'hB;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_874 =
      _GEN_873
      | (dis_ld_val_1
           ? ~_GEN_726 & ldq_11_bits_addr_valid
           : ~_GEN_654 & ldq_11_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_875 = _GEN_272 & ldq_idx == 4'hC;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_876 =
      _GEN_875
      | (dis_ld_val_1
           ? ~_GEN_729 & ldq_12_bits_addr_valid
           : ~_GEN_655 & ldq_12_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_877 = _GEN_272 & ldq_idx == 4'hD;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_878 =
      _GEN_877
      | (dis_ld_val_1
           ? ~_GEN_732 & ldq_13_bits_addr_valid
           : ~_GEN_656 & ldq_13_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_879 = _GEN_272 & ldq_idx == 4'hE;	// lsu.scala:220:29, :304:5, :305:44, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_880 =
      _GEN_879
      | (dis_ld_val_1
           ? ~_GEN_735 & ldq_14_bits_addr_valid
           : ~_GEN_657 & ldq_14_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _GEN_881 = _GEN_272 & (&ldq_idx);	// lsu.scala:220:29, :304:5, :766:39, :773:43, :780:45, :836:5, :837:24, :838:45
    _GEN_882 =
      _GEN_881
      | (dis_ld_val_1
           ? ~_GEN_737 & ldq_15_bits_addr_valid
           : ~_GEN_658 & ldq_15_bits_addr_valid);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :836:5, :838:45
    _ldq_bits_addr_is_uncacheable_T_1 = ~_dtlb_io_resp_0_cacheable & ~exe_tlb_miss_0;	// lsu.scala:249:20, :708:58, :711:43, :842:{71,74}
    stq_idx = _stq_idx_T ? io_core_exe_0_req_bits_uop_stq_idx : stq_retry_idx;	// lsu.scala:422:30, :660:56, :850:24
    _GEN_883 = _GEN_278 & stq_idx == 4'h0;	// lsu.scala:304:5, :848:67, :849:5, :850:24, :853:36
    _GEN_884 = _GEN_883 ? ~pf_st_0 : _GEN_819 & _GEN_675 & stq_0_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_885 = _GEN_278 & stq_idx == 4'h1;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_886 = _GEN_885 ? ~pf_st_0 : _GEN_820 & _GEN_676 & stq_1_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_887 = _GEN_278 & stq_idx == 4'h2;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_888 = _GEN_887 ? ~pf_st_0 : _GEN_821 & _GEN_677 & stq_2_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_889 = _GEN_278 & stq_idx == 4'h3;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_890 = _GEN_889 ? ~pf_st_0 : _GEN_822 & _GEN_678 & stq_3_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_891 = _GEN_278 & stq_idx == 4'h4;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_892 = _GEN_891 ? ~pf_st_0 : _GEN_823 & _GEN_679 & stq_4_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_893 = _GEN_278 & stq_idx == 4'h5;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_894 = _GEN_893 ? ~pf_st_0 : _GEN_824 & _GEN_680 & stq_5_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_895 = _GEN_278 & stq_idx == 4'h6;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_896 = _GEN_895 ? ~pf_st_0 : _GEN_825 & _GEN_681 & stq_6_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_897 = _GEN_278 & stq_idx == 4'h7;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_898 = _GEN_897 ? ~pf_st_0 : _GEN_826 & _GEN_682 & stq_7_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_899 = _GEN_278 & stq_idx == 4'h8;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_900 = _GEN_899 ? ~pf_st_0 : _GEN_827 & _GEN_683 & stq_8_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_901 = _GEN_278 & stq_idx == 4'h9;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_902 = _GEN_901 ? ~pf_st_0 : _GEN_828 & _GEN_684 & stq_9_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_903 = _GEN_278 & stq_idx == 4'hA;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_904 = _GEN_903 ? ~pf_st_0 : _GEN_829 & _GEN_685 & stq_10_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_905 = _GEN_278 & stq_idx == 4'hB;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_906 = _GEN_905 ? ~pf_st_0 : _GEN_830 & _GEN_686 & stq_11_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_907 = _GEN_278 & stq_idx == 4'hC;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_908 = _GEN_907 ? ~pf_st_0 : _GEN_831 & _GEN_687 & stq_12_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_909 = _GEN_278 & stq_idx == 4'hD;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_910 = _GEN_909 ? ~pf_st_0 : _GEN_832 & _GEN_688 & stq_13_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_911 = _GEN_278 & stq_idx == 4'hE;	// lsu.scala:304:5, :305:44, :848:67, :849:5, :850:24, :853:36
    _GEN_912 = _GEN_911 ? ~pf_st_0 : _GEN_833 & _GEN_689 & stq_14_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_913 = _GEN_278 & (&stq_idx);	// lsu.scala:304:5, :848:67, :849:5, :850:24, :853:36
    _GEN_914 = _GEN_913 ? ~pf_st_0 : _GEN_834 & _GEN_690 & stq_15_bits_addr_valid;	// lsu.scala:211:16, :304:5, :321:5, :662:75, :849:5, :853:{36,39}
    _GEN_916 = _GEN_915 | _GEN_819 & _GEN_675 & stq_0_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_918 = _GEN_917 | _GEN_820 & _GEN_676 & stq_1_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_920 = _GEN_919 | _GEN_821 & _GEN_677 & stq_2_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_922 = _GEN_921 | _GEN_822 & _GEN_678 & stq_3_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_924 = _GEN_923 | _GEN_823 & _GEN_679 & stq_4_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_926 = _GEN_925 | _GEN_824 & _GEN_680 & stq_5_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_928 = _GEN_927 | _GEN_825 & _GEN_681 & stq_6_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_930 = _GEN_929 | _GEN_826 & _GEN_682 & stq_7_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_932 = _GEN_931 | _GEN_827 & _GEN_683 & stq_8_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_934 = _GEN_933 | _GEN_828 & _GEN_684 & stq_9_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_936 = _GEN_935 | _GEN_829 & _GEN_685 & stq_10_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_938 = _GEN_937 | _GEN_830 & _GEN_686 & stq_11_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_940 = _GEN_939 | _GEN_831 & _GEN_687 & stq_12_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_942 = _GEN_941 | _GEN_832 & _GEN_688 & stq_13_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_944 = _GEN_943 | _GEN_833 & _GEN_689 & stq_14_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    _GEN_946 = _GEN_945 | _GEN_834 & _GEN_690 & stq_15_bits_data_valid;	// lsu.scala:211:16, :304:5, :321:5, :869:5, :873:33
    l_forward_stq_idx =
      l_forwarders_0 ? wb_forward_stq_idx_0 : ldq_0_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_947 =
      ~ldq_0_bits_forward_std_val | l_forward_stq_idx != lcam_stq_idx_0
      & (l_forward_stq_idx < lcam_stq_idx_0
         ^ l_forward_stq_idx < ldq_0_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_0_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_948 = _GEN_286 & ~s1_executing_loads_0 & ldq_0_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_16 =
      ~_GEN_284 & (_GEN_289 ? _GEN_947 : _GEN_290 & searcher_is_older & _GEN_948);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_1 =
      l_forwarders_1_0 ? wb_forward_stq_idx_0 : ldq_1_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_963 =
      ~ldq_1_bits_forward_std_val | l_forward_stq_idx_1 != lcam_stq_idx_0
      & (l_forward_stq_idx_1 < lcam_stq_idx_0
         ^ l_forward_stq_idx_1 < ldq_1_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_1_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_964 = _GEN_297 & ~s1_executing_loads_1 & ldq_1_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_17 =
      ~_GEN_295 & (_GEN_299 ? _GEN_963 : _GEN_300 & searcher_is_older_1 & _GEN_964);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_2 =
      l_forwarders_2_0 ? wb_forward_stq_idx_0 : ldq_2_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_965 =
      ~ldq_2_bits_forward_std_val | l_forward_stq_idx_2 != lcam_stq_idx_0
      & (l_forward_stq_idx_2 < lcam_stq_idx_0
         ^ l_forward_stq_idx_2 < ldq_2_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_2_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_966 = _GEN_308 & ~s1_executing_loads_2 & ldq_2_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_18 =
      ~_GEN_306 & (_GEN_310 ? _GEN_965 : _GEN_311 & searcher_is_older_2 & _GEN_966);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_3 =
      l_forwarders_3_0 ? wb_forward_stq_idx_0 : ldq_3_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_967 =
      ~ldq_3_bits_forward_std_val | l_forward_stq_idx_3 != lcam_stq_idx_0
      & (l_forward_stq_idx_3 < lcam_stq_idx_0
         ^ l_forward_stq_idx_3 < ldq_3_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_3_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_968 = _GEN_319 & ~s1_executing_loads_3 & ldq_3_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_19 =
      ~_GEN_317 & (_GEN_321 ? _GEN_967 : _GEN_322 & searcher_is_older_3 & _GEN_968);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_4 =
      l_forwarders_4_0 ? wb_forward_stq_idx_0 : ldq_4_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_969 =
      ~ldq_4_bits_forward_std_val | l_forward_stq_idx_4 != lcam_stq_idx_0
      & (l_forward_stq_idx_4 < lcam_stq_idx_0
         ^ l_forward_stq_idx_4 < ldq_4_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_4_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_970 = _GEN_330 & ~s1_executing_loads_4 & ldq_4_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_20 =
      ~_GEN_328 & (_GEN_332 ? _GEN_969 : _GEN_333 & searcher_is_older_4 & _GEN_970);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_5 =
      l_forwarders_5_0 ? wb_forward_stq_idx_0 : ldq_5_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_971 =
      ~ldq_5_bits_forward_std_val | l_forward_stq_idx_5 != lcam_stq_idx_0
      & (l_forward_stq_idx_5 < lcam_stq_idx_0
         ^ l_forward_stq_idx_5 < ldq_5_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_5_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_972 = _GEN_341 & ~s1_executing_loads_5 & ldq_5_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_21 =
      ~_GEN_339 & (_GEN_343 ? _GEN_971 : _GEN_344 & searcher_is_older_5 & _GEN_972);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_6 =
      l_forwarders_6_0 ? wb_forward_stq_idx_0 : ldq_6_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_973 =
      ~ldq_6_bits_forward_std_val | l_forward_stq_idx_6 != lcam_stq_idx_0
      & (l_forward_stq_idx_6 < lcam_stq_idx_0
         ^ l_forward_stq_idx_6 < ldq_6_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_6_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_974 = _GEN_352 & ~s1_executing_loads_6 & ldq_6_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_22 =
      ~_GEN_350 & (_GEN_354 ? _GEN_973 : _GEN_355 & searcher_is_older_6 & _GEN_974);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_7 =
      l_forwarders_7_0 ? wb_forward_stq_idx_0 : ldq_7_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_975 =
      ~ldq_7_bits_forward_std_val | l_forward_stq_idx_7 != lcam_stq_idx_0
      & (l_forward_stq_idx_7 < lcam_stq_idx_0
         ^ l_forward_stq_idx_7 < ldq_7_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_7_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_976 = _GEN_363 & ~s1_executing_loads_7 & ldq_7_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_23 =
      ~_GEN_361 & (_GEN_365 ? _GEN_975 : _GEN_366 & searcher_is_older_7 & _GEN_976);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_8 =
      l_forwarders_8_0 ? wb_forward_stq_idx_0 : ldq_8_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_977 =
      ~ldq_8_bits_forward_std_val | l_forward_stq_idx_8 != lcam_stq_idx_0
      & (l_forward_stq_idx_8 < lcam_stq_idx_0
         ^ l_forward_stq_idx_8 < ldq_8_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_8_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_978 = _GEN_374 & ~s1_executing_loads_8 & ldq_8_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_24 =
      ~_GEN_372 & (_GEN_376 ? _GEN_977 : _GEN_377 & searcher_is_older_8 & _GEN_978);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_9 =
      l_forwarders_9_0 ? wb_forward_stq_idx_0 : ldq_9_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_979 =
      ~ldq_9_bits_forward_std_val | l_forward_stq_idx_9 != lcam_stq_idx_0
      & (l_forward_stq_idx_9 < lcam_stq_idx_0
         ^ l_forward_stq_idx_9 < ldq_9_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_9_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_980 = _GEN_385 & ~s1_executing_loads_9 & ldq_9_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_25 =
      ~_GEN_383 & (_GEN_387 ? _GEN_979 : _GEN_388 & searcher_is_older_9 & _GEN_980);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_10 =
      l_forwarders_10_0 ? wb_forward_stq_idx_0 : ldq_10_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_981 =
      ~ldq_10_bits_forward_std_val | l_forward_stq_idx_10 != lcam_stq_idx_0
      & (l_forward_stq_idx_10 < lcam_stq_idx_0
         ^ l_forward_stq_idx_10 < ldq_10_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_10_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_982 = _GEN_396 & ~s1_executing_loads_10 & ldq_10_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_26 =
      ~_GEN_394 & (_GEN_398 ? _GEN_981 : _GEN_399 & searcher_is_older_10 & _GEN_982);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_11 =
      l_forwarders_11_0 ? wb_forward_stq_idx_0 : ldq_11_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_983 =
      ~ldq_11_bits_forward_std_val | l_forward_stq_idx_11 != lcam_stq_idx_0
      & (l_forward_stq_idx_11 < lcam_stq_idx_0
         ^ l_forward_stq_idx_11 < ldq_11_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_11_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_984 = _GEN_407 & ~s1_executing_loads_11 & ldq_11_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_27 =
      ~_GEN_405 & (_GEN_409 ? _GEN_983 : _GEN_410 & searcher_is_older_11 & _GEN_984);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_12 =
      l_forwarders_12_0 ? wb_forward_stq_idx_0 : ldq_12_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_985 =
      ~ldq_12_bits_forward_std_val | l_forward_stq_idx_12 != lcam_stq_idx_0
      & (l_forward_stq_idx_12 < lcam_stq_idx_0
         ^ l_forward_stq_idx_12 < ldq_12_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_12_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_986 = _GEN_418 & ~s1_executing_loads_12 & ldq_12_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_28 =
      ~_GEN_416 & (_GEN_420 ? _GEN_985 : _GEN_421 & searcher_is_older_12 & _GEN_986);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_13 =
      l_forwarders_13_0 ? wb_forward_stq_idx_0 : ldq_13_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_987 =
      ~ldq_13_bits_forward_std_val | l_forward_stq_idx_13 != lcam_stq_idx_0
      & (l_forward_stq_idx_13 < lcam_stq_idx_0
         ^ l_forward_stq_idx_13 < ldq_13_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_13_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_988 = _GEN_429 & ~s1_executing_loads_13 & ldq_13_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_29 =
      ~_GEN_427 & (_GEN_431 ? _GEN_987 : _GEN_432 & searcher_is_older_13 & _GEN_988);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    l_forward_stq_idx_14 =
      l_forwarders_14_0 ? wb_forward_stq_idx_0 : ldq_14_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_989 =
      ~ldq_14_bits_forward_std_val | l_forward_stq_idx_14 != lcam_stq_idx_0
      & (l_forward_stq_idx_14 < lcam_stq_idx_0
         ^ l_forward_stq_idx_14 < ldq_14_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_14_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_990 = _GEN_440 & ~s1_executing_loads_14 & ldq_14_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_30 =
      ~_GEN_438 & (_GEN_442 ? _GEN_989 : _GEN_443 & searcher_is_older_14 & _GEN_990);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:72
    _GEN_991 =
      (_GEN_446 | ~_GEN_443 | searcher_is_older_14
       | ~(_GEN_444 & _GEN_445 & (&lcam_ldq_idx_0)))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13
         | ~(_GEN_433 & _GEN_434 & (&lcam_ldq_idx_0)))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12
         | ~(_GEN_422 & _GEN_423 & (&lcam_ldq_idx_0)))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11
         | ~(_GEN_411 & _GEN_412 & (&lcam_ldq_idx_0)))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10
         | ~(_GEN_400 & _GEN_401 & (&lcam_ldq_idx_0)))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9
         | ~(_GEN_389 & _GEN_390 & (&lcam_ldq_idx_0)))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8
         | ~(_GEN_378 & _GEN_379 & (&lcam_ldq_idx_0)))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7
         | ~(_GEN_367 & _GEN_368 & (&lcam_ldq_idx_0)))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6
         | ~(_GEN_356 & _GEN_357 & (&lcam_ldq_idx_0)))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5
         | ~(_GEN_345 & _GEN_346 & (&lcam_ldq_idx_0)))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4
         | ~(_GEN_334 & _GEN_335 & (&lcam_ldq_idx_0)))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3
         | ~(_GEN_323 & _GEN_324 & (&lcam_ldq_idx_0)))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2
         | ~(_GEN_312 & _GEN_313 & (&lcam_ldq_idx_0)))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1
         | ~(_GEN_301 & _GEN_302 & (&lcam_ldq_idx_0)))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & (&lcam_ldq_idx_0))) & s1_executing_loads_15;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:72
    l_forward_stq_idx_15 =
      l_forwarders_15_0 ? wb_forward_stq_idx_0 : ldq_15_bits_forward_stq_idx;	// lsu.scala:210:16, :1067:36, :1075:63, :1077:32
    _GEN_992 =
      ~ldq_15_bits_forward_std_val | l_forward_stq_idx_15 != lcam_stq_idx_0
      & (l_forward_stq_idx_15 < lcam_stq_idx_0
         ^ l_forward_stq_idx_15 < ldq_15_bits_youngest_stq_idx
         ^ lcam_stq_idx_0 < ldq_15_bits_youngest_stq_idx);	// lsu.scala:210:16, :1040:26, :1077:32, :1106:{15,39}, :1107:{31,52}, util.scala:363:{52,64,72,78}
    _GEN_993 = _GEN_451 & ~s1_executing_loads_15 & ldq_15_bits_observed;	// lsu.scala:210:16, :1056:35, :1098:57, :1120:{17,40}
    _temp_bits_WIRE_1_31 =
      ~_GEN_449 & (_GEN_453 ? _GEN_992 : _GEN_454 & searcher_is_older_15 & _GEN_993);	// lsu.scala:1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, util.scala:363:58
    _GEN_994 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & ~(|lcam_ldq_idx_0)))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14
         | ~(_GEN_444 & _GEN_445 & ~(|lcam_ldq_idx_0)))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13
         | ~(_GEN_433 & _GEN_434 & ~(|lcam_ldq_idx_0)))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12
         | ~(_GEN_422 & _GEN_423 & ~(|lcam_ldq_idx_0)))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11
         | ~(_GEN_411 & _GEN_412 & ~(|lcam_ldq_idx_0)))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10
         | ~(_GEN_400 & _GEN_401 & ~(|lcam_ldq_idx_0)))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9
         | ~(_GEN_389 & _GEN_390 & ~(|lcam_ldq_idx_0)))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8
         | ~(_GEN_378 & _GEN_379 & ~(|lcam_ldq_idx_0)))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7
         | ~(_GEN_367 & _GEN_368 & ~(|lcam_ldq_idx_0)))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6
         | ~(_GEN_356 & _GEN_357 & ~(|lcam_ldq_idx_0)))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5
         | ~(_GEN_345 & _GEN_346 & ~(|lcam_ldq_idx_0)))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4
         | ~(_GEN_334 & _GEN_335 & ~(|lcam_ldq_idx_0)))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3
         | ~(_GEN_323 & _GEN_324 & ~(|lcam_ldq_idx_0)))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2
         | ~(_GEN_312 & _GEN_313 & ~(|lcam_ldq_idx_0)))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1
         | ~(_GEN_301 & _GEN_302 & ~(|lcam_ldq_idx_0))) & s1_executing_loads_0;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_995 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_949))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_949))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_949))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_949))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_949))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_949))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_949))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_949))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_949))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_949))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_949))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_949))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_949))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_949))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_949))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_949)) & s1_executing_loads_1;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_996 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_950))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_950))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_950))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_950))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_950))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_950))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_950))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_950))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_950))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_950))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_950))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_950))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_950))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_950))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_950))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_950)) & s1_executing_loads_2;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_997 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_951))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_951))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_951))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_951))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_951))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_951))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_951))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_951))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_951))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_951))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_951))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_951))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_951))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_951))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_951))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_951)) & s1_executing_loads_3;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_998 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_952))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_952))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_952))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_952))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_952))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_952))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_952))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_952))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_952))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_952))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_952))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_952))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_952))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_952))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_952))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_952)) & s1_executing_loads_4;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_999 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_953))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_953))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_953))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_953))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_953))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_953))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_953))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_953))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_953))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_953))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_953))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_953))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_953))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_953))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_953))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_953)) & s1_executing_loads_5;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1000 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_954))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_954))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_954))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_954))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_954))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_954))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_954))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_954))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_954))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_954))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_954))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_954))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_954))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_954))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_954))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_954)) & s1_executing_loads_6;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1001 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_955))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_955))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_955))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_955))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_955))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_955))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_955))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_955))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_955))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_955))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_955))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_955))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_955))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_955))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_955))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_955)) & s1_executing_loads_7;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1002 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_956))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_956))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_956))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_956))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_956))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_956))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_956))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_956))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_956))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_956))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_956))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_956))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_956))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_956))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_956))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_956)) & s1_executing_loads_8;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1003 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_957))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_957))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_957))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_957))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_957))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_957))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_957))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_957))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_957))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_957))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_957))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_957))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_957))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_957))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_957))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_957)) & s1_executing_loads_9;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1004 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_958))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_958))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_958))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_958))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_958))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_958))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_958))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_958))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_958))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_958))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_958))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_958))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_958))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_958))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_958))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_958)) & s1_executing_loads_10;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1005 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_959))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_959))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_959))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_959))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_959))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_959))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_959))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_959))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_959))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_959))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_959))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_959))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_959))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_959))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_959))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_959)) & s1_executing_loads_11;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1006 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_960))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_960))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_960))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_960))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_960))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_960))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_960))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_960))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_960))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_960))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_960))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_960))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_960))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_960))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_960))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_960)) & s1_executing_loads_12;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1007 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_961))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_961))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_961))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_961))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_961))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_961))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_961))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_961))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_961))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_961))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_961))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_961))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_961))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_961))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_961))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_961)) & s1_executing_loads_13;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1008 =
      (_GEN_456 | ~_GEN_454 | searcher_is_older_15
       | ~(~(&lcam_ldq_idx_0) & _GEN_455 & _GEN_962))
      & (_GEN_446 | ~_GEN_443 | searcher_is_older_14 | ~(_GEN_444 & _GEN_445 & _GEN_962))
      & (_GEN_435 | ~_GEN_432 | searcher_is_older_13 | ~(_GEN_433 & _GEN_434 & _GEN_962))
      & (_GEN_424 | ~_GEN_421 | searcher_is_older_12 | ~(_GEN_422 & _GEN_423 & _GEN_962))
      & (_GEN_413 | ~_GEN_410 | searcher_is_older_11 | ~(_GEN_411 & _GEN_412 & _GEN_962))
      & (_GEN_402 | ~_GEN_399 | searcher_is_older_10 | ~(_GEN_400 & _GEN_401 & _GEN_962))
      & (_GEN_391 | ~_GEN_388 | searcher_is_older_9 | ~(_GEN_389 & _GEN_390 & _GEN_962))
      & (_GEN_380 | ~_GEN_377 | searcher_is_older_8 | ~(_GEN_378 & _GEN_379 & _GEN_962))
      & (_GEN_369 | ~_GEN_366 | searcher_is_older_7 | ~(_GEN_367 & _GEN_368 & _GEN_962))
      & (_GEN_358 | ~_GEN_355 | searcher_is_older_6 | ~(_GEN_356 & _GEN_357 & _GEN_962))
      & (_GEN_347 | ~_GEN_344 | searcher_is_older_5 | ~(_GEN_345 & _GEN_346 & _GEN_962))
      & (_GEN_336 | ~_GEN_333 | searcher_is_older_4 | ~(_GEN_334 & _GEN_335 & _GEN_962))
      & (_GEN_325 | ~_GEN_322 | searcher_is_older_3 | ~(_GEN_323 & _GEN_324 & _GEN_962))
      & (_GEN_314 | ~_GEN_311 | searcher_is_older_2 | ~(_GEN_312 & _GEN_313 & _GEN_962))
      & (_GEN_303 | ~_GEN_300 | searcher_is_older_1 | ~(_GEN_301 & _GEN_302 & _GEN_962))
      & (_GEN_292 | ~_GEN_290 | searcher_is_older
         | ~((|lcam_ldq_idx_0) & _GEN_291 & _GEN_962)) & s1_executing_loads_14;	// lsu.scala:1036:26, :1056:35, :1091:36, :1102:37, :1115:47, :1116:37, :1118:34, :1125:{38,47}, :1129:{56,73}, :1130:48, util.scala:363:{58,72}
    _GEN_1010 =
      _GEN_460
        ? (_GEN_1009
             ? (|lcam_ldq_idx_0) & _GEN_994
             : ~(_GEN_464 & ~(|lcam_ldq_idx_0)) & _GEN_994)
        : _GEN_994;	// lsu.scala:1036:26, :1091:36, :1102:37, :1116:37, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1011 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_949 & _GEN_995 : ~(_GEN_464 & _GEN_949) & _GEN_995)
        : _GEN_995;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1012 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_950 & _GEN_996 : ~(_GEN_464 & _GEN_950) & _GEN_996)
        : _GEN_996;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1013 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_951 & _GEN_997 : ~(_GEN_464 & _GEN_951) & _GEN_997)
        : _GEN_997;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1014 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_952 & _GEN_998 : ~(_GEN_464 & _GEN_952) & _GEN_998)
        : _GEN_998;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1015 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_953 & _GEN_999 : ~(_GEN_464 & _GEN_953) & _GEN_999)
        : _GEN_999;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1016 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_954 & _GEN_1000 : ~(_GEN_464 & _GEN_954) & _GEN_1000)
        : _GEN_1000;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1017 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_955 & _GEN_1001 : ~(_GEN_464 & _GEN_955) & _GEN_1001)
        : _GEN_1001;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1018 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_956 & _GEN_1002 : ~(_GEN_464 & _GEN_956) & _GEN_1002)
        : _GEN_1002;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1019 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_957 & _GEN_1003 : ~(_GEN_464 & _GEN_957) & _GEN_1003)
        : _GEN_1003;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1020 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_958 & _GEN_1004 : ~(_GEN_464 & _GEN_958) & _GEN_1004)
        : _GEN_1004;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1021 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_959 & _GEN_1005 : ~(_GEN_464 & _GEN_959) & _GEN_1005)
        : _GEN_1005;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1022 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_960 & _GEN_1006 : ~(_GEN_464 & _GEN_960) & _GEN_1006)
        : _GEN_1006;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1023 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_961 & _GEN_1007 : ~(_GEN_464 & _GEN_961) & _GEN_1007)
        : _GEN_1007;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1024 =
      _GEN_460
        ? (_GEN_1009 ? ~_GEN_962 & _GEN_1008 : ~(_GEN_464 & _GEN_962) & _GEN_1008)
        : _GEN_1008;	// lsu.scala:1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1025 =
      _GEN_460
        ? (_GEN_1009
             ? ~(&lcam_ldq_idx_0) & _GEN_991
             : ~(_GEN_464 & (&lcam_ldq_idx_0)) & _GEN_991)
        : _GEN_991;	// lsu.scala:1036:26, :1091:36, :1102:37, :1116:37, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1027 =
      _GEN_467
        ? (_GEN_1026
             ? (|lcam_ldq_idx_0) & _GEN_1010
             : ~(_GEN_471 & ~(|lcam_ldq_idx_0)) & _GEN_1010)
        : _GEN_1010;	// lsu.scala:1036:26, :1091:36, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1028 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_949 & _GEN_1011 : ~(_GEN_471 & _GEN_949) & _GEN_1011)
        : _GEN_1011;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1029 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_950 & _GEN_1012 : ~(_GEN_471 & _GEN_950) & _GEN_1012)
        : _GEN_1012;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1030 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_951 & _GEN_1013 : ~(_GEN_471 & _GEN_951) & _GEN_1013)
        : _GEN_1013;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1031 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_952 & _GEN_1014 : ~(_GEN_471 & _GEN_952) & _GEN_1014)
        : _GEN_1014;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1032 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_953 & _GEN_1015 : ~(_GEN_471 & _GEN_953) & _GEN_1015)
        : _GEN_1015;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1033 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_954 & _GEN_1016 : ~(_GEN_471 & _GEN_954) & _GEN_1016)
        : _GEN_1016;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1034 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_955 & _GEN_1017 : ~(_GEN_471 & _GEN_955) & _GEN_1017)
        : _GEN_1017;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1035 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_956 & _GEN_1018 : ~(_GEN_471 & _GEN_956) & _GEN_1018)
        : _GEN_1018;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1036 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_957 & _GEN_1019 : ~(_GEN_471 & _GEN_957) & _GEN_1019)
        : _GEN_1019;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1037 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_958 & _GEN_1020 : ~(_GEN_471 & _GEN_958) & _GEN_1020)
        : _GEN_1020;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1038 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_959 & _GEN_1021 : ~(_GEN_471 & _GEN_959) & _GEN_1021)
        : _GEN_1021;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1039 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_960 & _GEN_1022 : ~(_GEN_471 & _GEN_960) & _GEN_1022)
        : _GEN_1022;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1040 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_961 & _GEN_1023 : ~(_GEN_471 & _GEN_961) & _GEN_1023)
        : _GEN_1023;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1041 =
      _GEN_467
        ? (_GEN_1026 ? ~_GEN_962 & _GEN_1024 : ~(_GEN_471 & _GEN_962) & _GEN_1024)
        : _GEN_1024;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1042 =
      _GEN_467
        ? (_GEN_1026
             ? ~(&lcam_ldq_idx_0) & _GEN_1025
             : ~(_GEN_471 & (&lcam_ldq_idx_0)) & _GEN_1025)
        : _GEN_1025;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1044 =
      _GEN_474
        ? (_GEN_1043
             ? (|lcam_ldq_idx_0) & _GEN_1027
             : ~(_GEN_478 & ~(|lcam_ldq_idx_0)) & _GEN_1027)
        : _GEN_1027;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1045 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_949 & _GEN_1028 : ~(_GEN_478 & _GEN_949) & _GEN_1028)
        : _GEN_1028;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1046 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_950 & _GEN_1029 : ~(_GEN_478 & _GEN_950) & _GEN_1029)
        : _GEN_1029;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1047 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_951 & _GEN_1030 : ~(_GEN_478 & _GEN_951) & _GEN_1030)
        : _GEN_1030;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1048 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_952 & _GEN_1031 : ~(_GEN_478 & _GEN_952) & _GEN_1031)
        : _GEN_1031;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1049 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_953 & _GEN_1032 : ~(_GEN_478 & _GEN_953) & _GEN_1032)
        : _GEN_1032;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1050 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_954 & _GEN_1033 : ~(_GEN_478 & _GEN_954) & _GEN_1033)
        : _GEN_1033;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1051 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_955 & _GEN_1034 : ~(_GEN_478 & _GEN_955) & _GEN_1034)
        : _GEN_1034;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1052 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_956 & _GEN_1035 : ~(_GEN_478 & _GEN_956) & _GEN_1035)
        : _GEN_1035;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1053 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_957 & _GEN_1036 : ~(_GEN_478 & _GEN_957) & _GEN_1036)
        : _GEN_1036;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1054 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_958 & _GEN_1037 : ~(_GEN_478 & _GEN_958) & _GEN_1037)
        : _GEN_1037;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1055 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_959 & _GEN_1038 : ~(_GEN_478 & _GEN_959) & _GEN_1038)
        : _GEN_1038;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1056 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_960 & _GEN_1039 : ~(_GEN_478 & _GEN_960) & _GEN_1039)
        : _GEN_1039;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1057 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_961 & _GEN_1040 : ~(_GEN_478 & _GEN_961) & _GEN_1040)
        : _GEN_1040;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1058 =
      _GEN_474
        ? (_GEN_1043 ? ~_GEN_962 & _GEN_1041 : ~(_GEN_478 & _GEN_962) & _GEN_1041)
        : _GEN_1041;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1059 =
      _GEN_474
        ? (_GEN_1043
             ? ~(&lcam_ldq_idx_0) & _GEN_1042
             : ~(_GEN_478 & (&lcam_ldq_idx_0)) & _GEN_1042)
        : _GEN_1042;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1061 =
      _GEN_481
        ? (_GEN_1060
             ? (|lcam_ldq_idx_0) & _GEN_1044
             : ~(_GEN_485 & ~(|lcam_ldq_idx_0)) & _GEN_1044)
        : _GEN_1044;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1062 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_949 & _GEN_1045 : ~(_GEN_485 & _GEN_949) & _GEN_1045)
        : _GEN_1045;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1063 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_950 & _GEN_1046 : ~(_GEN_485 & _GEN_950) & _GEN_1046)
        : _GEN_1046;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1064 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_951 & _GEN_1047 : ~(_GEN_485 & _GEN_951) & _GEN_1047)
        : _GEN_1047;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1065 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_952 & _GEN_1048 : ~(_GEN_485 & _GEN_952) & _GEN_1048)
        : _GEN_1048;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1066 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_953 & _GEN_1049 : ~(_GEN_485 & _GEN_953) & _GEN_1049)
        : _GEN_1049;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1067 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_954 & _GEN_1050 : ~(_GEN_485 & _GEN_954) & _GEN_1050)
        : _GEN_1050;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1068 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_955 & _GEN_1051 : ~(_GEN_485 & _GEN_955) & _GEN_1051)
        : _GEN_1051;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1069 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_956 & _GEN_1052 : ~(_GEN_485 & _GEN_956) & _GEN_1052)
        : _GEN_1052;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1070 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_957 & _GEN_1053 : ~(_GEN_485 & _GEN_957) & _GEN_1053)
        : _GEN_1053;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1071 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_958 & _GEN_1054 : ~(_GEN_485 & _GEN_958) & _GEN_1054)
        : _GEN_1054;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1072 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_959 & _GEN_1055 : ~(_GEN_485 & _GEN_959) & _GEN_1055)
        : _GEN_1055;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1073 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_960 & _GEN_1056 : ~(_GEN_485 & _GEN_960) & _GEN_1056)
        : _GEN_1056;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1074 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_961 & _GEN_1057 : ~(_GEN_485 & _GEN_961) & _GEN_1057)
        : _GEN_1057;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1075 =
      _GEN_481
        ? (_GEN_1060 ? ~_GEN_962 & _GEN_1058 : ~(_GEN_485 & _GEN_962) & _GEN_1058)
        : _GEN_1058;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1076 =
      _GEN_481
        ? (_GEN_1060
             ? ~(&lcam_ldq_idx_0) & _GEN_1059
             : ~(_GEN_485 & (&lcam_ldq_idx_0)) & _GEN_1059)
        : _GEN_1059;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1078 =
      _GEN_488
        ? (_GEN_1077
             ? (|lcam_ldq_idx_0) & _GEN_1061
             : ~(_GEN_492 & ~(|lcam_ldq_idx_0)) & _GEN_1061)
        : _GEN_1061;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1079 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_949 & _GEN_1062 : ~(_GEN_492 & _GEN_949) & _GEN_1062)
        : _GEN_1062;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1080 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_950 & _GEN_1063 : ~(_GEN_492 & _GEN_950) & _GEN_1063)
        : _GEN_1063;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1081 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_951 & _GEN_1064 : ~(_GEN_492 & _GEN_951) & _GEN_1064)
        : _GEN_1064;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1082 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_952 & _GEN_1065 : ~(_GEN_492 & _GEN_952) & _GEN_1065)
        : _GEN_1065;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1083 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_953 & _GEN_1066 : ~(_GEN_492 & _GEN_953) & _GEN_1066)
        : _GEN_1066;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1084 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_954 & _GEN_1067 : ~(_GEN_492 & _GEN_954) & _GEN_1067)
        : _GEN_1067;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1085 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_955 & _GEN_1068 : ~(_GEN_492 & _GEN_955) & _GEN_1068)
        : _GEN_1068;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1086 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_956 & _GEN_1069 : ~(_GEN_492 & _GEN_956) & _GEN_1069)
        : _GEN_1069;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1087 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_957 & _GEN_1070 : ~(_GEN_492 & _GEN_957) & _GEN_1070)
        : _GEN_1070;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1088 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_958 & _GEN_1071 : ~(_GEN_492 & _GEN_958) & _GEN_1071)
        : _GEN_1071;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1089 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_959 & _GEN_1072 : ~(_GEN_492 & _GEN_959) & _GEN_1072)
        : _GEN_1072;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1090 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_960 & _GEN_1073 : ~(_GEN_492 & _GEN_960) & _GEN_1073)
        : _GEN_1073;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1091 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_961 & _GEN_1074 : ~(_GEN_492 & _GEN_961) & _GEN_1074)
        : _GEN_1074;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1092 =
      _GEN_488
        ? (_GEN_1077 ? ~_GEN_962 & _GEN_1075 : ~(_GEN_492 & _GEN_962) & _GEN_1075)
        : _GEN_1075;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1093 =
      _GEN_488
        ? (_GEN_1077
             ? ~(&lcam_ldq_idx_0) & _GEN_1076
             : ~(_GEN_492 & (&lcam_ldq_idx_0)) & _GEN_1076)
        : _GEN_1076;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1095 =
      _GEN_495
        ? (_GEN_1094
             ? (|lcam_ldq_idx_0) & _GEN_1078
             : ~(_GEN_499 & ~(|lcam_ldq_idx_0)) & _GEN_1078)
        : _GEN_1078;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1096 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_949 & _GEN_1079 : ~(_GEN_499 & _GEN_949) & _GEN_1079)
        : _GEN_1079;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1097 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_950 & _GEN_1080 : ~(_GEN_499 & _GEN_950) & _GEN_1080)
        : _GEN_1080;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1098 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_951 & _GEN_1081 : ~(_GEN_499 & _GEN_951) & _GEN_1081)
        : _GEN_1081;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1099 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_952 & _GEN_1082 : ~(_GEN_499 & _GEN_952) & _GEN_1082)
        : _GEN_1082;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1100 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_953 & _GEN_1083 : ~(_GEN_499 & _GEN_953) & _GEN_1083)
        : _GEN_1083;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1101 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_954 & _GEN_1084 : ~(_GEN_499 & _GEN_954) & _GEN_1084)
        : _GEN_1084;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1102 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_955 & _GEN_1085 : ~(_GEN_499 & _GEN_955) & _GEN_1085)
        : _GEN_1085;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1103 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_956 & _GEN_1086 : ~(_GEN_499 & _GEN_956) & _GEN_1086)
        : _GEN_1086;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1104 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_957 & _GEN_1087 : ~(_GEN_499 & _GEN_957) & _GEN_1087)
        : _GEN_1087;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1105 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_958 & _GEN_1088 : ~(_GEN_499 & _GEN_958) & _GEN_1088)
        : _GEN_1088;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1106 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_959 & _GEN_1089 : ~(_GEN_499 & _GEN_959) & _GEN_1089)
        : _GEN_1089;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1107 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_960 & _GEN_1090 : ~(_GEN_499 & _GEN_960) & _GEN_1090)
        : _GEN_1090;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1108 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_961 & _GEN_1091 : ~(_GEN_499 & _GEN_961) & _GEN_1091)
        : _GEN_1091;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1109 =
      _GEN_495
        ? (_GEN_1094 ? ~_GEN_962 & _GEN_1092 : ~(_GEN_499 & _GEN_962) & _GEN_1092)
        : _GEN_1092;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1110 =
      _GEN_495
        ? (_GEN_1094
             ? ~(&lcam_ldq_idx_0) & _GEN_1093
             : ~(_GEN_499 & (&lcam_ldq_idx_0)) & _GEN_1093)
        : _GEN_1093;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1112 =
      _GEN_502
        ? (_GEN_1111
             ? (|lcam_ldq_idx_0) & _GEN_1095
             : ~(_GEN_506 & ~(|lcam_ldq_idx_0)) & _GEN_1095)
        : _GEN_1095;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1113 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_949 & _GEN_1096 : ~(_GEN_506 & _GEN_949) & _GEN_1096)
        : _GEN_1096;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1114 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_950 & _GEN_1097 : ~(_GEN_506 & _GEN_950) & _GEN_1097)
        : _GEN_1097;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1115 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_951 & _GEN_1098 : ~(_GEN_506 & _GEN_951) & _GEN_1098)
        : _GEN_1098;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1116 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_952 & _GEN_1099 : ~(_GEN_506 & _GEN_952) & _GEN_1099)
        : _GEN_1099;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1117 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_953 & _GEN_1100 : ~(_GEN_506 & _GEN_953) & _GEN_1100)
        : _GEN_1100;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1118 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_954 & _GEN_1101 : ~(_GEN_506 & _GEN_954) & _GEN_1101)
        : _GEN_1101;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1119 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_955 & _GEN_1102 : ~(_GEN_506 & _GEN_955) & _GEN_1102)
        : _GEN_1102;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1120 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_956 & _GEN_1103 : ~(_GEN_506 & _GEN_956) & _GEN_1103)
        : _GEN_1103;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1121 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_957 & _GEN_1104 : ~(_GEN_506 & _GEN_957) & _GEN_1104)
        : _GEN_1104;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1122 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_958 & _GEN_1105 : ~(_GEN_506 & _GEN_958) & _GEN_1105)
        : _GEN_1105;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1123 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_959 & _GEN_1106 : ~(_GEN_506 & _GEN_959) & _GEN_1106)
        : _GEN_1106;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1124 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_960 & _GEN_1107 : ~(_GEN_506 & _GEN_960) & _GEN_1107)
        : _GEN_1107;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1125 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_961 & _GEN_1108 : ~(_GEN_506 & _GEN_961) & _GEN_1108)
        : _GEN_1108;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1126 =
      _GEN_502
        ? (_GEN_1111 ? ~_GEN_962 & _GEN_1109 : ~(_GEN_506 & _GEN_962) & _GEN_1109)
        : _GEN_1109;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1127 =
      _GEN_502
        ? (_GEN_1111
             ? ~(&lcam_ldq_idx_0) & _GEN_1110
             : ~(_GEN_506 & (&lcam_ldq_idx_0)) & _GEN_1110)
        : _GEN_1110;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1129 =
      _GEN_509
        ? (_GEN_1128
             ? (|lcam_ldq_idx_0) & _GEN_1112
             : ~(_GEN_513 & ~(|lcam_ldq_idx_0)) & _GEN_1112)
        : _GEN_1112;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1130 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_949 & _GEN_1113 : ~(_GEN_513 & _GEN_949) & _GEN_1113)
        : _GEN_1113;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1131 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_950 & _GEN_1114 : ~(_GEN_513 & _GEN_950) & _GEN_1114)
        : _GEN_1114;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1132 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_951 & _GEN_1115 : ~(_GEN_513 & _GEN_951) & _GEN_1115)
        : _GEN_1115;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1133 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_952 & _GEN_1116 : ~(_GEN_513 & _GEN_952) & _GEN_1116)
        : _GEN_1116;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1134 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_953 & _GEN_1117 : ~(_GEN_513 & _GEN_953) & _GEN_1117)
        : _GEN_1117;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1135 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_954 & _GEN_1118 : ~(_GEN_513 & _GEN_954) & _GEN_1118)
        : _GEN_1118;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1136 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_955 & _GEN_1119 : ~(_GEN_513 & _GEN_955) & _GEN_1119)
        : _GEN_1119;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1137 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_956 & _GEN_1120 : ~(_GEN_513 & _GEN_956) & _GEN_1120)
        : _GEN_1120;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1138 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_957 & _GEN_1121 : ~(_GEN_513 & _GEN_957) & _GEN_1121)
        : _GEN_1121;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1139 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_958 & _GEN_1122 : ~(_GEN_513 & _GEN_958) & _GEN_1122)
        : _GEN_1122;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1140 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_959 & _GEN_1123 : ~(_GEN_513 & _GEN_959) & _GEN_1123)
        : _GEN_1123;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1141 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_960 & _GEN_1124 : ~(_GEN_513 & _GEN_960) & _GEN_1124)
        : _GEN_1124;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1142 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_961 & _GEN_1125 : ~(_GEN_513 & _GEN_961) & _GEN_1125)
        : _GEN_1125;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1143 =
      _GEN_509
        ? (_GEN_1128 ? ~_GEN_962 & _GEN_1126 : ~(_GEN_513 & _GEN_962) & _GEN_1126)
        : _GEN_1126;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1144 =
      _GEN_509
        ? (_GEN_1128
             ? ~(&lcam_ldq_idx_0) & _GEN_1127
             : ~(_GEN_513 & (&lcam_ldq_idx_0)) & _GEN_1127)
        : _GEN_1127;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1146 =
      _GEN_516
        ? (_GEN_1145
             ? (|lcam_ldq_idx_0) & _GEN_1129
             : ~(_GEN_520 & ~(|lcam_ldq_idx_0)) & _GEN_1129)
        : _GEN_1129;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1147 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_949 & _GEN_1130 : ~(_GEN_520 & _GEN_949) & _GEN_1130)
        : _GEN_1130;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1148 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_950 & _GEN_1131 : ~(_GEN_520 & _GEN_950) & _GEN_1131)
        : _GEN_1131;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1149 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_951 & _GEN_1132 : ~(_GEN_520 & _GEN_951) & _GEN_1132)
        : _GEN_1132;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1150 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_952 & _GEN_1133 : ~(_GEN_520 & _GEN_952) & _GEN_1133)
        : _GEN_1133;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1151 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_953 & _GEN_1134 : ~(_GEN_520 & _GEN_953) & _GEN_1134)
        : _GEN_1134;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1152 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_954 & _GEN_1135 : ~(_GEN_520 & _GEN_954) & _GEN_1135)
        : _GEN_1135;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1153 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_955 & _GEN_1136 : ~(_GEN_520 & _GEN_955) & _GEN_1136)
        : _GEN_1136;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1154 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_956 & _GEN_1137 : ~(_GEN_520 & _GEN_956) & _GEN_1137)
        : _GEN_1137;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1155 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_957 & _GEN_1138 : ~(_GEN_520 & _GEN_957) & _GEN_1138)
        : _GEN_1138;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1156 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_958 & _GEN_1139 : ~(_GEN_520 & _GEN_958) & _GEN_1139)
        : _GEN_1139;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1157 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_959 & _GEN_1140 : ~(_GEN_520 & _GEN_959) & _GEN_1140)
        : _GEN_1140;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1158 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_960 & _GEN_1141 : ~(_GEN_520 & _GEN_960) & _GEN_1141)
        : _GEN_1141;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1159 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_961 & _GEN_1142 : ~(_GEN_520 & _GEN_961) & _GEN_1142)
        : _GEN_1142;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1160 =
      _GEN_516
        ? (_GEN_1145 ? ~_GEN_962 & _GEN_1143 : ~(_GEN_520 & _GEN_962) & _GEN_1143)
        : _GEN_1143;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1161 =
      _GEN_516
        ? (_GEN_1145
             ? ~(&lcam_ldq_idx_0) & _GEN_1144
             : ~(_GEN_520 & (&lcam_ldq_idx_0)) & _GEN_1144)
        : _GEN_1144;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1163 =
      _GEN_523
        ? (_GEN_1162
             ? (|lcam_ldq_idx_0) & _GEN_1146
             : ~(_GEN_527 & ~(|lcam_ldq_idx_0)) & _GEN_1146)
        : _GEN_1146;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1164 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_949 & _GEN_1147 : ~(_GEN_527 & _GEN_949) & _GEN_1147)
        : _GEN_1147;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1165 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_950 & _GEN_1148 : ~(_GEN_527 & _GEN_950) & _GEN_1148)
        : _GEN_1148;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1166 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_951 & _GEN_1149 : ~(_GEN_527 & _GEN_951) & _GEN_1149)
        : _GEN_1149;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1167 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_952 & _GEN_1150 : ~(_GEN_527 & _GEN_952) & _GEN_1150)
        : _GEN_1150;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1168 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_953 & _GEN_1151 : ~(_GEN_527 & _GEN_953) & _GEN_1151)
        : _GEN_1151;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1169 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_954 & _GEN_1152 : ~(_GEN_527 & _GEN_954) & _GEN_1152)
        : _GEN_1152;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1170 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_955 & _GEN_1153 : ~(_GEN_527 & _GEN_955) & _GEN_1153)
        : _GEN_1153;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1171 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_956 & _GEN_1154 : ~(_GEN_527 & _GEN_956) & _GEN_1154)
        : _GEN_1154;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1172 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_957 & _GEN_1155 : ~(_GEN_527 & _GEN_957) & _GEN_1155)
        : _GEN_1155;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1173 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_958 & _GEN_1156 : ~(_GEN_527 & _GEN_958) & _GEN_1156)
        : _GEN_1156;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1174 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_959 & _GEN_1157 : ~(_GEN_527 & _GEN_959) & _GEN_1157)
        : _GEN_1157;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1175 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_960 & _GEN_1158 : ~(_GEN_527 & _GEN_960) & _GEN_1158)
        : _GEN_1158;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1176 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_961 & _GEN_1159 : ~(_GEN_527 & _GEN_961) & _GEN_1159)
        : _GEN_1159;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1177 =
      _GEN_523
        ? (_GEN_1162 ? ~_GEN_962 & _GEN_1160 : ~(_GEN_527 & _GEN_962) & _GEN_1160)
        : _GEN_1160;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1178 =
      _GEN_523
        ? (_GEN_1162
             ? ~(&lcam_ldq_idx_0) & _GEN_1161
             : ~(_GEN_527 & (&lcam_ldq_idx_0)) & _GEN_1161)
        : _GEN_1161;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1180 =
      _GEN_530
        ? (_GEN_1179
             ? (|lcam_ldq_idx_0) & _GEN_1163
             : ~(_GEN_534 & ~(|lcam_ldq_idx_0)) & _GEN_1163)
        : _GEN_1163;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1181 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_949 & _GEN_1164 : ~(_GEN_534 & _GEN_949) & _GEN_1164)
        : _GEN_1164;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1182 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_950 & _GEN_1165 : ~(_GEN_534 & _GEN_950) & _GEN_1165)
        : _GEN_1165;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1183 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_951 & _GEN_1166 : ~(_GEN_534 & _GEN_951) & _GEN_1166)
        : _GEN_1166;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1184 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_952 & _GEN_1167 : ~(_GEN_534 & _GEN_952) & _GEN_1167)
        : _GEN_1167;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1185 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_953 & _GEN_1168 : ~(_GEN_534 & _GEN_953) & _GEN_1168)
        : _GEN_1168;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1186 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_954 & _GEN_1169 : ~(_GEN_534 & _GEN_954) & _GEN_1169)
        : _GEN_1169;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1187 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_955 & _GEN_1170 : ~(_GEN_534 & _GEN_955) & _GEN_1170)
        : _GEN_1170;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1188 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_956 & _GEN_1171 : ~(_GEN_534 & _GEN_956) & _GEN_1171)
        : _GEN_1171;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1189 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_957 & _GEN_1172 : ~(_GEN_534 & _GEN_957) & _GEN_1172)
        : _GEN_1172;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1190 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_958 & _GEN_1173 : ~(_GEN_534 & _GEN_958) & _GEN_1173)
        : _GEN_1173;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1191 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_959 & _GEN_1174 : ~(_GEN_534 & _GEN_959) & _GEN_1174)
        : _GEN_1174;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1192 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_960 & _GEN_1175 : ~(_GEN_534 & _GEN_960) & _GEN_1175)
        : _GEN_1175;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1193 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_961 & _GEN_1176 : ~(_GEN_534 & _GEN_961) & _GEN_1176)
        : _GEN_1176;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1194 =
      _GEN_530
        ? (_GEN_1179 ? ~_GEN_962 & _GEN_1177 : ~(_GEN_534 & _GEN_962) & _GEN_1177)
        : _GEN_1177;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1195 =
      _GEN_530
        ? (_GEN_1179
             ? ~(&lcam_ldq_idx_0) & _GEN_1178
             : ~(_GEN_534 & (&lcam_ldq_idx_0)) & _GEN_1178)
        : _GEN_1178;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1197 =
      _GEN_537
        ? (_GEN_1196
             ? (|lcam_ldq_idx_0) & _GEN_1180
             : ~(_GEN_541 & ~(|lcam_ldq_idx_0)) & _GEN_1180)
        : _GEN_1180;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1198 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_949 & _GEN_1181 : ~(_GEN_541 & _GEN_949) & _GEN_1181)
        : _GEN_1181;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1199 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_950 & _GEN_1182 : ~(_GEN_541 & _GEN_950) & _GEN_1182)
        : _GEN_1182;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1200 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_951 & _GEN_1183 : ~(_GEN_541 & _GEN_951) & _GEN_1183)
        : _GEN_1183;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1201 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_952 & _GEN_1184 : ~(_GEN_541 & _GEN_952) & _GEN_1184)
        : _GEN_1184;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1202 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_953 & _GEN_1185 : ~(_GEN_541 & _GEN_953) & _GEN_1185)
        : _GEN_1185;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1203 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_954 & _GEN_1186 : ~(_GEN_541 & _GEN_954) & _GEN_1186)
        : _GEN_1186;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1204 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_955 & _GEN_1187 : ~(_GEN_541 & _GEN_955) & _GEN_1187)
        : _GEN_1187;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1205 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_956 & _GEN_1188 : ~(_GEN_541 & _GEN_956) & _GEN_1188)
        : _GEN_1188;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1206 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_957 & _GEN_1189 : ~(_GEN_541 & _GEN_957) & _GEN_1189)
        : _GEN_1189;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1207 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_958 & _GEN_1190 : ~(_GEN_541 & _GEN_958) & _GEN_1190)
        : _GEN_1190;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1208 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_959 & _GEN_1191 : ~(_GEN_541 & _GEN_959) & _GEN_1191)
        : _GEN_1191;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1209 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_960 & _GEN_1192 : ~(_GEN_541 & _GEN_960) & _GEN_1192)
        : _GEN_1192;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1210 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_961 & _GEN_1193 : ~(_GEN_541 & _GEN_961) & _GEN_1193)
        : _GEN_1193;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1211 =
      _GEN_537
        ? (_GEN_1196 ? ~_GEN_962 & _GEN_1194 : ~(_GEN_541 & _GEN_962) & _GEN_1194)
        : _GEN_1194;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1212 =
      _GEN_537
        ? (_GEN_1196
             ? ~(&lcam_ldq_idx_0) & _GEN_1195
             : ~(_GEN_541 & (&lcam_ldq_idx_0)) & _GEN_1195)
        : _GEN_1195;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1214 =
      _GEN_544
        ? (_GEN_1213
             ? (|lcam_ldq_idx_0) & _GEN_1197
             : ~(_GEN_548 & ~(|lcam_ldq_idx_0)) & _GEN_1197)
        : _GEN_1197;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1215 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_949 & _GEN_1198 : ~(_GEN_548 & _GEN_949) & _GEN_1198)
        : _GEN_1198;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1216 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_950 & _GEN_1199 : ~(_GEN_548 & _GEN_950) & _GEN_1199)
        : _GEN_1199;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1217 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_951 & _GEN_1200 : ~(_GEN_548 & _GEN_951) & _GEN_1200)
        : _GEN_1200;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1218 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_952 & _GEN_1201 : ~(_GEN_548 & _GEN_952) & _GEN_1201)
        : _GEN_1201;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1219 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_953 & _GEN_1202 : ~(_GEN_548 & _GEN_953) & _GEN_1202)
        : _GEN_1202;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1220 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_954 & _GEN_1203 : ~(_GEN_548 & _GEN_954) & _GEN_1203)
        : _GEN_1203;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1221 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_955 & _GEN_1204 : ~(_GEN_548 & _GEN_955) & _GEN_1204)
        : _GEN_1204;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1222 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_956 & _GEN_1205 : ~(_GEN_548 & _GEN_956) & _GEN_1205)
        : _GEN_1205;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1223 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_957 & _GEN_1206 : ~(_GEN_548 & _GEN_957) & _GEN_1206)
        : _GEN_1206;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1224 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_958 & _GEN_1207 : ~(_GEN_548 & _GEN_958) & _GEN_1207)
        : _GEN_1207;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1225 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_959 & _GEN_1208 : ~(_GEN_548 & _GEN_959) & _GEN_1208)
        : _GEN_1208;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1226 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_960 & _GEN_1209 : ~(_GEN_548 & _GEN_960) & _GEN_1209)
        : _GEN_1209;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1227 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_961 & _GEN_1210 : ~(_GEN_548 & _GEN_961) & _GEN_1210)
        : _GEN_1210;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1228 =
      _GEN_544
        ? (_GEN_1213 ? ~_GEN_962 & _GEN_1211 : ~(_GEN_548 & _GEN_962) & _GEN_1211)
        : _GEN_1211;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1229 =
      _GEN_544
        ? (_GEN_1213
             ? ~(&lcam_ldq_idx_0) & _GEN_1212
             : ~(_GEN_548 & (&lcam_ldq_idx_0)) & _GEN_1212)
        : _GEN_1212;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1231 =
      _GEN_551
        ? (_GEN_1230
             ? (|lcam_ldq_idx_0) & _GEN_1214
             : ~(_GEN_555 & ~(|lcam_ldq_idx_0)) & _GEN_1214)
        : _GEN_1214;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1232 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_949 & _GEN_1215 : ~(_GEN_555 & _GEN_949) & _GEN_1215)
        : _GEN_1215;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1233 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_950 & _GEN_1216 : ~(_GEN_555 & _GEN_950) & _GEN_1216)
        : _GEN_1216;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1234 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_951 & _GEN_1217 : ~(_GEN_555 & _GEN_951) & _GEN_1217)
        : _GEN_1217;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1235 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_952 & _GEN_1218 : ~(_GEN_555 & _GEN_952) & _GEN_1218)
        : _GEN_1218;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1236 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_953 & _GEN_1219 : ~(_GEN_555 & _GEN_953) & _GEN_1219)
        : _GEN_1219;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1237 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_954 & _GEN_1220 : ~(_GEN_555 & _GEN_954) & _GEN_1220)
        : _GEN_1220;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1238 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_955 & _GEN_1221 : ~(_GEN_555 & _GEN_955) & _GEN_1221)
        : _GEN_1221;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1239 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_956 & _GEN_1222 : ~(_GEN_555 & _GEN_956) & _GEN_1222)
        : _GEN_1222;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1240 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_957 & _GEN_1223 : ~(_GEN_555 & _GEN_957) & _GEN_1223)
        : _GEN_1223;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1241 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_958 & _GEN_1224 : ~(_GEN_555 & _GEN_958) & _GEN_1224)
        : _GEN_1224;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1242 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_959 & _GEN_1225 : ~(_GEN_555 & _GEN_959) & _GEN_1225)
        : _GEN_1225;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1243 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_960 & _GEN_1226 : ~(_GEN_555 & _GEN_960) & _GEN_1226)
        : _GEN_1226;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1244 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_961 & _GEN_1227 : ~(_GEN_555 & _GEN_961) & _GEN_1227)
        : _GEN_1227;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1245 =
      _GEN_551
        ? (_GEN_1230 ? ~_GEN_962 & _GEN_1228 : ~(_GEN_555 & _GEN_962) & _GEN_1228)
        : _GEN_1228;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1246 =
      _GEN_551
        ? (_GEN_1230
             ? ~(&lcam_ldq_idx_0) & _GEN_1229
             : ~(_GEN_555 & (&lcam_ldq_idx_0)) & _GEN_1229)
        : _GEN_1229;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1248 =
      _GEN_558
        ? (_GEN_1247
             ? (|lcam_ldq_idx_0) & _GEN_1231
             : ~(_GEN_562 & ~(|lcam_ldq_idx_0)) & _GEN_1231)
        : _GEN_1231;	// lsu.scala:1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1249 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_949 & _GEN_1232 : ~(_GEN_562 & _GEN_949) & _GEN_1232)
        : _GEN_1232;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1250 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_950 & _GEN_1233 : ~(_GEN_562 & _GEN_950) & _GEN_1233)
        : _GEN_1233;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1251 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_951 & _GEN_1234 : ~(_GEN_562 & _GEN_951) & _GEN_1234)
        : _GEN_1234;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1252 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_952 & _GEN_1235 : ~(_GEN_562 & _GEN_952) & _GEN_1235)
        : _GEN_1235;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1253 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_953 & _GEN_1236 : ~(_GEN_562 & _GEN_953) & _GEN_1236)
        : _GEN_1236;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1254 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_954 & _GEN_1237 : ~(_GEN_562 & _GEN_954) & _GEN_1237)
        : _GEN_1237;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1255 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_955 & _GEN_1238 : ~(_GEN_562 & _GEN_955) & _GEN_1238)
        : _GEN_1238;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1256 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_956 & _GEN_1239 : ~(_GEN_562 & _GEN_956) & _GEN_1239)
        : _GEN_1239;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1257 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_957 & _GEN_1240 : ~(_GEN_562 & _GEN_957) & _GEN_1240)
        : _GEN_1240;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1258 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_958 & _GEN_1241 : ~(_GEN_562 & _GEN_958) & _GEN_1241)
        : _GEN_1241;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1259 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_959 & _GEN_1242 : ~(_GEN_562 & _GEN_959) & _GEN_1242)
        : _GEN_1242;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1260 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_960 & _GEN_1243 : ~(_GEN_562 & _GEN_960) & _GEN_1243)
        : _GEN_1243;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1261 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_961 & _GEN_1244 : ~(_GEN_562 & _GEN_961) & _GEN_1244)
        : _GEN_1244;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1262 =
      _GEN_558
        ? (_GEN_1247 ? ~_GEN_962 & _GEN_1245 : ~(_GEN_562 & _GEN_962) & _GEN_1245)
        : _GEN_1245;	// lsu.scala:1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    _GEN_1263 =
      _GEN_558
        ? (_GEN_1247
             ? ~(&lcam_ldq_idx_0) & _GEN_1246
             : ~(_GEN_562 & (&lcam_ldq_idx_0)) & _GEN_1246)
        : _GEN_1246;	// lsu.scala:1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46
    mem_forward_valid_0 =
      _GEN_1265[_forwarding_age_logic_0_io_forwarding_idx]
      & (io_core_brupdate_b1_mispredict_mask
         & (do_st_search_0
              ? (_lcam_stq_idx_T
                   ? mem_stq_incoming_e_0_bits_uop_br_mask
                   : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_br_mask : 12'h0)
              : do_ld_search_0
                  ? (fired_load_incoming_REG
                       ? mem_ldq_incoming_e_0_bits_uop_br_mask
                       : fired_load_retry_REG
                           ? mem_ldq_retry_e_bits_uop_br_mask
                           : fired_load_wakeup_REG
                               ? mem_ldq_wakeup_e_bits_uop_br_mask
                               : 12'h0)
                  : 12'h0)) == 12'h0 & ~io_core_exception & ~REG_1;	// lsu.scala:669:22, :894:51, :901:51, :902:51, :904:51, :909:37, :910:37, :911:37, :912:37, :913:37, :915:33, :916:33, :917:33, :919:{33,57}, :921:33, :1014:108, :1016:106, :1029:37, :1030:37, :1178:57, :1187:86, :1189:{53,56,64}, util.scala:118:{51,59}
    _l_idx_T_53 =
      _temp_bits_WIRE_1_25 & _temp_bits_T_18
        ? 5'h9
        : _temp_bits_WIRE_1_26 & _temp_bits_T_20
            ? 5'hA
            : _temp_bits_WIRE_1_27 & _temp_bits_T_22
                ? 5'hB
                : _temp_bits_WIRE_1_28 & _temp_bits_T_24
                    ? 5'hC
                    : _temp_bits_WIRE_1_29 & _temp_bits_T_26
                        ? 5'hD
                        : _temp_bits_WIRE_1_30 & _temp_bits_T_28
                            ? 5'hE
                            : _temp_bits_WIRE_1_31
                                ? 5'hF
                                : _temp_bits_WIRE_1_16
                                    ? 5'h10
                                    : _temp_bits_WIRE_1_17
                                        ? 5'h11
                                        : _temp_bits_WIRE_1_18
                                            ? 5'h12
                                            : _temp_bits_WIRE_1_19
                                                ? 5'h13
                                                : _temp_bits_WIRE_1_20
                                                    ? 5'h14
                                                    : _temp_bits_WIRE_1_21
                                                        ? 5'h15
                                                        : _temp_bits_WIRE_1_22
                                                            ? 5'h16
                                                            : _temp_bits_WIRE_1_23
                                                                ? 5'h17
                                                                : _temp_bits_WIRE_1_24
                                                                    ? 5'h18
                                                                    : _temp_bits_WIRE_1_25
                                                                        ? 5'h19
                                                                        : _temp_bits_WIRE_1_26
                                                                            ? 5'h1A
                                                                            : _temp_bits_WIRE_1_27
                                                                                ? 5'h1B
                                                                                : _temp_bits_WIRE_1_28
                                                                                    ? 5'h1C
                                                                                    : _temp_bits_WIRE_1_29
                                                                                        ? 5'h1D
                                                                                        : {4'hF,
                                                                                           ~_temp_bits_WIRE_1_30};	// Mux.scala:47:69, lsu.scala:305:44, :1091:36, :1102:37, :1229:21, util.scala:351:72
    l_idx =
      _temp_bits_WIRE_1_16 & _temp_bits_T
        ? 4'h0
        : _temp_bits_WIRE_1_17 & _temp_bits_T_2
            ? 4'h1
            : _temp_bits_WIRE_1_18 & _temp_bits_T_4
                ? 4'h2
                : _temp_bits_WIRE_1_19 & _temp_bits_T_6
                    ? 4'h3
                    : _temp_bits_WIRE_1_20 & _temp_bits_T_8
                        ? 4'h4
                        : _temp_bits_WIRE_1_21 & _temp_bits_T_10
                            ? 4'h5
                            : _temp_bits_WIRE_1_22 & _temp_bits_T_12
                                ? 4'h6
                                : _temp_bits_WIRE_1_23 & ~(ldq_head[3])
                                    ? 4'h7
                                    : _temp_bits_WIRE_1_24 & _temp_bits_T_16
                                        ? 4'h8
                                        : _l_idx_T_53[3:0];	// Mux.scala:47:69, lsu.scala:215:29, :305:44, :1091:36, :1102:37, :1229:21, util.scala:351:72
    ld_xcpt_valid =
      _temp_bits_WIRE_1_16 | _temp_bits_WIRE_1_17 | _temp_bits_WIRE_1_18
      | _temp_bits_WIRE_1_19 | _temp_bits_WIRE_1_20 | _temp_bits_WIRE_1_21
      | _temp_bits_WIRE_1_22 | _temp_bits_WIRE_1_23 | _temp_bits_WIRE_1_24
      | _temp_bits_WIRE_1_25 | _temp_bits_WIRE_1_26 | _temp_bits_WIRE_1_27
      | _temp_bits_WIRE_1_28 | _temp_bits_WIRE_1_29 | _temp_bits_WIRE_1_30
      | _temp_bits_WIRE_1_31;	// lsu.scala:1091:36, :1102:37, :1238:44
    use_mem_xcpt =
      mem_xcpt_valids_0
      & (mem_xcpt_uops_0_rob_idx < _GEN_140[l_idx]
         ^ mem_xcpt_uops_0_rob_idx < io_core_rob_head_idx
         ^ _GEN_140[l_idx] < io_core_rob_head_idx) | ~ld_xcpt_valid;	// Mux.scala:47:69, lsu.scala:465:79, :667:32, :671:32, :1238:44, :1241:{38,115,118}, util.scala:363:{52,64,72,78}
    xcpt_uop_br_mask = use_mem_xcpt ? mem_xcpt_uops_0_br_mask : _GEN_102[l_idx];	// Mux.scala:47:69, lsu.scala:264:49, :671:32, :1241:115, :1243:21, util.scala:363:52
    _GEN_1267 = _GEN_591 & _GEN_1266 & ~(|wb_forward_ldq_idx_0);	// lsu.scala:1065:36, :1075:88, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1268 = _GEN_590 | ~_GEN_1267;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1269 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h1;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1270 = _GEN_590 | ~_GEN_1269;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1271 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h2;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1272 = _GEN_590 | ~_GEN_1271;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1273 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h3;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1274 = _GEN_590 | ~_GEN_1273;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1275 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h4;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1276 = _GEN_590 | ~_GEN_1275;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1277 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h5;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1278 = _GEN_590 | ~_GEN_1277;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1279 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h6;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1280 = _GEN_590 | ~_GEN_1279;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1281 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h7;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1282 = _GEN_590 | ~_GEN_1281;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1283 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h8;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1284 = _GEN_590 | ~_GEN_1283;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1285 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'h9;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1286 = _GEN_590 | ~_GEN_1285;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1287 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'hA;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1288 = _GEN_590 | ~_GEN_1287;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1289 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'hB;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1290 = _GEN_590 | ~_GEN_1289;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1291 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'hC;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1292 = _GEN_590 | ~_GEN_1291;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1293 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'hD;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1294 = _GEN_590 | ~_GEN_1293;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1295 = _GEN_591 & _GEN_1266 & wb_forward_ldq_idx_0 == 4'hE;	// lsu.scala:305:44, :1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1296 = _GEN_590 | ~_GEN_1295;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1297 = _GEN_591 & _GEN_1266 & (&wb_forward_ldq_idx_0);	// lsu.scala:1065:36, :1306:5, :1347:38, :1348:5, :1369:{24,33}, :1370:35
    _GEN_1298 = _GEN_590 | ~_GEN_1297;	// lsu.scala:1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35
    _GEN_1299 = stq_0_valid & (|_GEN_605);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1300 = stq_1_valid & (|_GEN_606);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1301 = stq_2_valid & (|_GEN_607);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1302 = stq_3_valid & (|_GEN_608);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1303 = stq_4_valid & (|_GEN_609);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1304 = stq_5_valid & (|_GEN_610);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1305 = stq_6_valid & (|_GEN_611);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1306 = stq_7_valid & (|_GEN_612);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1307 = stq_8_valid & (|_GEN_613);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1308 = stq_9_valid & (|_GEN_614);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1309 = stq_10_valid & (|_GEN_615);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1310 = stq_11_valid & (|_GEN_616);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1311 = stq_12_valid & (|_GEN_617);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1312 = stq_13_valid & (|_GEN_618);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1313 = stq_14_valid & (|_GEN_619);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1314 = stq_15_valid & (|_GEN_620);	// lsu.scala:211:16, :304:5, :1404:5, :1408:7, :1409:32, util.scala:118:{51,59}
    _GEN_1315 =
      ldq_0_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_0_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1316 =
      ldq_1_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_1_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1317 =
      ldq_2_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_2_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1318 =
      ldq_3_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_3_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1319 =
      ldq_4_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_4_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1320 =
      ldq_5_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_5_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1321 =
      ldq_6_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_6_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1322 =
      ldq_7_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_7_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1323 =
      ldq_8_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_8_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1324 =
      ldq_9_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_9_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1325 =
      ldq_10_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_10_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1326 =
      ldq_11_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_11_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1327 =
      ldq_12_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_12_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1328 =
      ldq_13_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_13_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1329 =
      ldq_14_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_14_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1330 =
      ldq_15_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_15_bits_uop_br_mask));	// lsu.scala:210:16, :304:5, :1424:5, :1427:7, :1428:32, util.scala:118:{51,59}
    _GEN_1362 = _GEN_1331 | _GEN_1315;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1364 = _GEN_1333 | _GEN_1316;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1365 = _GEN_1335 | _GEN_1317;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1366 = _GEN_1337 | _GEN_1318;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1367 = _GEN_1339 | _GEN_1319;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1368 = _GEN_1341 | _GEN_1320;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1369 = _GEN_1343 | _GEN_1321;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1370 = _GEN_1345 | _GEN_1322;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1371 = _GEN_1347 | _GEN_1323;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1372 = _GEN_1349 | _GEN_1324;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1373 = _GEN_1351 | _GEN_1325;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1374 = _GEN_1353 | _GEN_1326;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1375 = _GEN_1355 | _GEN_1327;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1376 = _GEN_1357 | _GEN_1328;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1377 = _GEN_1359 | _GEN_1329;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1456:31, :1462:38
    _GEN_1378 = (&idx) | _GEN_1330;	// lsu.scala:304:5, :1424:5, :1427:7, :1428:32, :1453:18, :1456:31, :1462:38
    _GEN_1426 = stq_head == 4'h0;	// lsu.scala:217:29, :1506:35
    _GEN_1427 = _GEN_1426 | _GEN_1299;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1428 = stq_head == 4'h1;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1429 = _GEN_1428 | _GEN_1300;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1430 = stq_head == 4'h2;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1431 = _GEN_1430 | _GEN_1301;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1432 = stq_head == 4'h3;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1433 = _GEN_1432 | _GEN_1302;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1434 = stq_head == 4'h4;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1435 = _GEN_1434 | _GEN_1303;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1436 = stq_head == 4'h5;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1437 = _GEN_1436 | _GEN_1304;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1438 = stq_head == 4'h6;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1439 = _GEN_1438 | _GEN_1305;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1440 = stq_head == 4'h7;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1441 = _GEN_1440 | _GEN_1306;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1442 = stq_head == 4'h8;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1443 = _GEN_1442 | _GEN_1307;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1444 = stq_head == 4'h9;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1445 = _GEN_1444 | _GEN_1308;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1446 = stq_head == 4'hA;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1447 = _GEN_1446 | _GEN_1309;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1448 = stq_head == 4'hB;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1449 = _GEN_1448 | _GEN_1310;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1450 = stq_head == 4'hC;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1451 = _GEN_1450 | _GEN_1311;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1452 = stq_head == 4'hD;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1453 = _GEN_1452 | _GEN_1312;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1454 = stq_head == 4'hE;	// lsu.scala:217:29, :305:44, :1506:35
    _GEN_1455 = _GEN_1454 | _GEN_1313;	// lsu.scala:304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1456 = (&stq_head) | _GEN_1314;	// lsu.scala:217:29, :304:5, :1404:5, :1408:7, :1409:32, :1506:35
    _GEN_1457 = clear_store & _GEN_1426;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1458 = clear_store & _GEN_1428;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1459 = clear_store & _GEN_1430;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1460 = clear_store & _GEN_1432;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1461 = clear_store & _GEN_1434;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1462 = clear_store & _GEN_1436;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1463 = clear_store & _GEN_1438;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1464 = clear_store & _GEN_1440;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1465 = clear_store & _GEN_1442;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1466 = clear_store & _GEN_1444;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1467 = clear_store & _GEN_1446;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1468 = clear_store & _GEN_1448;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1469 = clear_store & _GEN_1450;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1470 = clear_store & _GEN_1452;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1471 = clear_store & _GEN_1454;	// lsu.scala:1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1472 = clear_store & (&stq_head);	// lsu.scala:217:29, :1306:5, :1495:3, :1500:17, :1505:3, :1506:35, :1509:35
    _GEN_1473 = ~(|hella_state) & io_hellacache_req_valid;	// Decoupled.scala:40:37, lsu.scala:242:38, :593:24, :1527:21
    _GEN_1474 = ~(|hella_state) & _GEN_1473;	// Decoupled.scala:40:37, lsu.scala:242:38, :243:34, :593:24, :1527:{21,34}, :1529:37, :1530:19
    _GEN_1475 = (|hella_state) & _GEN_1;	// lsu.scala:242:38, :244:34, :593:24, :803:26, :1527:34, :1533:38
    _GEN_1476 = reset | io_core_exception;	// lsu.scala:1596:22
    _GEN_1477 = _GEN_1476 & reset;	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1603:16
    _GEN_1478 = ~stq_0_bits_committed & ~stq_0_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1479 = _GEN_1476 & (reset | _GEN_1478);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1480 = ~stq_1_bits_committed & ~stq_1_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1481 = _GEN_1476 & (reset | _GEN_1480);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1482 = ~stq_2_bits_committed & ~stq_2_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1483 = _GEN_1476 & (reset | _GEN_1482);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1484 = ~stq_3_bits_committed & ~stq_3_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1485 = _GEN_1476 & (reset | _GEN_1484);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1486 = ~stq_4_bits_committed & ~stq_4_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1487 = _GEN_1476 & (reset | _GEN_1486);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1488 = ~stq_5_bits_committed & ~stq_5_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1489 = _GEN_1476 & (reset | _GEN_1488);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1490 = ~stq_6_bits_committed & ~stq_6_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1491 = _GEN_1476 & (reset | _GEN_1490);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1492 = ~stq_7_bits_committed & ~stq_7_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1493 = _GEN_1476 & (reset | _GEN_1492);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1494 = ~stq_8_bits_committed & ~stq_8_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1495 = _GEN_1476 & (reset | _GEN_1494);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1496 = ~stq_9_bits_committed & ~stq_9_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1497 = _GEN_1476 & (reset | _GEN_1496);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1498 = ~stq_10_bits_committed & ~stq_10_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1499 = _GEN_1476 & (reset | _GEN_1498);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1500 = ~stq_11_bits_committed & ~stq_11_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1501 = _GEN_1476 & (reset | _GEN_1500);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1502 = ~stq_12_bits_committed & ~stq_12_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1503 = _GEN_1476 & (reset | _GEN_1502);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1504 = ~stq_13_bits_committed & ~stq_13_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1505 = _GEN_1476 & (reset | _GEN_1504);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1506 = ~stq_14_bits_committed & ~stq_14_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1507 = _GEN_1476 & (reset | _GEN_1506);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    _GEN_1508 = ~stq_15_bits_committed & ~stq_15_bits_succeeded;	// lsu.scala:211:16, :1622:{15,38,41}
    _GEN_1509 = _GEN_1476 & (reset | _GEN_1508);	// lsu.scala:1505:3, :1596:22, :1597:3, :1602:5, :1610:32, :1622:38, :1623:9, :1624:34
    ldq_0_valid <=
      ~_GEN_1476 & _GEN_1410
      & (_GEN_1363 ? ~_GEN_1315 & _GEN_694 : ~_GEN_1362 & _GEN_694);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_739) begin	// lsu.scala:304:5, :306:44
      ldq_0_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_0_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_0_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_0_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_0_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_0_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_643) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_0_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_0_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_0_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_0_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_0_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_0_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_0_valid)	// lsu.scala:210:16
      ldq_0_bits_uop_br_mask <=
        ldq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_739)	// lsu.scala:304:5, :306:44
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_643)	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_851) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_0_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_0_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_0_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_0_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_0_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_0_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_0_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_0_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_0_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_0_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_0_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_739)	// lsu.scala:304:5, :306:44
      ldq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_643)	// lsu.scala:210:16, :304:5, :305:44
      ldq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_755)	// lsu.scala:210:16, :304:5, :306:44
      ldq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_0_bits_uop_ppred_busy <= ~_GEN_755 & ldq_0_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_0_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h0
      | (_GEN_739
           ? io_core_dis_uops_1_bits_exception
           : _GEN_643 ? io_core_dis_uops_0_bits_exception : ldq_0_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_0_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1410
      & (_GEN_1363 ? ~_GEN_1315 & _GEN_852 : ~_GEN_1362 & _GEN_852);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_0_bits_executed <=
      ~_GEN_1476 & _GEN_1410 & _GEN_1379
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_573))
      & ((_GEN_565
            ? (_GEN_1264
                 ? (|lcam_ldq_idx_0) & _GEN_1248
                 : ~(_GEN_569 & ~(|lcam_ldq_idx_0)) & _GEN_1248)
            : _GEN_1248)
         | (dis_ld_val_1
              ? ~_GEN_693 & ldq_0_bits_executed
              : ~_GEN_643 & ldq_0_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1036:26, :1125:38, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_0_bits_succeeded <=
      _GEN_1410 & _GEN_1379
      & (_GEN_1268
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h0
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_693 & ldq_0_bits_succeeded
                    : ~_GEN_643 & ldq_0_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_0_bits_order_fail <=
      _GEN_1410 & _GEN_1379
      & (_GEN_284
           ? _GEN_771
           : _GEN_289
               ? _GEN_947 | _GEN_771
               : _GEN_290 & searcher_is_older & _GEN_948 | _GEN_771);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_0_bits_observed <=
      _GEN_284
      | (dis_ld_val_1
           ? ~_GEN_693 & ldq_0_bits_observed
           : ~_GEN_643 & ldq_0_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_0_bits_forward_std_val <=
      _GEN_1410 & _GEN_1379
      & (~_GEN_590 & _GEN_1267
         | (dis_ld_val_1
              ? ~_GEN_693 & ldq_0_bits_forward_std_val
              : ~_GEN_643 & ldq_0_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1268) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_0_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_1_valid <=
      ~_GEN_1476 & _GEN_1411
      & (_GEN_1363 ? ~_GEN_1316 & _GEN_697 : ~_GEN_1364 & _GEN_697);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_740) begin	// lsu.scala:304:5, :306:44
      ldq_1_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_1_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_1_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_1_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_1_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_1_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_644) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_1_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_1_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_1_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_1_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_1_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_1_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_1_valid)	// lsu.scala:210:16
      ldq_1_bits_uop_br_mask <=
        ldq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_740)	// lsu.scala:304:5, :306:44
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_644)	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_853) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_1_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_1_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_1_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_1_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_1_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_1_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_1_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_1_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_1_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_1_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_1_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_740)	// lsu.scala:304:5, :306:44
      ldq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_644)	// lsu.scala:210:16, :304:5, :305:44
      ldq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_756)	// lsu.scala:210:16, :304:5, :306:44
      ldq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_1_bits_uop_ppred_busy <= ~_GEN_756 & ldq_1_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_1_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h1
      | (_GEN_740
           ? io_core_dis_uops_1_bits_exception
           : _GEN_644 ? io_core_dis_uops_0_bits_exception : ldq_1_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_1_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1411
      & (_GEN_1363 ? ~_GEN_1316 & _GEN_854 : ~_GEN_1364 & _GEN_854);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_1_bits_executed <=
      ~_GEN_1476 & _GEN_1411 & _GEN_1380
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_574))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_949 & _GEN_1249 : ~(_GEN_569 & _GEN_949) & _GEN_1249)
            : _GEN_1249)
         | (dis_ld_val_1
              ? ~_GEN_696 & ldq_1_bits_executed
              : ~_GEN_644 & ldq_1_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_1_bits_succeeded <=
      _GEN_1411 & _GEN_1380
      & (_GEN_1270
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h1
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_696 & ldq_1_bits_succeeded
                    : ~_GEN_644 & ldq_1_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_1_bits_order_fail <=
      _GEN_1411 & _GEN_1380
      & (_GEN_295
           ? _GEN_772
           : _GEN_299
               ? _GEN_963 | _GEN_772
               : _GEN_300 & searcher_is_older_1 & _GEN_964 | _GEN_772);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_1_bits_observed <=
      _GEN_295
      | (dis_ld_val_1
           ? ~_GEN_696 & ldq_1_bits_observed
           : ~_GEN_644 & ldq_1_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_1_bits_forward_std_val <=
      _GEN_1411 & _GEN_1380
      & (~_GEN_590 & _GEN_1269
         | (dis_ld_val_1
              ? ~_GEN_696 & ldq_1_bits_forward_std_val
              : ~_GEN_644 & ldq_1_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1270) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_1_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_2_valid <=
      ~_GEN_1476 & _GEN_1412
      & (_GEN_1363 ? ~_GEN_1317 & _GEN_700 : ~_GEN_1365 & _GEN_700);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_741) begin	// lsu.scala:304:5, :306:44
      ldq_2_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_2_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_2_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_2_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_2_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_2_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_645) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_2_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_2_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_2_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_2_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_2_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_2_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_2_valid)	// lsu.scala:210:16
      ldq_2_bits_uop_br_mask <=
        ldq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_741)	// lsu.scala:304:5, :306:44
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_645)	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_855) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_2_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_2_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_2_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_2_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_2_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_2_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_2_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_2_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_2_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_2_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_2_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_741)	// lsu.scala:304:5, :306:44
      ldq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_645)	// lsu.scala:210:16, :304:5, :305:44
      ldq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_757)	// lsu.scala:210:16, :304:5, :306:44
      ldq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_2_bits_uop_ppred_busy <= ~_GEN_757 & ldq_2_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_2_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h2
      | (_GEN_741
           ? io_core_dis_uops_1_bits_exception
           : _GEN_645 ? io_core_dis_uops_0_bits_exception : ldq_2_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_2_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1412
      & (_GEN_1363 ? ~_GEN_1317 & _GEN_856 : ~_GEN_1365 & _GEN_856);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_2_bits_executed <=
      ~_GEN_1476 & _GEN_1412 & _GEN_1381
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_575))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_950 & _GEN_1250 : ~(_GEN_569 & _GEN_950) & _GEN_1250)
            : _GEN_1250)
         | (dis_ld_val_1
              ? ~_GEN_699 & ldq_2_bits_executed
              : ~_GEN_645 & ldq_2_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_2_bits_succeeded <=
      _GEN_1412 & _GEN_1381
      & (_GEN_1272
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h2
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_699 & ldq_2_bits_succeeded
                    : ~_GEN_645 & ldq_2_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_2_bits_order_fail <=
      _GEN_1412 & _GEN_1381
      & (_GEN_306
           ? _GEN_773
           : _GEN_310
               ? _GEN_965 | _GEN_773
               : _GEN_311 & searcher_is_older_2 & _GEN_966 | _GEN_773);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_2_bits_observed <=
      _GEN_306
      | (dis_ld_val_1
           ? ~_GEN_699 & ldq_2_bits_observed
           : ~_GEN_645 & ldq_2_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_2_bits_forward_std_val <=
      _GEN_1412 & _GEN_1381
      & (~_GEN_590 & _GEN_1271
         | (dis_ld_val_1
              ? ~_GEN_699 & ldq_2_bits_forward_std_val
              : ~_GEN_645 & ldq_2_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1272) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_2_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_3_valid <=
      ~_GEN_1476 & _GEN_1413
      & (_GEN_1363 ? ~_GEN_1318 & _GEN_703 : ~_GEN_1366 & _GEN_703);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_742) begin	// lsu.scala:304:5, :306:44
      ldq_3_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_3_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_3_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_3_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_3_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_3_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_646) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_3_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_3_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_3_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_3_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_3_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_3_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_3_valid)	// lsu.scala:210:16
      ldq_3_bits_uop_br_mask <=
        ldq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_742)	// lsu.scala:304:5, :306:44
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_646)	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_857) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_3_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_3_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_3_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_3_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_3_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_3_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_3_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_3_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_3_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_3_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_3_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_742)	// lsu.scala:304:5, :306:44
      ldq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_646)	// lsu.scala:210:16, :304:5, :305:44
      ldq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_758)	// lsu.scala:210:16, :304:5, :306:44
      ldq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_3_bits_uop_ppred_busy <= ~_GEN_758 & ldq_3_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_3_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h3
      | (_GEN_742
           ? io_core_dis_uops_1_bits_exception
           : _GEN_646 ? io_core_dis_uops_0_bits_exception : ldq_3_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_3_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1413
      & (_GEN_1363 ? ~_GEN_1318 & _GEN_858 : ~_GEN_1366 & _GEN_858);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_3_bits_executed <=
      ~_GEN_1476 & _GEN_1413 & _GEN_1382
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_576))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_951 & _GEN_1251 : ~(_GEN_569 & _GEN_951) & _GEN_1251)
            : _GEN_1251)
         | (dis_ld_val_1
              ? ~_GEN_702 & ldq_3_bits_executed
              : ~_GEN_646 & ldq_3_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_3_bits_succeeded <=
      _GEN_1413 & _GEN_1382
      & (_GEN_1274
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h3
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_702 & ldq_3_bits_succeeded
                    : ~_GEN_646 & ldq_3_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_3_bits_order_fail <=
      _GEN_1413 & _GEN_1382
      & (_GEN_317
           ? _GEN_774
           : _GEN_321
               ? _GEN_967 | _GEN_774
               : _GEN_322 & searcher_is_older_3 & _GEN_968 | _GEN_774);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_3_bits_observed <=
      _GEN_317
      | (dis_ld_val_1
           ? ~_GEN_702 & ldq_3_bits_observed
           : ~_GEN_646 & ldq_3_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_3_bits_forward_std_val <=
      _GEN_1413 & _GEN_1382
      & (~_GEN_590 & _GEN_1273
         | (dis_ld_val_1
              ? ~_GEN_702 & ldq_3_bits_forward_std_val
              : ~_GEN_646 & ldq_3_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1274) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_3_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_4_valid <=
      ~_GEN_1476 & _GEN_1414
      & (_GEN_1363 ? ~_GEN_1319 & _GEN_706 : ~_GEN_1367 & _GEN_706);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_743) begin	// lsu.scala:304:5, :306:44
      ldq_4_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_4_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_4_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_4_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_4_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_4_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_647) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_4_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_4_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_4_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_4_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_4_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_4_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_4_valid)	// lsu.scala:210:16
      ldq_4_bits_uop_br_mask <=
        ldq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_743)	// lsu.scala:304:5, :306:44
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_647)	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_859) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_4_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_4_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_4_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_4_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_4_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_4_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_4_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_4_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_4_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_4_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_4_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_743)	// lsu.scala:304:5, :306:44
      ldq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_647)	// lsu.scala:210:16, :304:5, :305:44
      ldq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_759)	// lsu.scala:210:16, :304:5, :306:44
      ldq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_4_bits_uop_ppred_busy <= ~_GEN_759 & ldq_4_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_4_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h4
      | (_GEN_743
           ? io_core_dis_uops_1_bits_exception
           : _GEN_647 ? io_core_dis_uops_0_bits_exception : ldq_4_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_4_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1414
      & (_GEN_1363 ? ~_GEN_1319 & _GEN_860 : ~_GEN_1367 & _GEN_860);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_4_bits_executed <=
      ~_GEN_1476 & _GEN_1414 & _GEN_1383
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_577))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_952 & _GEN_1252 : ~(_GEN_569 & _GEN_952) & _GEN_1252)
            : _GEN_1252)
         | (dis_ld_val_1
              ? ~_GEN_705 & ldq_4_bits_executed
              : ~_GEN_647 & ldq_4_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_4_bits_succeeded <=
      _GEN_1414 & _GEN_1383
      & (_GEN_1276
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h4
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_705 & ldq_4_bits_succeeded
                    : ~_GEN_647 & ldq_4_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_4_bits_order_fail <=
      _GEN_1414 & _GEN_1383
      & (_GEN_328
           ? _GEN_775
           : _GEN_332
               ? _GEN_969 | _GEN_775
               : _GEN_333 & searcher_is_older_4 & _GEN_970 | _GEN_775);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_4_bits_observed <=
      _GEN_328
      | (dis_ld_val_1
           ? ~_GEN_705 & ldq_4_bits_observed
           : ~_GEN_647 & ldq_4_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_4_bits_forward_std_val <=
      _GEN_1414 & _GEN_1383
      & (~_GEN_590 & _GEN_1275
         | (dis_ld_val_1
              ? ~_GEN_705 & ldq_4_bits_forward_std_val
              : ~_GEN_647 & ldq_4_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1276) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_4_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_5_valid <=
      ~_GEN_1476 & _GEN_1415
      & (_GEN_1363 ? ~_GEN_1320 & _GEN_709 : ~_GEN_1368 & _GEN_709);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_744) begin	// lsu.scala:304:5, :306:44
      ldq_5_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_5_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_5_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_5_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_5_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_5_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_648) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_5_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_5_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_5_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_5_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_5_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_5_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_5_valid)	// lsu.scala:210:16
      ldq_5_bits_uop_br_mask <=
        ldq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_744)	// lsu.scala:304:5, :306:44
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_648)	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_861) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_5_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_5_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_5_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_5_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_5_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_5_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_5_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_5_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_5_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_5_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_5_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_744)	// lsu.scala:304:5, :306:44
      ldq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_648)	// lsu.scala:210:16, :304:5, :305:44
      ldq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_760)	// lsu.scala:210:16, :304:5, :306:44
      ldq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_5_bits_uop_ppred_busy <= ~_GEN_760 & ldq_5_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_5_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h5
      | (_GEN_744
           ? io_core_dis_uops_1_bits_exception
           : _GEN_648 ? io_core_dis_uops_0_bits_exception : ldq_5_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_5_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1415
      & (_GEN_1363 ? ~_GEN_1320 & _GEN_862 : ~_GEN_1368 & _GEN_862);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_5_bits_executed <=
      ~_GEN_1476 & _GEN_1415 & _GEN_1384
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_578))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_953 & _GEN_1253 : ~(_GEN_569 & _GEN_953) & _GEN_1253)
            : _GEN_1253)
         | (dis_ld_val_1
              ? ~_GEN_708 & ldq_5_bits_executed
              : ~_GEN_648 & ldq_5_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_5_bits_succeeded <=
      _GEN_1415 & _GEN_1384
      & (_GEN_1278
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h5
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_708 & ldq_5_bits_succeeded
                    : ~_GEN_648 & ldq_5_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_5_bits_order_fail <=
      _GEN_1415 & _GEN_1384
      & (_GEN_339
           ? _GEN_776
           : _GEN_343
               ? _GEN_971 | _GEN_776
               : _GEN_344 & searcher_is_older_5 & _GEN_972 | _GEN_776);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_5_bits_observed <=
      _GEN_339
      | (dis_ld_val_1
           ? ~_GEN_708 & ldq_5_bits_observed
           : ~_GEN_648 & ldq_5_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_5_bits_forward_std_val <=
      _GEN_1415 & _GEN_1384
      & (~_GEN_590 & _GEN_1277
         | (dis_ld_val_1
              ? ~_GEN_708 & ldq_5_bits_forward_std_val
              : ~_GEN_648 & ldq_5_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1278) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_5_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_6_valid <=
      ~_GEN_1476 & _GEN_1416
      & (_GEN_1363 ? ~_GEN_1321 & _GEN_712 : ~_GEN_1369 & _GEN_712);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_745) begin	// lsu.scala:304:5, :306:44
      ldq_6_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_6_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_6_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_6_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_6_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_6_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_649) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_6_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_6_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_6_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_6_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_6_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_6_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_6_valid)	// lsu.scala:210:16
      ldq_6_bits_uop_br_mask <=
        ldq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_745)	// lsu.scala:304:5, :306:44
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_649)	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_863) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_6_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_6_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_6_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_6_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_6_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_6_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_6_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_6_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_6_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_6_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_6_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_745)	// lsu.scala:304:5, :306:44
      ldq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_649)	// lsu.scala:210:16, :304:5, :305:44
      ldq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_761)	// lsu.scala:210:16, :304:5, :306:44
      ldq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_6_bits_uop_ppred_busy <= ~_GEN_761 & ldq_6_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_6_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h6
      | (_GEN_745
           ? io_core_dis_uops_1_bits_exception
           : _GEN_649 ? io_core_dis_uops_0_bits_exception : ldq_6_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_6_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1416
      & (_GEN_1363 ? ~_GEN_1321 & _GEN_864 : ~_GEN_1369 & _GEN_864);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_6_bits_executed <=
      ~_GEN_1476 & _GEN_1416 & _GEN_1385
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_579))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_954 & _GEN_1254 : ~(_GEN_569 & _GEN_954) & _GEN_1254)
            : _GEN_1254)
         | (dis_ld_val_1
              ? ~_GEN_711 & ldq_6_bits_executed
              : ~_GEN_649 & ldq_6_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_6_bits_succeeded <=
      _GEN_1416 & _GEN_1385
      & (_GEN_1280
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h6
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_711 & ldq_6_bits_succeeded
                    : ~_GEN_649 & ldq_6_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_6_bits_order_fail <=
      _GEN_1416 & _GEN_1385
      & (_GEN_350
           ? _GEN_777
           : _GEN_354
               ? _GEN_973 | _GEN_777
               : _GEN_355 & searcher_is_older_6 & _GEN_974 | _GEN_777);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_6_bits_observed <=
      _GEN_350
      | (dis_ld_val_1
           ? ~_GEN_711 & ldq_6_bits_observed
           : ~_GEN_649 & ldq_6_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_6_bits_forward_std_val <=
      _GEN_1416 & _GEN_1385
      & (~_GEN_590 & _GEN_1279
         | (dis_ld_val_1
              ? ~_GEN_711 & ldq_6_bits_forward_std_val
              : ~_GEN_649 & ldq_6_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1280) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_6_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_7_valid <=
      ~_GEN_1476 & _GEN_1417
      & (_GEN_1363 ? ~_GEN_1322 & _GEN_715 : ~_GEN_1370 & _GEN_715);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_746) begin	// lsu.scala:304:5, :306:44
      ldq_7_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_7_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_7_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_7_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_7_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_7_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_650) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_7_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_7_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_7_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_7_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_7_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_7_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_7_valid)	// lsu.scala:210:16
      ldq_7_bits_uop_br_mask <=
        ldq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_746)	// lsu.scala:304:5, :306:44
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_650)	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_865) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_7_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_7_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_7_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_7_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_7_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_7_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_7_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_7_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_7_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_7_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_7_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_746)	// lsu.scala:304:5, :306:44
      ldq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_650)	// lsu.scala:210:16, :304:5, :305:44
      ldq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_762)	// lsu.scala:210:16, :304:5, :306:44
      ldq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_7_bits_uop_ppred_busy <= ~_GEN_762 & ldq_7_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_7_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h7
      | (_GEN_746
           ? io_core_dis_uops_1_bits_exception
           : _GEN_650 ? io_core_dis_uops_0_bits_exception : ldq_7_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_7_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1417
      & (_GEN_1363 ? ~_GEN_1322 & _GEN_866 : ~_GEN_1370 & _GEN_866);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_7_bits_executed <=
      ~_GEN_1476 & _GEN_1417 & _GEN_1386
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_580))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_955 & _GEN_1255 : ~(_GEN_569 & _GEN_955) & _GEN_1255)
            : _GEN_1255)
         | (dis_ld_val_1
              ? ~_GEN_714 & ldq_7_bits_executed
              : ~_GEN_650 & ldq_7_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_7_bits_succeeded <=
      _GEN_1417 & _GEN_1386
      & (_GEN_1282
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h7
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_714 & ldq_7_bits_succeeded
                    : ~_GEN_650 & ldq_7_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_7_bits_order_fail <=
      _GEN_1417 & _GEN_1386
      & (_GEN_361
           ? _GEN_778
           : _GEN_365
               ? _GEN_975 | _GEN_778
               : _GEN_366 & searcher_is_older_7 & _GEN_976 | _GEN_778);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_7_bits_observed <=
      _GEN_361
      | (dis_ld_val_1
           ? ~_GEN_714 & ldq_7_bits_observed
           : ~_GEN_650 & ldq_7_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_7_bits_forward_std_val <=
      _GEN_1417 & _GEN_1386
      & (~_GEN_590 & _GEN_1281
         | (dis_ld_val_1
              ? ~_GEN_714 & ldq_7_bits_forward_std_val
              : ~_GEN_650 & ldq_7_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1282) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_7_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_8_valid <=
      ~_GEN_1476 & _GEN_1418
      & (_GEN_1363 ? ~_GEN_1323 & _GEN_718 : ~_GEN_1371 & _GEN_718);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_747) begin	// lsu.scala:304:5, :306:44
      ldq_8_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_8_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_8_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_8_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_8_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_8_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_651) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_8_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_8_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_8_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_8_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_8_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_8_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_8_valid)	// lsu.scala:210:16
      ldq_8_bits_uop_br_mask <=
        ldq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_747)	// lsu.scala:304:5, :306:44
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_651)	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_867) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_8_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_8_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_8_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_8_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_8_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_8_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_8_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_8_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_8_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_8_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_8_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_747)	// lsu.scala:304:5, :306:44
      ldq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_651)	// lsu.scala:210:16, :304:5, :305:44
      ldq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_763)	// lsu.scala:210:16, :304:5, :306:44
      ldq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_8_bits_uop_ppred_busy <= ~_GEN_763 & ldq_8_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_8_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h8
      | (_GEN_747
           ? io_core_dis_uops_1_bits_exception
           : _GEN_651 ? io_core_dis_uops_0_bits_exception : ldq_8_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_8_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1418
      & (_GEN_1363 ? ~_GEN_1323 & _GEN_868 : ~_GEN_1371 & _GEN_868);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_8_bits_executed <=
      ~_GEN_1476 & _GEN_1418 & _GEN_1387
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_581))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_956 & _GEN_1256 : ~(_GEN_569 & _GEN_956) & _GEN_1256)
            : _GEN_1256)
         | (dis_ld_val_1
              ? ~_GEN_717 & ldq_8_bits_executed
              : ~_GEN_651 & ldq_8_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_8_bits_succeeded <=
      _GEN_1418 & _GEN_1387
      & (_GEN_1284
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h8
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_717 & ldq_8_bits_succeeded
                    : ~_GEN_651 & ldq_8_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_8_bits_order_fail <=
      _GEN_1418 & _GEN_1387
      & (_GEN_372
           ? _GEN_779
           : _GEN_376
               ? _GEN_977 | _GEN_779
               : _GEN_377 & searcher_is_older_8 & _GEN_978 | _GEN_779);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_8_bits_observed <=
      _GEN_372
      | (dis_ld_val_1
           ? ~_GEN_717 & ldq_8_bits_observed
           : ~_GEN_651 & ldq_8_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_8_bits_forward_std_val <=
      _GEN_1418 & _GEN_1387
      & (~_GEN_590 & _GEN_1283
         | (dis_ld_val_1
              ? ~_GEN_717 & ldq_8_bits_forward_std_val
              : ~_GEN_651 & ldq_8_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1284) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_8_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_9_valid <=
      ~_GEN_1476 & _GEN_1419
      & (_GEN_1363 ? ~_GEN_1324 & _GEN_721 : ~_GEN_1372 & _GEN_721);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_748) begin	// lsu.scala:304:5, :306:44
      ldq_9_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_9_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_9_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_9_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_9_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_9_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_652) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_9_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_9_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_9_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_9_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_9_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_9_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_9_valid)	// lsu.scala:210:16
      ldq_9_bits_uop_br_mask <=
        ldq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_748)	// lsu.scala:304:5, :306:44
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_652)	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_869) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_9_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_9_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_9_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_9_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_9_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_9_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_9_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_9_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_9_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_9_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_9_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_748)	// lsu.scala:304:5, :306:44
      ldq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_652)	// lsu.scala:210:16, :304:5, :305:44
      ldq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_764)	// lsu.scala:210:16, :304:5, :306:44
      ldq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_9_bits_uop_ppred_busy <= ~_GEN_764 & ldq_9_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_9_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'h9
      | (_GEN_748
           ? io_core_dis_uops_1_bits_exception
           : _GEN_652 ? io_core_dis_uops_0_bits_exception : ldq_9_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_9_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1419
      & (_GEN_1363 ? ~_GEN_1324 & _GEN_870 : ~_GEN_1372 & _GEN_870);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_9_bits_executed <=
      ~_GEN_1476 & _GEN_1419 & _GEN_1388
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_582))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_957 & _GEN_1257 : ~(_GEN_569 & _GEN_957) & _GEN_1257)
            : _GEN_1257)
         | (dis_ld_val_1
              ? ~_GEN_720 & ldq_9_bits_executed
              : ~_GEN_652 & ldq_9_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_9_bits_succeeded <=
      _GEN_1419 & _GEN_1388
      & (_GEN_1286
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'h9
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_720 & ldq_9_bits_succeeded
                    : ~_GEN_652 & ldq_9_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_9_bits_order_fail <=
      _GEN_1419 & _GEN_1388
      & (_GEN_383
           ? _GEN_780
           : _GEN_387
               ? _GEN_979 | _GEN_780
               : _GEN_388 & searcher_is_older_9 & _GEN_980 | _GEN_780);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_9_bits_observed <=
      _GEN_383
      | (dis_ld_val_1
           ? ~_GEN_720 & ldq_9_bits_observed
           : ~_GEN_652 & ldq_9_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_9_bits_forward_std_val <=
      _GEN_1419 & _GEN_1388
      & (~_GEN_590 & _GEN_1285
         | (dis_ld_val_1
              ? ~_GEN_720 & ldq_9_bits_forward_std_val
              : ~_GEN_652 & ldq_9_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1286) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_9_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_10_valid <=
      ~_GEN_1476 & _GEN_1420
      & (_GEN_1363 ? ~_GEN_1325 & _GEN_724 : ~_GEN_1373 & _GEN_724);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_749) begin	// lsu.scala:304:5, :306:44
      ldq_10_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_10_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_10_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_10_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_10_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_10_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_653) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_10_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_10_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_10_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_10_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_10_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_10_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_10_valid)	// lsu.scala:210:16
      ldq_10_bits_uop_br_mask <=
        ldq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_749)	// lsu.scala:304:5, :306:44
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_653)	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_871) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_10_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_10_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_10_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_10_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_10_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_10_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_10_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_10_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_10_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_10_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_10_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_749)	// lsu.scala:304:5, :306:44
      ldq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_653)	// lsu.scala:210:16, :304:5, :305:44
      ldq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_765)	// lsu.scala:210:16, :304:5, :306:44
      ldq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_10_bits_uop_ppred_busy <= ~_GEN_765 & ldq_10_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_10_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'hA
      | (_GEN_749
           ? io_core_dis_uops_1_bits_exception
           : _GEN_653 ? io_core_dis_uops_0_bits_exception : ldq_10_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_10_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1420
      & (_GEN_1363 ? ~_GEN_1325 & _GEN_872 : ~_GEN_1373 & _GEN_872);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_10_bits_executed <=
      ~_GEN_1476 & _GEN_1420 & _GEN_1389
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_583))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_958 & _GEN_1258 : ~(_GEN_569 & _GEN_958) & _GEN_1258)
            : _GEN_1258)
         | (dis_ld_val_1
              ? ~_GEN_723 & ldq_10_bits_executed
              : ~_GEN_653 & ldq_10_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_10_bits_succeeded <=
      _GEN_1420 & _GEN_1389
      & (_GEN_1288
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'hA
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_723 & ldq_10_bits_succeeded
                    : ~_GEN_653 & ldq_10_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_10_bits_order_fail <=
      _GEN_1420 & _GEN_1389
      & (_GEN_394
           ? _GEN_781
           : _GEN_398
               ? _GEN_981 | _GEN_781
               : _GEN_399 & searcher_is_older_10 & _GEN_982 | _GEN_781);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_10_bits_observed <=
      _GEN_394
      | (dis_ld_val_1
           ? ~_GEN_723 & ldq_10_bits_observed
           : ~_GEN_653 & ldq_10_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_10_bits_forward_std_val <=
      _GEN_1420 & _GEN_1389
      & (~_GEN_590 & _GEN_1287
         | (dis_ld_val_1
              ? ~_GEN_723 & ldq_10_bits_forward_std_val
              : ~_GEN_653 & ldq_10_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1288) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_10_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_11_valid <=
      ~_GEN_1476 & _GEN_1421
      & (_GEN_1363 ? ~_GEN_1326 & _GEN_727 : ~_GEN_1374 & _GEN_727);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_750) begin	// lsu.scala:304:5, :306:44
      ldq_11_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_11_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_11_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_11_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_11_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_11_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_654) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_11_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_11_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_11_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_11_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_11_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_11_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_11_valid)	// lsu.scala:210:16
      ldq_11_bits_uop_br_mask <=
        ldq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_750)	// lsu.scala:304:5, :306:44
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_654)	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_873) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_11_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_11_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_11_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_11_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_11_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_11_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_11_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_11_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_11_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_11_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_11_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_750)	// lsu.scala:304:5, :306:44
      ldq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_654)	// lsu.scala:210:16, :304:5, :305:44
      ldq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_766)	// lsu.scala:210:16, :304:5, :306:44
      ldq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_11_bits_uop_ppred_busy <= ~_GEN_766 & ldq_11_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_11_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'hB
      | (_GEN_750
           ? io_core_dis_uops_1_bits_exception
           : _GEN_654 ? io_core_dis_uops_0_bits_exception : ldq_11_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_11_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1421
      & (_GEN_1363 ? ~_GEN_1326 & _GEN_874 : ~_GEN_1374 & _GEN_874);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_11_bits_executed <=
      ~_GEN_1476 & _GEN_1421 & _GEN_1390
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_584))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_959 & _GEN_1259 : ~(_GEN_569 & _GEN_959) & _GEN_1259)
            : _GEN_1259)
         | (dis_ld_val_1
              ? ~_GEN_726 & ldq_11_bits_executed
              : ~_GEN_654 & ldq_11_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_11_bits_succeeded <=
      _GEN_1421 & _GEN_1390
      & (_GEN_1290
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'hB
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_726 & ldq_11_bits_succeeded
                    : ~_GEN_654 & ldq_11_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_11_bits_order_fail <=
      _GEN_1421 & _GEN_1390
      & (_GEN_405
           ? _GEN_782
           : _GEN_409
               ? _GEN_983 | _GEN_782
               : _GEN_410 & searcher_is_older_11 & _GEN_984 | _GEN_782);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_11_bits_observed <=
      _GEN_405
      | (dis_ld_val_1
           ? ~_GEN_726 & ldq_11_bits_observed
           : ~_GEN_654 & ldq_11_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_11_bits_forward_std_val <=
      _GEN_1421 & _GEN_1390
      & (~_GEN_590 & _GEN_1289
         | (dis_ld_val_1
              ? ~_GEN_726 & ldq_11_bits_forward_std_val
              : ~_GEN_654 & ldq_11_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1290) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_11_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_12_valid <=
      ~_GEN_1476 & _GEN_1422
      & (_GEN_1363 ? ~_GEN_1327 & _GEN_730 : ~_GEN_1375 & _GEN_730);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_751) begin	// lsu.scala:304:5, :306:44
      ldq_12_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_12_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_12_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_12_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_12_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_12_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_655) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_12_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_12_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_12_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_12_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_12_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_12_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_12_valid)	// lsu.scala:210:16
      ldq_12_bits_uop_br_mask <=
        ldq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_751)	// lsu.scala:304:5, :306:44
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_655)	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_875) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_12_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_12_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_12_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_12_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_12_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_12_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_12_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_12_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_12_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_12_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_12_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_751)	// lsu.scala:304:5, :306:44
      ldq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_655)	// lsu.scala:210:16, :304:5, :305:44
      ldq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_767)	// lsu.scala:210:16, :304:5, :306:44
      ldq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_12_bits_uop_ppred_busy <= ~_GEN_767 & ldq_12_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_12_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'hC
      | (_GEN_751
           ? io_core_dis_uops_1_bits_exception
           : _GEN_655 ? io_core_dis_uops_0_bits_exception : ldq_12_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_12_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1422
      & (_GEN_1363 ? ~_GEN_1327 & _GEN_876 : ~_GEN_1375 & _GEN_876);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_12_bits_executed <=
      ~_GEN_1476 & _GEN_1422 & _GEN_1391
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_585))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_960 & _GEN_1260 : ~(_GEN_569 & _GEN_960) & _GEN_1260)
            : _GEN_1260)
         | (dis_ld_val_1
              ? ~_GEN_729 & ldq_12_bits_executed
              : ~_GEN_655 & ldq_12_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_12_bits_succeeded <=
      _GEN_1422 & _GEN_1391
      & (_GEN_1292
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'hC
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_729 & ldq_12_bits_succeeded
                    : ~_GEN_655 & ldq_12_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_12_bits_order_fail <=
      _GEN_1422 & _GEN_1391
      & (_GEN_416
           ? _GEN_783
           : _GEN_420
               ? _GEN_985 | _GEN_783
               : _GEN_421 & searcher_is_older_12 & _GEN_986 | _GEN_783);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_12_bits_observed <=
      _GEN_416
      | (dis_ld_val_1
           ? ~_GEN_729 & ldq_12_bits_observed
           : ~_GEN_655 & ldq_12_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_12_bits_forward_std_val <=
      _GEN_1422 & _GEN_1391
      & (~_GEN_590 & _GEN_1291
         | (dis_ld_val_1
              ? ~_GEN_729 & ldq_12_bits_forward_std_val
              : ~_GEN_655 & ldq_12_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1292) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_12_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_13_valid <=
      ~_GEN_1476 & _GEN_1423
      & (_GEN_1363 ? ~_GEN_1328 & _GEN_733 : ~_GEN_1376 & _GEN_733);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_752) begin	// lsu.scala:304:5, :306:44
      ldq_13_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_13_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_13_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_13_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_13_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_13_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_656) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_13_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_13_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_13_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_13_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_13_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_13_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_13_valid)	// lsu.scala:210:16
      ldq_13_bits_uop_br_mask <=
        ldq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_752)	// lsu.scala:304:5, :306:44
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_656)	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_877) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_13_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_13_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_13_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_13_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_13_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_13_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_13_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_13_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_13_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_13_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_13_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_752)	// lsu.scala:304:5, :306:44
      ldq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_656)	// lsu.scala:210:16, :304:5, :305:44
      ldq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_768)	// lsu.scala:210:16, :304:5, :306:44
      ldq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_13_bits_uop_ppred_busy <= ~_GEN_768 & ldq_13_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_13_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'hD
      | (_GEN_752
           ? io_core_dis_uops_1_bits_exception
           : _GEN_656 ? io_core_dis_uops_0_bits_exception : ldq_13_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_13_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1423
      & (_GEN_1363 ? ~_GEN_1328 & _GEN_878 : ~_GEN_1376 & _GEN_878);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_13_bits_executed <=
      ~_GEN_1476 & _GEN_1423 & _GEN_1392
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_586))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_961 & _GEN_1261 : ~(_GEN_569 & _GEN_961) & _GEN_1261)
            : _GEN_1261)
         | (dis_ld_val_1
              ? ~_GEN_732 & ldq_13_bits_executed
              : ~_GEN_656 & ldq_13_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_13_bits_succeeded <=
      _GEN_1423 & _GEN_1392
      & (_GEN_1294
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'hD
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_732 & ldq_13_bits_succeeded
                    : ~_GEN_656 & ldq_13_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_13_bits_order_fail <=
      _GEN_1423 & _GEN_1392
      & (_GEN_427
           ? _GEN_784
           : _GEN_431
               ? _GEN_987 | _GEN_784
               : _GEN_432 & searcher_is_older_13 & _GEN_988 | _GEN_784);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_13_bits_observed <=
      _GEN_427
      | (dis_ld_val_1
           ? ~_GEN_732 & ldq_13_bits_observed
           : ~_GEN_656 & ldq_13_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_13_bits_forward_std_val <=
      _GEN_1423 & _GEN_1392
      & (~_GEN_590 & _GEN_1293
         | (dis_ld_val_1
              ? ~_GEN_732 & ldq_13_bits_forward_std_val
              : ~_GEN_656 & ldq_13_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1294) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_13_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_14_valid <=
      ~_GEN_1476 & _GEN_1424
      & (_GEN_1363 ? ~_GEN_1329 & _GEN_736 : ~_GEN_1377 & _GEN_736);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_753) begin	// lsu.scala:304:5, :306:44
      ldq_14_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_14_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_14_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_14_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_14_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_14_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_657) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_14_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_14_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_14_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_14_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_14_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_14_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_14_valid)	// lsu.scala:210:16
      ldq_14_bits_uop_br_mask <=
        ldq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_753)	// lsu.scala:304:5, :306:44
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_657)	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_879) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_14_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_14_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_14_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_14_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_14_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_14_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_14_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_14_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_14_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_14_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_14_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_753)	// lsu.scala:304:5, :306:44
      ldq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_657)	// lsu.scala:210:16, :304:5, :305:44
      ldq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_769)	// lsu.scala:210:16, :304:5, :306:44
      ldq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_14_bits_uop_ppred_busy <= ~_GEN_769 & ldq_14_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_14_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 4'hE
      | (_GEN_753
           ? io_core_dis_uops_1_bits_exception
           : _GEN_657 ? io_core_dis_uops_0_bits_exception : ldq_14_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_14_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1424
      & (_GEN_1363 ? ~_GEN_1329 & _GEN_880 : ~_GEN_1377 & _GEN_880);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_14_bits_executed <=
      ~_GEN_1476 & _GEN_1424 & _GEN_1393
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_587))
      & ((_GEN_565
            ? (_GEN_1264 ? ~_GEN_962 & _GEN_1262 : ~(_GEN_569 & _GEN_962) & _GEN_1262)
            : _GEN_1262)
         | (dis_ld_val_1
              ? ~_GEN_735 & ldq_14_bits_executed
              : ~_GEN_657 & ldq_14_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_14_bits_succeeded <=
      _GEN_1424 & _GEN_1393
      & (_GEN_1296
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & io_dmem_resp_0_bits_uop_ldq_idx == 4'hE
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_735 & ldq_14_bits_succeeded
                    : ~_GEN_657 & ldq_14_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_14_bits_order_fail <=
      _GEN_1424 & _GEN_1393
      & (_GEN_438
           ? _GEN_785
           : _GEN_442
               ? _GEN_989 | _GEN_785
               : _GEN_443 & searcher_is_older_14 & _GEN_990 | _GEN_785);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:72
    ldq_14_bits_observed <=
      _GEN_438
      | (dis_ld_val_1
           ? ~_GEN_735 & ldq_14_bits_observed
           : ~_GEN_657 & ldq_14_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_14_bits_forward_std_val <=
      _GEN_1424 & _GEN_1393
      & (~_GEN_590 & _GEN_1295
         | (dis_ld_val_1
              ? ~_GEN_735 & ldq_14_bits_forward_std_val
              : ~_GEN_657 & ldq_14_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1296) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_14_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    ldq_15_valid <=
      ~_GEN_1476 & _GEN_1425
      & (_GEN_1363 ? ~_GEN_1330 & _GEN_738 : ~_GEN_1378 & _GEN_738);	// lsu.scala:210:16, :304:5, :305:44, :1424:5, :1427:7, :1428:32, :1455:5, :1457:31, :1462:38, :1596:22, :1597:3, :1634:30
    if (_GEN_754) begin	// lsu.scala:304:5, :306:44
      ldq_15_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:210:16
      ldq_15_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:210:16
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:210:16
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;	// lsu.scala:210:16
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:210:16
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:210:16
      ldq_15_bits_uop_taken <= io_core_dis_uops_1_bits_taken;	// lsu.scala:210:16
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:210:16
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:210:16
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:210:16
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:210:16
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;	// lsu.scala:210:16
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;	// lsu.scala:210:16
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;	// lsu.scala:210:16
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_15_bits_st_dep_mask <= _GEN_691;	// lsu.scala:210:16, :336:31
      if (dis_st_val)	// lsu.scala:302:85
        ldq_15_bits_youngest_stq_idx <= _GEN_96;	// lsu.scala:210:16, util.scala:203:14
      else	// lsu.scala:302:85
        ldq_15_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else if (_GEN_658) begin	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:210:16
      ldq_15_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:210:16
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:210:16
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;	// lsu.scala:210:16
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;	// lsu.scala:210:16
      ldq_15_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;	// lsu.scala:210:16
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;	// lsu.scala:210:16
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:210:16
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;	// lsu.scala:210:16
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:210:16
      ldq_15_bits_uop_taken <= io_core_dis_uops_0_bits_taken;	// lsu.scala:210:16
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:210:16
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:210:16
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:210:16
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;	// lsu.scala:210:16
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:210:16
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:210:16
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:210:16
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;	// lsu.scala:210:16
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;	// lsu.scala:210:16
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;	// lsu.scala:210:16
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;	// lsu.scala:210:16
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;	// lsu.scala:210:16
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;	// lsu.scala:210:16
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:210:16
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;	// lsu.scala:210:16
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:210:16
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;	// lsu.scala:210:16
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;	// lsu.scala:210:16
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;	// lsu.scala:210:16
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:210:16
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:210:16
      ldq_15_bits_st_dep_mask <= next_live_store_mask;	// lsu.scala:210:16, :260:33
      ldq_15_bits_youngest_stq_idx <= stq_tail;	// lsu.scala:210:16, :218:29
    end
    else	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_st_dep_mask <=
        (_GEN_642 | ~_ldq_15_bits_st_dep_mask_T) & ldq_15_bits_st_dep_mask;	// lsu.scala:210:16, :260:{33,71}, :277:5, :278:{31,60}
    if (ldq_15_valid)	// lsu.scala:210:16
      ldq_15_bits_uop_br_mask <=
        ldq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:210:16, util.scala:85:27, :89:21
    else if (_GEN_754)	// lsu.scala:304:5, :306:44
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:210:16
    else if (_GEN_658)	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:210:16
    if (_GEN_881) begin	// lsu.scala:304:5, :836:5, :838:45
      if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
        ldq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:210:16
      else if (will_fire_load_retry_0)	// lsu.scala:535:65
        ldq_15_bits_uop_pdst <= _GEN_146;	// lsu.scala:210:16, :465:79
      else if (will_fire_sta_retry_0)	// lsu.scala:536:61
        ldq_15_bits_uop_pdst <= _GEN_199;	// lsu.scala:210:16, :478:79
      else	// lsu.scala:536:61
        ldq_15_bits_uop_pdst <= 7'h0;	// lsu.scala:210:16
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          ldq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:210:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          ldq_15_bits_addr_bits <= _GEN_269;	// lsu.scala:210:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          ldq_15_bits_addr_bits <= _GEN_191;	// lsu.scala:210:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          ldq_15_bits_addr_bits <= _GEN_200;	// lsu.scala:210:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          ldq_15_bits_addr_bits <= hella_req_addr;	// lsu.scala:210:16, :243:34
        else	// lsu.scala:535:65
          ldq_15_bits_addr_bits <= 40'h0;	// lsu.scala:210:16
      end
      else	// lsu.scala:708:58
        ldq_15_bits_addr_bits <= _GEN_270;	// lsu.scala:210:16, :768:30
      ldq_15_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:210:16, :708:58
      ldq_15_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;	// lsu.scala:210:16, :842:71
    end
    else if (_GEN_754)	// lsu.scala:304:5, :306:44
      ldq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:210:16
    else if (_GEN_658)	// lsu.scala:210:16, :304:5, :305:44
      ldq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:210:16
    if (_GEN_770)	// lsu.scala:210:16, :304:5, :306:44
      ldq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:210:16
    ldq_15_bits_uop_ppred_busy <= ~_GEN_770 & ldq_15_bits_uop_ppred_busy;	// lsu.scala:210:16, :304:5, :306:44
    ldq_15_bits_uop_exception <=
      mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & (&mem_xcpt_uops_0_ldq_idx)
      | (_GEN_754
           ? io_core_dis_uops_1_bits_exception
           : _GEN_658 ? io_core_dis_uops_0_bits_exception : ldq_15_bits_uop_exception);	// lsu.scala:210:16, :304:5, :305:44, :306:44, :667:32, :671:32, :717:5, :723:7, :724:58
    ldq_15_bits_addr_valid <=
      ~_GEN_1476 & _GEN_1425
      & (_GEN_1363 ? ~_GEN_1330 & _GEN_882 : ~_GEN_1378 & _GEN_882);	// lsu.scala:210:16, :304:5, :836:5, :838:45, :1424:5, :1427:7, :1428:32, :1429:32, :1455:5, :1457:31, :1462:38, :1463:38, :1596:22, :1597:3, :1634:30, :1635:30
    ldq_15_bits_executed <=
      ~_GEN_1476 & _GEN_1425 & _GEN_1394
      & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
         | ~(io_dmem_nack_0_bits_uop_uses_ldq & (&io_dmem_nack_0_bits_uop_ldq_idx)))
      & ((_GEN_565
            ? (_GEN_1264
                 ? ~(&lcam_ldq_idx_0) & _GEN_1263
                 : ~(_GEN_569 & (&lcam_ldq_idx_0)) & _GEN_1263)
            : _GEN_1263)
         | (dis_ld_val_1
              ? ~_GEN_737 & ldq_15_bits_executed
              : ~_GEN_658 & ldq_15_bits_executed));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :311:44, :1036:26, :1091:36, :1130:48, :1148:{45,72}, :1150:9, :1154:46, :1157:9, :1162:37, :1163:9, :1166:46, :1174:{30,53}, :1284:5, :1287:7, :1291:7, :1293:62, :1455:5, :1457:31, :1596:22, :1597:3, :1634:30, :1636:30
    ldq_15_bits_succeeded <=
      _GEN_1425 & _GEN_1394
      & (_GEN_1298
           ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq
              & (&io_dmem_resp_0_bits_uop_ldq_idx)
                ? _ldq_bits_succeeded_T
                : dis_ld_val_1
                    ? ~_GEN_737 & ldq_15_bits_succeeded
                    : ~_GEN_658 & ldq_15_bits_succeeded)
           : _GEN_600);	// AMOALU.scala:10:17, lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :312:44, :1284:5, :1306:5, :1308:7, :1324:{42,72}, :1344:5, :1348:5, :1455:5, :1457:31
    ldq_15_bits_order_fail <=
      _GEN_1425 & _GEN_1394
      & (_GEN_449
           ? _GEN_786
           : _GEN_453
               ? _GEN_992 | _GEN_786
               : _GEN_454 & searcher_is_older_15 & _GEN_993 | _GEN_786);	// lsu.scala:210:16, :304:5, :313:44, :1090:34, :1091:36, :1101:131, :1102:37, :1106:39, :1107:76, :1108:34, :1115:47, :1116:37, :1118:34, :1120:40, :1121:34, :1122:36, :1284:5, :1455:5, :1457:31, util.scala:363:58
    ldq_15_bits_observed <=
      _GEN_449
      | (dis_ld_val_1
           ? ~_GEN_737 & ldq_15_bits_observed
           : ~_GEN_658 & ldq_15_bits_observed);	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :314:44, :1090:34, :1091:36, :1094:30
    ldq_15_bits_forward_std_val <=
      _GEN_1425 & _GEN_1394
      & (~_GEN_590 & _GEN_1297
         | (dis_ld_val_1
              ? ~_GEN_737 & ldq_15_bits_forward_std_val
              : ~_GEN_658 & ldq_15_bits_forward_std_val));	// lsu.scala:210:16, :301:85, :304:5, :305:44, :310:44, :315:44, :1284:5, :1306:5, :1343:30, :1344:5, :1348:5, :1369:33, :1370:35, :1455:5, :1457:31
    if (_GEN_1298) begin	// lsu.scala:210:16, :1306:5, :1344:5, :1348:5
    end
    else	// lsu.scala:210:16, :1344:5, :1348:5
      ldq_15_bits_forward_stq_idx <= wb_forward_stq_idx_0;	// lsu.scala:210:16, :1067:36
    stq_0_valid <=
      ~_GEN_1479 & (clear_store ? ~_GEN_1427 & _GEN_788 : ~_GEN_1299 & _GEN_788);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    if (_GEN_1477) begin	// lsu.scala:1505:3, :1597:3, :1602:5, :1603:16
      stq_0_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_0_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_0_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_0_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_0_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_0_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_0_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_0_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_0_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_0_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_0_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_0_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_0_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_0_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_0_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_1_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_1_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_1_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_1_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_1_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_1_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_1_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_1_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_1_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_1_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_1_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_1_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_1_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_1_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_2_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_2_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_2_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_2_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_2_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_2_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_2_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_2_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_2_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_2_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_2_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_2_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_2_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_2_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_3_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_3_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_3_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_3_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_3_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_3_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_3_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_3_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_3_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_3_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_3_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_3_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_3_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_3_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_4_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_4_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_4_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_4_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_4_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_4_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_4_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_4_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_4_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_4_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_4_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_4_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_4_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_4_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_5_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_5_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_5_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_5_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_5_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_5_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_5_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_5_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_5_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_5_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_5_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_5_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_5_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_5_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_6_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_6_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_6_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_6_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_6_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_6_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_6_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_6_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_6_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_6_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_6_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_6_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_6_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_6_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_7_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_7_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_7_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_7_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_7_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_7_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_7_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_7_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_7_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_7_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_7_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_7_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_7_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_7_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_8_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_8_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_8_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_8_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_8_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_8_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_8_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_8_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_8_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_8_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_8_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_8_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_8_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_8_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_9_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_9_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_9_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_9_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_9_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_9_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_9_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_9_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_9_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_9_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_9_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_9_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_9_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_9_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_10_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_10_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_10_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_10_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_10_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_10_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_10_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_10_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_10_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_10_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_10_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_10_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_10_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_10_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_11_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_11_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_11_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_11_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_11_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_11_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_11_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_11_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_11_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_11_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_11_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_11_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_11_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_11_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_12_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_12_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_12_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_12_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_12_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_12_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_12_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_12_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_12_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_12_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_12_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_12_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_12_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_12_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_13_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_13_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_13_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_13_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_13_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_13_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_13_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_13_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_13_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_13_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_13_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_13_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_13_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_13_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_14_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_14_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_14_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_14_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_14_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_14_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_14_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_14_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_14_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_14_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_14_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_14_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_14_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_14_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_uopc <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_inst <= 32'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_inst <= 32'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_pc <= 40'h0;	// lsu.scala:211:16
      stq_15_bits_uop_iq_type <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_fu_code <= 10'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_br_type <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_op1_sel <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_op2_sel <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_imm_sel <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_op_fcn <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ctrl_csr_cmd <= 3'h0;	// lsu.scala:211:16
      stq_15_bits_uop_iw_state <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_br_mask <= 12'h0;	// lsu.scala:211:16
      stq_15_bits_uop_br_tag <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ftq_idx <= 5'h0;	// lsu.scala:211:16
      stq_15_bits_uop_pc_lob <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_imm_packed <= 20'h0;	// lsu.scala:211:16
      stq_15_bits_uop_csr_addr <= 12'h0;	// lsu.scala:211:16
      stq_15_bits_uop_rob_idx <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ldq_idx <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_stq_idx <= 4'h0;	// lsu.scala:211:16
      stq_15_bits_uop_rxq_idx <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_prs1 <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_prs2 <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_prs3 <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      stq_15_bits_uop_stale_pdst <= 7'h0;	// lsu.scala:211:16
      stq_15_bits_uop_exc_cause <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:211:16, :249:20
      stq_15_bits_uop_mem_cmd <= 5'h0;	// lsu.scala:211:16
      stq_15_bits_uop_mem_size <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_ldst <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs1 <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs2 <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs3 <= 6'h0;	// lsu.scala:211:16
      stq_15_bits_uop_dst_rtype <= 2'h2;	// lsu.scala:211:16, util.scala:351:72
      stq_15_bits_uop_lrs1_rtype <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_lrs2_rtype <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_fsrc <= 2'h0;	// lsu.scala:211:16
      stq_15_bits_uop_debug_tsrc <= 2'h0;	// lsu.scala:211:16
      stq_head <= 4'h0;	// lsu.scala:217:29
      stq_commit_head <= 4'h0;	// lsu.scala:219:29
      stq_execute_head <= 4'h0;	// lsu.scala:220:29
    end
    else begin	// lsu.scala:1505:3, :1597:3, :1602:5, :1603:16
      if (_GEN_819) begin	// lsu.scala:304:5, :321:5
        if (_GEN_675) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_0_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_0_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_0_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_0_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_0_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_0_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_0_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_0_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_0_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_0_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_0_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_0_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_0_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_0_valid)	// lsu.scala:211:16
        stq_0_bits_uop_br_mask <=
          stq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_819) begin	// lsu.scala:304:5, :321:5
        if (_GEN_675) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_819) begin	// lsu.scala:304:5, :321:5
        if (_GEN_675) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_0_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_0_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_0_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_0_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_0_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_0_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_0_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_0_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_0_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_0_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_0_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_883) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_0_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_0_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_0_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_819) begin	// lsu.scala:304:5, :321:5
        if (_GEN_675) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_819) begin	// lsu.scala:304:5, :321:5
        if (_GEN_675) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_0_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_0_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_0_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_0_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_0_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
      end
      if (dis_ld_val_1) begin	// lsu.scala:301:85
        if (_GEN_675) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_676) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_677) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_678) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_679) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_680) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_681) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_682) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_683) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_684) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_685) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_686) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_687) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_688) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_689) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_690) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      end
      else begin	// lsu.scala:301:85
        if (_GEN_787 | ~_GEN_675)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_0_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_789 | ~_GEN_676)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_1_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_791 | ~_GEN_677)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_2_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_793 | ~_GEN_678)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_3_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_795 | ~_GEN_679)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_4_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_797 | ~_GEN_680)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_5_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_799 | ~_GEN_681)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_6_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_801 | ~_GEN_682)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_7_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_803 | ~_GEN_683)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_8_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_805 | ~_GEN_684)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_9_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_807 | ~_GEN_685)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_10_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_809 | ~_GEN_686)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_11_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_811 | ~_GEN_687)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_12_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_813 | ~_GEN_688)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_13_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_815 | ~_GEN_689)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_14_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
        if (_GEN_817 | ~_GEN_690)	// lsu.scala:211:16, :304:5, :321:5, :322:39, :323:39
          stq_15_bits_uop_ppred <= 5'h0;	// lsu.scala:211:16
      end
      if (_GEN_819) begin	// lsu.scala:304:5, :321:5
        if (_GEN_675) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_0_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_0_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_0_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_0_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_0_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_0_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_0_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_0_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_0_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_0_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_0_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_0_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_820) begin	// lsu.scala:304:5, :321:5
        if (_GEN_676) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_1_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_1_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_1_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_1_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_1_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_1_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_1_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_1_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_1_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_1_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_1_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_1_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_1_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_1_valid)	// lsu.scala:211:16
        stq_1_bits_uop_br_mask <=
          stq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_820) begin	// lsu.scala:304:5, :321:5
        if (_GEN_676) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_820) begin	// lsu.scala:304:5, :321:5
        if (_GEN_676) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_1_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_1_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_1_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_1_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_1_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_1_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_1_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_1_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_1_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_1_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_1_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_885) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_1_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_1_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_1_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_820) begin	// lsu.scala:304:5, :321:5
        if (_GEN_676) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_820) begin	// lsu.scala:304:5, :321:5
        if (_GEN_676) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_1_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_1_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_1_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_1_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_1_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_1_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_1_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_1_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_1_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_1_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_1_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_1_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_1_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_1_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_1_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_1_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_1_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_1_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_821) begin	// lsu.scala:304:5, :321:5
        if (_GEN_677) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_2_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_2_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_2_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_2_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_2_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_2_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_2_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_2_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_2_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_2_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_2_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_2_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_2_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_2_valid)	// lsu.scala:211:16
        stq_2_bits_uop_br_mask <=
          stq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_821) begin	// lsu.scala:304:5, :321:5
        if (_GEN_677) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_821) begin	// lsu.scala:304:5, :321:5
        if (_GEN_677) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_2_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_2_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_2_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_2_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_2_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_2_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_2_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_2_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_2_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_2_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_2_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_887) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_2_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_2_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_2_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_821) begin	// lsu.scala:304:5, :321:5
        if (_GEN_677) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_821) begin	// lsu.scala:304:5, :321:5
        if (_GEN_677) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_2_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_2_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_2_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_2_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_2_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_2_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_2_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_2_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_2_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_2_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_2_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_2_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_2_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_2_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_2_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_2_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_2_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_2_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_822) begin	// lsu.scala:304:5, :321:5
        if (_GEN_678) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_3_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_3_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_3_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_3_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_3_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_3_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_3_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_3_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_3_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_3_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_3_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_3_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_3_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_3_valid)	// lsu.scala:211:16
        stq_3_bits_uop_br_mask <=
          stq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_822) begin	// lsu.scala:304:5, :321:5
        if (_GEN_678) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_822) begin	// lsu.scala:304:5, :321:5
        if (_GEN_678) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_3_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_3_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_3_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_3_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_3_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_3_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_3_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_3_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_3_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_3_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_3_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_889) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_3_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_3_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_3_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_822) begin	// lsu.scala:304:5, :321:5
        if (_GEN_678) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_822) begin	// lsu.scala:304:5, :321:5
        if (_GEN_678) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_3_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_3_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_3_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_3_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_3_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_3_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_3_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_3_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_3_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_3_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_3_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_3_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_3_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_3_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_3_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_3_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_3_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_3_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_823) begin	// lsu.scala:304:5, :321:5
        if (_GEN_679) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_4_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_4_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_4_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_4_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_4_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_4_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_4_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_4_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_4_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_4_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_4_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_4_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_4_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_4_valid)	// lsu.scala:211:16
        stq_4_bits_uop_br_mask <=
          stq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_823) begin	// lsu.scala:304:5, :321:5
        if (_GEN_679) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_823) begin	// lsu.scala:304:5, :321:5
        if (_GEN_679) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_4_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_4_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_4_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_4_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_4_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_4_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_4_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_4_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_4_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_4_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_4_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_891) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_4_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_4_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_4_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_823) begin	// lsu.scala:304:5, :321:5
        if (_GEN_679) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_823) begin	// lsu.scala:304:5, :321:5
        if (_GEN_679) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_4_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_4_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_4_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_4_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_4_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_4_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_4_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_4_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_4_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_4_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_4_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_4_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_4_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_4_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_4_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_4_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_4_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_4_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_824) begin	// lsu.scala:304:5, :321:5
        if (_GEN_680) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_5_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_5_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_5_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_5_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_5_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_5_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_5_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_5_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_5_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_5_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_5_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_5_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_5_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_5_valid)	// lsu.scala:211:16
        stq_5_bits_uop_br_mask <=
          stq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_824) begin	// lsu.scala:304:5, :321:5
        if (_GEN_680) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_824) begin	// lsu.scala:304:5, :321:5
        if (_GEN_680) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_5_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_5_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_5_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_5_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_5_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_5_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_5_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_5_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_5_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_5_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_5_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_893) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_5_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_5_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_5_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_824) begin	// lsu.scala:304:5, :321:5
        if (_GEN_680) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_824) begin	// lsu.scala:304:5, :321:5
        if (_GEN_680) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_5_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_5_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_5_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_5_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_5_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_5_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_5_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_5_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_5_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_5_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_5_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_5_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_5_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_5_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_5_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_5_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_5_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_5_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_825) begin	// lsu.scala:304:5, :321:5
        if (_GEN_681) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_6_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_6_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_6_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_6_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_6_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_6_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_6_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_6_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_6_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_6_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_6_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_6_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_6_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_6_valid)	// lsu.scala:211:16
        stq_6_bits_uop_br_mask <=
          stq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_825) begin	// lsu.scala:304:5, :321:5
        if (_GEN_681) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_825) begin	// lsu.scala:304:5, :321:5
        if (_GEN_681) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_6_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_6_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_6_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_6_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_6_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_6_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_6_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_6_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_6_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_6_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_6_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_895) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_6_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_6_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_6_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_825) begin	// lsu.scala:304:5, :321:5
        if (_GEN_681) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_825) begin	// lsu.scala:304:5, :321:5
        if (_GEN_681) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_6_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_6_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_6_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_6_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_6_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_6_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_6_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_6_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_6_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_6_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_6_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_6_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_6_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_6_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_6_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_6_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_6_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_6_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_826) begin	// lsu.scala:304:5, :321:5
        if (_GEN_682) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_7_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_7_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_7_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_7_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_7_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_7_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_7_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_7_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_7_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_7_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_7_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_7_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_7_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_7_valid)	// lsu.scala:211:16
        stq_7_bits_uop_br_mask <=
          stq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_826) begin	// lsu.scala:304:5, :321:5
        if (_GEN_682) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_826) begin	// lsu.scala:304:5, :321:5
        if (_GEN_682) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_7_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_7_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_7_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_7_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_7_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_7_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_7_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_7_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_7_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_7_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_7_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_897) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_7_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_7_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_7_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_826) begin	// lsu.scala:304:5, :321:5
        if (_GEN_682) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_826) begin	// lsu.scala:304:5, :321:5
        if (_GEN_682) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_7_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_7_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_7_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_7_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_7_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_7_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_7_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_7_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_7_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_7_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_7_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_7_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_7_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_7_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_7_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_7_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_7_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_7_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_827) begin	// lsu.scala:304:5, :321:5
        if (_GEN_683) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_8_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_8_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_8_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_8_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_8_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_8_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_8_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_8_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_8_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_8_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_8_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_8_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_8_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_8_valid)	// lsu.scala:211:16
        stq_8_bits_uop_br_mask <=
          stq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_827) begin	// lsu.scala:304:5, :321:5
        if (_GEN_683) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_827) begin	// lsu.scala:304:5, :321:5
        if (_GEN_683) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_8_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_8_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_8_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_8_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_8_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_8_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_8_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_8_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_8_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_8_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_8_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_899) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_8_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_8_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_8_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_827) begin	// lsu.scala:304:5, :321:5
        if (_GEN_683) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_827) begin	// lsu.scala:304:5, :321:5
        if (_GEN_683) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_8_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_8_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_8_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_8_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_8_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_8_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_8_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_8_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_8_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_8_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_8_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_8_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_8_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_8_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_8_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_8_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_8_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_8_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_828) begin	// lsu.scala:304:5, :321:5
        if (_GEN_684) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_9_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_9_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_9_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_9_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_9_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_9_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_9_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_9_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_9_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_9_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_9_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_9_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_9_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_9_valid)	// lsu.scala:211:16
        stq_9_bits_uop_br_mask <=
          stq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_828) begin	// lsu.scala:304:5, :321:5
        if (_GEN_684) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_828) begin	// lsu.scala:304:5, :321:5
        if (_GEN_684) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_9_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_9_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_9_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_9_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_9_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_9_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_9_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_9_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_9_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_9_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_9_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_901) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_9_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_9_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_9_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_828) begin	// lsu.scala:304:5, :321:5
        if (_GEN_684) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_828) begin	// lsu.scala:304:5, :321:5
        if (_GEN_684) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_9_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_9_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_9_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_9_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_9_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_9_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_9_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_9_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_9_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_9_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_9_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_9_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_9_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_9_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_9_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_9_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_9_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_9_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_829) begin	// lsu.scala:304:5, :321:5
        if (_GEN_685) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_10_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_10_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_10_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_10_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_10_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_10_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_10_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_10_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_10_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_10_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_10_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_10_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_10_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_10_valid)	// lsu.scala:211:16
        stq_10_bits_uop_br_mask <=
          stq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_829) begin	// lsu.scala:304:5, :321:5
        if (_GEN_685) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_829) begin	// lsu.scala:304:5, :321:5
        if (_GEN_685) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_10_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_10_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_10_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_10_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_10_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_10_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_10_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_10_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_10_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_10_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_10_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_903) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_10_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_10_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_10_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_829) begin	// lsu.scala:304:5, :321:5
        if (_GEN_685) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_829) begin	// lsu.scala:304:5, :321:5
        if (_GEN_685) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_10_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_10_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_10_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_10_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_10_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_10_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_10_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_10_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_10_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_10_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_10_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_10_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_10_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_10_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_10_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_10_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_10_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_10_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_830) begin	// lsu.scala:304:5, :321:5
        if (_GEN_686) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_11_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_11_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_11_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_11_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_11_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_11_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_11_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_11_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_11_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_11_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_11_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_11_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_11_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_11_valid)	// lsu.scala:211:16
        stq_11_bits_uop_br_mask <=
          stq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_830) begin	// lsu.scala:304:5, :321:5
        if (_GEN_686) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_830) begin	// lsu.scala:304:5, :321:5
        if (_GEN_686) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_11_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_11_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_11_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_11_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_11_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_11_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_11_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_11_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_11_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_11_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_11_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_905) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_11_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_11_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_11_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_830) begin	// lsu.scala:304:5, :321:5
        if (_GEN_686) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_830) begin	// lsu.scala:304:5, :321:5
        if (_GEN_686) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_11_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_11_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_11_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_11_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_11_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_11_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_11_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_11_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_11_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_11_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_11_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_11_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_11_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_11_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_11_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_11_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_11_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_11_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_831) begin	// lsu.scala:304:5, :321:5
        if (_GEN_687) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_12_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_12_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_12_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_12_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_12_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_12_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_12_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_12_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_12_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_12_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_12_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_12_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_12_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_12_valid)	// lsu.scala:211:16
        stq_12_bits_uop_br_mask <=
          stq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_831) begin	// lsu.scala:304:5, :321:5
        if (_GEN_687) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_831) begin	// lsu.scala:304:5, :321:5
        if (_GEN_687) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_12_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_12_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_12_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_12_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_12_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_12_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_12_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_12_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_12_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_12_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_12_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_907) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_12_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_12_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_12_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_831) begin	// lsu.scala:304:5, :321:5
        if (_GEN_687) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_831) begin	// lsu.scala:304:5, :321:5
        if (_GEN_687) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_12_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_12_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_12_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_12_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_12_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_12_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_12_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_12_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_12_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_12_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_12_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_12_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_12_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_12_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_12_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_12_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_12_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_12_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_832) begin	// lsu.scala:304:5, :321:5
        if (_GEN_688) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_13_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_13_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_13_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_13_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_13_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_13_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_13_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_13_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_13_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_13_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_13_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_13_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_13_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_13_valid)	// lsu.scala:211:16
        stq_13_bits_uop_br_mask <=
          stq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_832) begin	// lsu.scala:304:5, :321:5
        if (_GEN_688) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_832) begin	// lsu.scala:304:5, :321:5
        if (_GEN_688) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_13_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_13_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_13_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_13_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_13_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_13_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_13_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_13_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_13_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_13_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_13_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_909) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_13_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_13_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_13_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_832) begin	// lsu.scala:304:5, :321:5
        if (_GEN_688) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_832) begin	// lsu.scala:304:5, :321:5
        if (_GEN_688) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_13_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_13_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_13_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_13_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_13_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_13_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_13_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_13_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_13_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_13_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_13_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_13_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_13_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_13_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_13_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_13_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_13_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_13_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_833) begin	// lsu.scala:304:5, :321:5
        if (_GEN_689) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_14_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_14_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_14_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_14_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_14_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_14_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_14_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_14_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_14_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_14_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_14_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_14_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_14_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_14_valid)	// lsu.scala:211:16
        stq_14_bits_uop_br_mask <=
          stq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_833) begin	// lsu.scala:304:5, :321:5
        if (_GEN_689) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_833) begin	// lsu.scala:304:5, :321:5
        if (_GEN_689) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_14_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_14_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_14_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_14_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_14_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_14_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_14_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_14_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_14_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_14_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_14_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_911) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_14_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_14_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_14_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_833) begin	// lsu.scala:304:5, :321:5
        if (_GEN_689) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_833) begin	// lsu.scala:304:5, :321:5
        if (_GEN_689) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_14_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_14_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_14_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_14_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_14_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_14_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_14_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_14_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_14_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_14_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_14_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_14_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_14_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_14_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_14_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_14_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_14_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_14_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (_GEN_834) begin	// lsu.scala:304:5, :321:5
        if (_GEN_690) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_15_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;	// lsu.scala:211:16
          stq_15_bits_uop_inst <= io_core_dis_uops_0_bits_inst;	// lsu.scala:211:16
          stq_15_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;	// lsu.scala:211:16
          stq_15_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;	// lsu.scala:211:16
          stq_15_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;	// lsu.scala:211:16
          stq_15_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;	// lsu.scala:211:16
          stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;	// lsu.scala:211:16
          stq_15_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;	// lsu.scala:211:16
        stq_15_bits_uop_inst <= io_core_dis_uops_1_bits_inst;	// lsu.scala:211:16
        stq_15_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;	// lsu.scala:211:16
        stq_15_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;	// lsu.scala:211:16
        stq_15_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;	// lsu.scala:211:16
        stq_15_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;	// lsu.scala:211:16
        stq_15_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;	// lsu.scala:211:16
      end
      if (stq_15_valid)	// lsu.scala:211:16
        stq_15_bits_uop_br_mask <=
          stq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:211:16, util.scala:85:27, :89:21
      else if (_GEN_834) begin	// lsu.scala:304:5, :321:5
        if (_GEN_690) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;	// lsu.scala:211:16
      if (_GEN_834) begin	// lsu.scala:304:5, :321:5
        if (_GEN_690) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_15_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;	// lsu.scala:211:16
          stq_15_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;	// lsu.scala:211:16
          stq_15_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;	// lsu.scala:211:16
          stq_15_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;	// lsu.scala:211:16
          stq_15_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;	// lsu.scala:211:16
          stq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;	// lsu.scala:211:16
          stq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;	// lsu.scala:211:16
          stq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;	// lsu.scala:211:16
          stq_15_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;	// lsu.scala:211:16
        stq_15_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;	// lsu.scala:211:16
        stq_15_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;	// lsu.scala:211:16
        stq_15_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;	// lsu.scala:211:16
        stq_15_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;	// lsu.scala:211:16
        stq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;	// lsu.scala:211:16
        stq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;	// lsu.scala:211:16
        stq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;	// lsu.scala:211:16
        stq_15_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;	// lsu.scala:211:16
      end
      if (_GEN_913) begin	// lsu.scala:304:5, :849:5, :853:36
        if (_exe_tlb_uop_T_2)	// lsu.scala:599:53
          stq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:211:16
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_15_bits_uop_pdst <= _GEN_146;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_15_bits_uop_pdst <= _GEN_199;	// lsu.scala:211:16, :478:79
        else	// lsu.scala:536:61
          stq_15_bits_uop_pdst <= 7'h0;	// lsu.scala:211:16
      end
      else if (_GEN_834) begin	// lsu.scala:304:5, :321:5
        if (_GEN_690) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else	// lsu.scala:211:16, :304:5, :321:5
          stq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;	// lsu.scala:211:16
      end
      else	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;	// lsu.scala:211:16
      if (_GEN_834) begin	// lsu.scala:304:5, :321:5
        if (_GEN_690) begin	// lsu.scala:211:16, :304:5, :321:5
        end
        else begin	// lsu.scala:211:16, :304:5, :321:5
          stq_15_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;	// lsu.scala:211:16
          stq_15_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;	// lsu.scala:211:16
          stq_15_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;	// lsu.scala:211:16
          stq_15_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;	// lsu.scala:211:16
          stq_15_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;	// lsu.scala:211:16
          stq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;	// lsu.scala:211:16
          stq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;	// lsu.scala:211:16
          stq_15_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;	// lsu.scala:211:16
          stq_15_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;	// lsu.scala:211:16
          stq_15_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;	// lsu.scala:211:16
          stq_15_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;	// lsu.scala:211:16
          stq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;	// lsu.scala:211:16
          stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;	// lsu.scala:211:16
          stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;	// lsu.scala:211:16
          stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;	// lsu.scala:211:16
          stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;	// lsu.scala:211:16
        end
      end
      else begin	// lsu.scala:304:5, :321:5
        stq_15_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;	// lsu.scala:211:16
        stq_15_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;	// lsu.scala:211:16
        stq_15_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;	// lsu.scala:211:16
        stq_15_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;	// lsu.scala:211:16
        stq_15_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;	// lsu.scala:211:16
        stq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;	// lsu.scala:211:16
        stq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;	// lsu.scala:211:16
        stq_15_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;	// lsu.scala:211:16
        stq_15_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;	// lsu.scala:211:16
        stq_15_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;	// lsu.scala:211:16
        stq_15_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;	// lsu.scala:211:16
        stq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;	// lsu.scala:211:16
        stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;	// lsu.scala:211:16
        stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;	// lsu.scala:211:16
        stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;	// lsu.scala:211:16
        stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;	// lsu.scala:211:16
      end
      if (clear_store)	// lsu.scala:1495:3, :1500:17
        stq_head <= stq_head + 4'h1;	// lsu.scala:217:29, :305:44, util.scala:203:14
      if (commit_store_1)	// lsu.scala:1451:49
        stq_commit_head <= _GEN_622 + 4'h1;	// lsu.scala:219:29, :305:44, :1482:31, util.scala:203:14
      else if (commit_store)	// lsu.scala:1451:49
        stq_commit_head <= _GEN_621;	// lsu.scala:219:29, util.scala:203:14
      if (clear_store & _GEN_634)	// lsu.scala:1284:5, :1494:29, :1495:3, :1500:17, :1505:3, :1514:5, :1515:24
        stq_execute_head <= stq_execute_head + 4'h1;	// lsu.scala:220:29, :305:44, util.scala:203:14
      else if (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella
               | io_dmem_nack_0_bits_uop_uses_ldq
               | io_dmem_nack_0_bits_uop_stq_idx < stq_head ^ stq_execute_head < stq_head
               ^ io_dmem_nack_0_bits_uop_stq_idx >= stq_execute_head) begin	// lsu.scala:217:29, :220:29, :766:39, :1174:30, :1284:5, :1287:7, :1291:7, :1299:86, util.scala:363:{52,64,78}
        if (_GEN_272 | ~(will_fire_store_commit_0 & dmem_req_fire_0)) begin	// lsu.scala:220:29, :535:65, :752:55, :766:39, :773:43, :780:45, :789:{44,50}
        end
        else	// lsu.scala:220:29, :766:39, :773:43, :780:45
          stq_execute_head <= stq_execute_head + 4'h1;	// lsu.scala:220:29, :305:44, util.scala:203:14
      end
      else	// lsu.scala:766:39, :1284:5, :1287:7
        stq_execute_head <= io_dmem_nack_0_bits_uop_stq_idx;	// lsu.scala:220:29
    end
    stq_0_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675
                ? stq_0_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675
                ? stq_0_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675
                ? stq_0_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_819 & _GEN_675 & stq_0_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h0
         | (_GEN_819
              ? (_GEN_675 ? stq_0_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675
                ? stq_0_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675
                ? stq_0_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_819
           ? (_GEN_675 ? stq_0_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_0_bits_addr_valid <=
      ~_GEN_1479 & (clear_store ? ~_GEN_1427 & _GEN_884 : ~_GEN_1299 & _GEN_884);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_883) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_0_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_0_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_0_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_0_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_0_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_0_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_0_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_0_bits_data_valid <=
      ~_GEN_1479 & (clear_store ? ~_GEN_1427 & _GEN_916 : ~_GEN_1299 & _GEN_916);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_915) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_0_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_0_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_0_bits_committed <=
      ~_GEN_1457
      & (commit_store_1 ? _GEN_1395 | _GEN_1332 | _GEN_835 : _GEN_1332 | _GEN_835);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_0_bits_succeeded <=
      ~_GEN_1457
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h0
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h0)) & _GEN_819
         & _GEN_675 & stq_0_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_1_valid <=
      ~_GEN_1481 & (clear_store ? ~_GEN_1429 & _GEN_790 : ~_GEN_1300 & _GEN_790);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_1_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676
                ? stq_1_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676
                ? stq_1_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676
                ? stq_1_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_820 & _GEN_676 & stq_1_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h1
         | (_GEN_820
              ? (_GEN_676 ? stq_1_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676
                ? stq_1_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676
                ? stq_1_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_820
           ? (_GEN_676 ? stq_1_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_1_bits_addr_valid <=
      ~_GEN_1481 & (clear_store ? ~_GEN_1429 & _GEN_886 : ~_GEN_1300 & _GEN_886);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_885) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_1_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_1_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_1_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_1_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_1_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_1_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_1_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_1_bits_data_valid <=
      ~_GEN_1481 & (clear_store ? ~_GEN_1429 & _GEN_918 : ~_GEN_1300 & _GEN_918);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_917) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_1_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_1_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_1_bits_committed <=
      ~_GEN_1458
      & (commit_store_1 ? _GEN_1396 | _GEN_1334 | _GEN_836 : _GEN_1334 | _GEN_836);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_1_bits_succeeded <=
      ~_GEN_1458
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h1
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h1)) & _GEN_820
         & _GEN_676 & stq_1_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_2_valid <=
      ~_GEN_1483 & (clear_store ? ~_GEN_1431 & _GEN_792 : ~_GEN_1301 & _GEN_792);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_2_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677
                ? stq_2_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677
                ? stq_2_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677
                ? stq_2_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_821 & _GEN_677 & stq_2_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h2
         | (_GEN_821
              ? (_GEN_677 ? stq_2_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677
                ? stq_2_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677
                ? stq_2_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_821
           ? (_GEN_677 ? stq_2_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_2_bits_addr_valid <=
      ~_GEN_1483 & (clear_store ? ~_GEN_1431 & _GEN_888 : ~_GEN_1301 & _GEN_888);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_887) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_2_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_2_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_2_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_2_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_2_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_2_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_2_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_2_bits_data_valid <=
      ~_GEN_1483 & (clear_store ? ~_GEN_1431 & _GEN_920 : ~_GEN_1301 & _GEN_920);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_919) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_2_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_2_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_2_bits_committed <=
      ~_GEN_1459
      & (commit_store_1 ? _GEN_1397 | _GEN_1336 | _GEN_837 : _GEN_1336 | _GEN_837);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_2_bits_succeeded <=
      ~_GEN_1459
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h2
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h2)) & _GEN_821
         & _GEN_677 & stq_2_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_3_valid <=
      ~_GEN_1485 & (clear_store ? ~_GEN_1433 & _GEN_794 : ~_GEN_1302 & _GEN_794);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_3_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678
                ? stq_3_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678
                ? stq_3_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678
                ? stq_3_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_822 & _GEN_678 & stq_3_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h3
         | (_GEN_822
              ? (_GEN_678 ? stq_3_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678
                ? stq_3_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678
                ? stq_3_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_822
           ? (_GEN_678 ? stq_3_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_3_bits_addr_valid <=
      ~_GEN_1485 & (clear_store ? ~_GEN_1433 & _GEN_890 : ~_GEN_1302 & _GEN_890);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_889) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_3_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_3_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_3_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_3_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_3_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_3_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_3_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_3_bits_data_valid <=
      ~_GEN_1485 & (clear_store ? ~_GEN_1433 & _GEN_922 : ~_GEN_1302 & _GEN_922);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_921) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_3_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_3_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_3_bits_committed <=
      ~_GEN_1460
      & (commit_store_1 ? _GEN_1398 | _GEN_1338 | _GEN_838 : _GEN_1338 | _GEN_838);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_3_bits_succeeded <=
      ~_GEN_1460
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h3
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h3)) & _GEN_822
         & _GEN_678 & stq_3_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_4_valid <=
      ~_GEN_1487 & (clear_store ? ~_GEN_1435 & _GEN_796 : ~_GEN_1303 & _GEN_796);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_4_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679
                ? stq_4_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679
                ? stq_4_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679
                ? stq_4_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_823 & _GEN_679 & stq_4_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h4
         | (_GEN_823
              ? (_GEN_679 ? stq_4_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679
                ? stq_4_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679
                ? stq_4_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_823
           ? (_GEN_679 ? stq_4_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_4_bits_addr_valid <=
      ~_GEN_1487 & (clear_store ? ~_GEN_1435 & _GEN_892 : ~_GEN_1303 & _GEN_892);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_891) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_4_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_4_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_4_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_4_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_4_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_4_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_4_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_4_bits_data_valid <=
      ~_GEN_1487 & (clear_store ? ~_GEN_1435 & _GEN_924 : ~_GEN_1303 & _GEN_924);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_923) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_4_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_4_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_4_bits_committed <=
      ~_GEN_1461
      & (commit_store_1 ? _GEN_1399 | _GEN_1340 | _GEN_839 : _GEN_1340 | _GEN_839);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_4_bits_succeeded <=
      ~_GEN_1461
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h4
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h4)) & _GEN_823
         & _GEN_679 & stq_4_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_5_valid <=
      ~_GEN_1489 & (clear_store ? ~_GEN_1437 & _GEN_798 : ~_GEN_1304 & _GEN_798);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_5_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680
                ? stq_5_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680
                ? stq_5_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680
                ? stq_5_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_824 & _GEN_680 & stq_5_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h5
         | (_GEN_824
              ? (_GEN_680 ? stq_5_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680
                ? stq_5_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680
                ? stq_5_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_824
           ? (_GEN_680 ? stq_5_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_5_bits_addr_valid <=
      ~_GEN_1489 & (clear_store ? ~_GEN_1437 & _GEN_894 : ~_GEN_1304 & _GEN_894);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_893) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_5_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_5_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_5_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_5_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_5_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_5_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_5_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_5_bits_data_valid <=
      ~_GEN_1489 & (clear_store ? ~_GEN_1437 & _GEN_926 : ~_GEN_1304 & _GEN_926);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_925) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_5_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_5_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_5_bits_committed <=
      ~_GEN_1462
      & (commit_store_1 ? _GEN_1400 | _GEN_1342 | _GEN_840 : _GEN_1342 | _GEN_840);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_5_bits_succeeded <=
      ~_GEN_1462
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h5
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h5)) & _GEN_824
         & _GEN_680 & stq_5_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_6_valid <=
      ~_GEN_1491 & (clear_store ? ~_GEN_1439 & _GEN_800 : ~_GEN_1305 & _GEN_800);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_6_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681
                ? stq_6_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681
                ? stq_6_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681
                ? stq_6_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_825 & _GEN_681 & stq_6_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h6
         | (_GEN_825
              ? (_GEN_681 ? stq_6_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681
                ? stq_6_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681
                ? stq_6_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_825
           ? (_GEN_681 ? stq_6_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_6_bits_addr_valid <=
      ~_GEN_1491 & (clear_store ? ~_GEN_1439 & _GEN_896 : ~_GEN_1305 & _GEN_896);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_895) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_6_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_6_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_6_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_6_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_6_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_6_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_6_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_6_bits_data_valid <=
      ~_GEN_1491 & (clear_store ? ~_GEN_1439 & _GEN_928 : ~_GEN_1305 & _GEN_928);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_927) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_6_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_6_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_6_bits_committed <=
      ~_GEN_1463
      & (commit_store_1 ? _GEN_1401 | _GEN_1344 | _GEN_841 : _GEN_1344 | _GEN_841);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_6_bits_succeeded <=
      ~_GEN_1463
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h6
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h6)) & _GEN_825
         & _GEN_681 & stq_6_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_7_valid <=
      ~_GEN_1493 & (clear_store ? ~_GEN_1441 & _GEN_802 : ~_GEN_1306 & _GEN_802);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_7_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682
                ? stq_7_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682
                ? stq_7_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682
                ? stq_7_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_826 & _GEN_682 & stq_7_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h7
         | (_GEN_826
              ? (_GEN_682 ? stq_7_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682
                ? stq_7_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682
                ? stq_7_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_826
           ? (_GEN_682 ? stq_7_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_7_bits_addr_valid <=
      ~_GEN_1493 & (clear_store ? ~_GEN_1441 & _GEN_898 : ~_GEN_1306 & _GEN_898);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_897) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_7_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_7_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_7_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_7_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_7_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_7_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_7_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_7_bits_data_valid <=
      ~_GEN_1493 & (clear_store ? ~_GEN_1441 & _GEN_930 : ~_GEN_1306 & _GEN_930);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_929) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_7_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_7_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_7_bits_committed <=
      ~_GEN_1464
      & (commit_store_1 ? _GEN_1402 | _GEN_1346 | _GEN_842 : _GEN_1346 | _GEN_842);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_7_bits_succeeded <=
      ~_GEN_1464
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h7
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h7)) & _GEN_826
         & _GEN_682 & stq_7_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_8_valid <=
      ~_GEN_1495 & (clear_store ? ~_GEN_1443 & _GEN_804 : ~_GEN_1307 & _GEN_804);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_8_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683
                ? stq_8_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683
                ? stq_8_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683
                ? stq_8_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_827 & _GEN_683 & stq_8_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h8
         | (_GEN_827
              ? (_GEN_683 ? stq_8_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683
                ? stq_8_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683
                ? stq_8_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_827
           ? (_GEN_683 ? stq_8_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_8_bits_addr_valid <=
      ~_GEN_1495 & (clear_store ? ~_GEN_1443 & _GEN_900 : ~_GEN_1307 & _GEN_900);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_899) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_8_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_8_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_8_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_8_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_8_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_8_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_8_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_8_bits_data_valid <=
      ~_GEN_1495 & (clear_store ? ~_GEN_1443 & _GEN_932 : ~_GEN_1307 & _GEN_932);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_931) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_8_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_8_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_8_bits_committed <=
      ~_GEN_1465
      & (commit_store_1 ? _GEN_1403 | _GEN_1348 | _GEN_843 : _GEN_1348 | _GEN_843);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_8_bits_succeeded <=
      ~_GEN_1465
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h8
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h8)) & _GEN_827
         & _GEN_683 & stq_8_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_9_valid <=
      ~_GEN_1497 & (clear_store ? ~_GEN_1445 & _GEN_806 : ~_GEN_1308 & _GEN_806);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_9_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684
                ? stq_9_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684
                ? stq_9_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684
                ? stq_9_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_828 & _GEN_684 & stq_9_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'h9
         | (_GEN_828
              ? (_GEN_684 ? stq_9_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684
                ? stq_9_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684
                ? stq_9_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_828
           ? (_GEN_684 ? stq_9_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_9_bits_addr_valid <=
      ~_GEN_1497 & (clear_store ? ~_GEN_1445 & _GEN_902 : ~_GEN_1308 & _GEN_902);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_901) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_9_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_9_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_9_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_9_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_9_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_9_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_9_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_9_bits_data_valid <=
      ~_GEN_1497 & (clear_store ? ~_GEN_1445 & _GEN_934 : ~_GEN_1308 & _GEN_934);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_933) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_9_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_9_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_9_bits_committed <=
      ~_GEN_1466
      & (commit_store_1 ? _GEN_1404 | _GEN_1350 | _GEN_844 : _GEN_1350 | _GEN_844);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_9_bits_succeeded <=
      ~_GEN_1466
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'h9
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'h9)) & _GEN_828
         & _GEN_684 & stq_9_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_10_valid <=
      ~_GEN_1499 & (clear_store ? ~_GEN_1447 & _GEN_808 : ~_GEN_1309 & _GEN_808);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_10_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_ctrl_fcn_dw
                : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_ctrl_is_sta
                : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_ctrl_is_std
                : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_829 & _GEN_685 & stq_10_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'hA
         | (_GEN_829
              ? (_GEN_685 ? stq_10_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_ldst_is_rs1
                : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685
                ? stq_10_bits_uop_bp_debug_if
                : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_829
           ? (_GEN_685 ? stq_10_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_10_bits_addr_valid <=
      ~_GEN_1499 & (clear_store ? ~_GEN_1447 & _GEN_904 : ~_GEN_1309 & _GEN_904);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_903) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_10_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_10_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_10_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_10_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_10_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_10_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_10_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_10_bits_data_valid <=
      ~_GEN_1499 & (clear_store ? ~_GEN_1447 & _GEN_936 : ~_GEN_1309 & _GEN_936);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_935) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_10_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_10_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_10_bits_committed <=
      ~_GEN_1467
      & (commit_store_1 ? _GEN_1405 | _GEN_1352 | _GEN_845 : _GEN_1352 | _GEN_845);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_10_bits_succeeded <=
      ~_GEN_1467
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'hA
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'hA)) & _GEN_829
         & _GEN_685 & stq_10_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_11_valid <=
      ~_GEN_1501 & (clear_store ? ~_GEN_1449 & _GEN_810 : ~_GEN_1310 & _GEN_810);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_11_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_ctrl_fcn_dw
                : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_ctrl_is_sta
                : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_ctrl_is_std
                : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_830 & _GEN_686 & stq_11_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'hB
         | (_GEN_830
              ? (_GEN_686 ? stq_11_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_ldst_is_rs1
                : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686
                ? stq_11_bits_uop_bp_debug_if
                : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_830
           ? (_GEN_686 ? stq_11_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_11_bits_addr_valid <=
      ~_GEN_1501 & (clear_store ? ~_GEN_1449 & _GEN_906 : ~_GEN_1310 & _GEN_906);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_905) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_11_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_11_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_11_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_11_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_11_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_11_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_11_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_11_bits_data_valid <=
      ~_GEN_1501 & (clear_store ? ~_GEN_1449 & _GEN_938 : ~_GEN_1310 & _GEN_938);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_937) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_11_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_11_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_11_bits_committed <=
      ~_GEN_1468
      & (commit_store_1 ? _GEN_1406 | _GEN_1354 | _GEN_846 : _GEN_1354 | _GEN_846);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_11_bits_succeeded <=
      ~_GEN_1468
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'hB
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'hB)) & _GEN_830
         & _GEN_686 & stq_11_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_12_valid <=
      ~_GEN_1503 & (clear_store ? ~_GEN_1451 & _GEN_812 : ~_GEN_1311 & _GEN_812);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_12_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_ctrl_fcn_dw
                : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_ctrl_is_sta
                : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_ctrl_is_std
                : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_831 & _GEN_687 & stq_12_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'hC
         | (_GEN_831
              ? (_GEN_687 ? stq_12_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_ldst_is_rs1
                : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687
                ? stq_12_bits_uop_bp_debug_if
                : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_831
           ? (_GEN_687 ? stq_12_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_12_bits_addr_valid <=
      ~_GEN_1503 & (clear_store ? ~_GEN_1451 & _GEN_908 : ~_GEN_1311 & _GEN_908);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_907) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_12_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_12_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_12_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_12_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_12_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_12_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_12_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_12_bits_data_valid <=
      ~_GEN_1503 & (clear_store ? ~_GEN_1451 & _GEN_940 : ~_GEN_1311 & _GEN_940);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_939) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_12_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_12_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_12_bits_committed <=
      ~_GEN_1469
      & (commit_store_1 ? _GEN_1407 | _GEN_1356 | _GEN_847 : _GEN_1356 | _GEN_847);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_12_bits_succeeded <=
      ~_GEN_1469
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'hC
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'hC)) & _GEN_831
         & _GEN_687 & stq_12_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_13_valid <=
      ~_GEN_1505 & (clear_store ? ~_GEN_1453 & _GEN_814 : ~_GEN_1312 & _GEN_814);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_13_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_ctrl_fcn_dw
                : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_ctrl_is_sta
                : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_ctrl_is_std
                : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_832 & _GEN_688 & stq_13_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'hD
         | (_GEN_832
              ? (_GEN_688 ? stq_13_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_ldst_is_rs1
                : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688
                ? stq_13_bits_uop_bp_debug_if
                : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_832
           ? (_GEN_688 ? stq_13_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_13_bits_addr_valid <=
      ~_GEN_1505 & (clear_store ? ~_GEN_1453 & _GEN_910 : ~_GEN_1312 & _GEN_910);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_909) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_13_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_13_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_13_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_13_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_13_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_13_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_13_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_13_bits_data_valid <=
      ~_GEN_1505 & (clear_store ? ~_GEN_1453 & _GEN_942 : ~_GEN_1312 & _GEN_942);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_941) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_13_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_13_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_13_bits_committed <=
      ~_GEN_1470
      & (commit_store_1 ? _GEN_1408 | _GEN_1358 | _GEN_848 : _GEN_1358 | _GEN_848);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_13_bits_succeeded <=
      ~_GEN_1470
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'hD
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'hD)) & _GEN_832
         & _GEN_688 & stq_13_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_14_valid <=
      ~_GEN_1507 & (clear_store ? ~_GEN_1455 & _GEN_816 : ~_GEN_1313 & _GEN_816);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_14_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_ctrl_fcn_dw
                : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_ctrl_is_sta
                : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_ctrl_is_std
                : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_833 & _GEN_689 & stq_14_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 4'hE
         | (_GEN_833
              ? (_GEN_689 ? stq_14_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :305:44, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_ldst_is_rs1
                : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689
                ? stq_14_bits_uop_bp_debug_if
                : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_833
           ? (_GEN_689 ? stq_14_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_14_bits_addr_valid <=
      ~_GEN_1507 & (clear_store ? ~_GEN_1455 & _GEN_912 : ~_GEN_1313 & _GEN_912);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_911) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_14_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_14_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_14_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_14_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_14_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_14_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_14_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_14_bits_data_valid <=
      ~_GEN_1507 & (clear_store ? ~_GEN_1455 & _GEN_944 : ~_GEN_1313 & _GEN_944);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_943) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_14_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_14_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_14_bits_committed <=
      ~_GEN_1471
      & (commit_store_1 ? _GEN_1409 | _GEN_1360 | _GEN_849 : _GEN_1360 | _GEN_849);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_14_bits_succeeded <=
      ~_GEN_1471
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 4'hE
         | (_GEN_272 | ~(will_fire_store_commit_0 & stq_execute_head == 4'hE)) & _GEN_833
         & _GEN_689 & stq_14_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :305:44, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    stq_15_valid <=
      ~_GEN_1509 & (clear_store ? ~_GEN_1456 & _GEN_818 : ~_GEN_1314 & _GEN_818);	// lsu.scala:211:16, :304:5, :321:5, :1404:5, :1408:7, :1409:32, :1495:3, :1500:17, :1505:3, :1506:35, :1597:3, :1602:5, :1610:32, :1623:9, :1624:34
    stq_15_bits_uop_is_rvc <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc)
           : io_core_dis_uops_1_bits_is_rvc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_fcn_dw <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_ctrl_fcn_dw
                : io_core_dis_uops_0_bits_ctrl_fcn_dw)
           : io_core_dis_uops_1_bits_ctrl_fcn_dw);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_is_load <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_ctrl_is_load
                : io_core_dis_uops_0_bits_ctrl_is_load)
           : io_core_dis_uops_1_bits_ctrl_is_load);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_is_sta <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_ctrl_is_sta
                : io_core_dis_uops_0_bits_ctrl_is_sta)
           : io_core_dis_uops_1_bits_ctrl_is_sta);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ctrl_is_std <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_ctrl_is_std
                : io_core_dis_uops_0_bits_ctrl_is_std)
           : io_core_dis_uops_1_bits_ctrl_is_std);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_iw_p1_poisoned <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_iw_p1_poisoned
                : io_core_dis_uops_0_bits_iw_p1_poisoned)
           : io_core_dis_uops_1_bits_iw_p1_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_iw_p2_poisoned <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_iw_p2_poisoned
                : io_core_dis_uops_0_bits_iw_p2_poisoned)
           : io_core_dis_uops_1_bits_iw_p2_poisoned);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_br <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_br : io_core_dis_uops_0_bits_is_br)
           : io_core_dis_uops_1_bits_is_br);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_jalr <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr)
           : io_core_dis_uops_1_bits_is_jalr);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_jal <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal)
           : io_core_dis_uops_1_bits_is_jal);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_sfb <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb)
           : io_core_dis_uops_1_bits_is_sfb);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_edge_inst <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst)
           : io_core_dis_uops_1_bits_edge_inst);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_taken <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_taken : io_core_dis_uops_0_bits_taken)
           : io_core_dis_uops_1_bits_taken);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_prs1_busy <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy)
           : io_core_dis_uops_1_bits_prs1_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_prs2_busy <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy)
           : io_core_dis_uops_1_bits_prs2_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_prs3_busy <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy)
           : io_core_dis_uops_1_bits_prs3_busy);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ppred_busy <=
      ~_GEN_1477 & _GEN_834 & _GEN_690 & stq_15_bits_uop_ppred_busy;	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_exception <=
      ~_GEN_1477
      & (mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & (&mem_xcpt_uops_0_stq_idx)
         | (_GEN_834
              ? (_GEN_690 ? stq_15_bits_uop_exception : io_core_dis_uops_0_bits_exception)
              : io_core_dis_uops_1_bits_exception));	// lsu.scala:211:16, :304:5, :321:5, :667:32, :671:32, :717:5, :723:7, :728:58, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_bypassable <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable)
           : io_core_dis_uops_1_bits_bypassable);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_mem_signed <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed)
           : io_core_dis_uops_1_bits_mem_signed);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_fence <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence)
           : io_core_dis_uops_1_bits_is_fence);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_fencei <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei)
           : io_core_dis_uops_1_bits_is_fencei);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_amo <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo)
           : io_core_dis_uops_1_bits_is_amo);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_uses_ldq <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq)
           : io_core_dis_uops_1_bits_uses_ldq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_uses_stq <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq)
           : io_core_dis_uops_1_bits_uses_stq);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_sys_pc2epc <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_is_sys_pc2epc
                : io_core_dis_uops_0_bits_is_sys_pc2epc)
           : io_core_dis_uops_1_bits_is_sys_pc2epc);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_is_unique <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique)
           : io_core_dis_uops_1_bits_is_unique);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_flush_on_commit <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_flush_on_commit
                : io_core_dis_uops_0_bits_flush_on_commit)
           : io_core_dis_uops_1_bits_flush_on_commit);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ldst_is_rs1 <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_ldst_is_rs1
                : io_core_dis_uops_0_bits_ldst_is_rs1)
           : io_core_dis_uops_1_bits_ldst_is_rs1);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_ldst_val <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val)
           : io_core_dis_uops_1_bits_ldst_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_frs3_en <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en)
           : io_core_dis_uops_1_bits_frs3_en);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_fp_val <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val)
           : io_core_dis_uops_1_bits_fp_val);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_fp_single <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single)
           : io_core_dis_uops_1_bits_fp_single);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_xcpt_pf_if <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if)
           : io_core_dis_uops_1_bits_xcpt_pf_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_xcpt_ae_if <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if)
           : io_core_dis_uops_1_bits_xcpt_ae_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_xcpt_ma_if <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if)
           : io_core_dis_uops_1_bits_xcpt_ma_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_bp_debug_if <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690
                ? stq_15_bits_uop_bp_debug_if
                : io_core_dis_uops_0_bits_bp_debug_if)
           : io_core_dis_uops_1_bits_bp_debug_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_uop_bp_xcpt_if <=
      ~_GEN_1477
      & (_GEN_834
           ? (_GEN_690 ? stq_15_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if)
           : io_core_dis_uops_1_bits_bp_xcpt_if);	// lsu.scala:211:16, :304:5, :321:5, :1505:3, :1597:3, :1602:5, :1603:16, :1613:32
    stq_15_bits_addr_valid <=
      ~_GEN_1509 & (clear_store ? ~_GEN_1456 & _GEN_914 : ~_GEN_1314 & _GEN_914);	// lsu.scala:211:16, :304:5, :849:5, :853:36, :1404:5, :1408:7, :1409:32, :1410:32, :1495:3, :1500:17, :1505:3, :1506:35, :1507:35, :1597:3, :1602:5, :1610:32, :1611:32, :1623:9, :1624:34, :1625:34
    if (_GEN_913) begin	// lsu.scala:304:5, :849:5, :853:36
      if (exe_tlb_miss_0) begin	// lsu.scala:708:58
        if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
          stq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;	// lsu.scala:211:16
        else if (will_fire_sfence_0)	// lsu.scala:536:61
          stq_15_bits_addr_bits <= _GEN_269;	// lsu.scala:211:16, :610:24
        else if (will_fire_load_retry_0)	// lsu.scala:535:65
          stq_15_bits_addr_bits <= _GEN_191;	// lsu.scala:211:16, :465:79
        else if (will_fire_sta_retry_0)	// lsu.scala:536:61
          stq_15_bits_addr_bits <= _GEN_200;	// lsu.scala:211:16, :478:79
        else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
          stq_15_bits_addr_bits <= hella_req_addr;	// lsu.scala:211:16, :243:34
        else	// lsu.scala:535:65
          stq_15_bits_addr_bits <= 40'h0;	// lsu.scala:211:16
      end
      else	// lsu.scala:708:58
        stq_15_bits_addr_bits <= _GEN_270;	// lsu.scala:211:16, :768:30
      stq_15_bits_addr_is_virtual <= exe_tlb_miss_0;	// lsu.scala:211:16, :708:58
    end
    stq_15_bits_data_valid <=
      ~_GEN_1509 & (clear_store ? ~_GEN_1456 & _GEN_946 : ~_GEN_1314 & _GEN_946);	// lsu.scala:211:16, :304:5, :869:5, :873:33, :1404:5, :1408:7, :1409:32, :1411:32, :1495:3, :1500:17, :1505:3, :1506:35, :1508:35, :1597:3, :1602:5, :1610:32, :1612:32, :1623:9, :1624:34, :1626:34
    if (_GEN_945) begin	// lsu.scala:304:5, :869:5, :873:33
      if (_stq_bits_data_bits_T)	// lsu.scala:868:37
        stq_15_bits_data_bits <= io_core_exe_0_req_bits_data;	// lsu.scala:211:16
      else	// lsu.scala:868:37
        stq_15_bits_data_bits <= io_core_fp_stdata_bits_data;	// lsu.scala:211:16
    end
    stq_15_bits_committed <=
      ~_GEN_1472
      & (commit_store_1 ? (&idx_1) | _GEN_1361 | _GEN_850 : _GEN_1361 | _GEN_850);	// lsu.scala:211:16, :304:5, :321:5, :1306:5, :1451:49, :1453:18, :1455:5, :1456:31, :1505:3, :1509:35, :1510:35
    stq_15_bits_succeeded <=
      ~_GEN_1472
      & (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq
         & io_dmem_resp_0_bits_uop_uses_stq & (&io_dmem_resp_0_bits_uop_stq_idx)
         | (_GEN_272 | ~(will_fire_store_commit_0 & (&stq_execute_head))) & _GEN_834
         & _GEN_690 & stq_15_bits_succeeded);	// lsu.scala:211:16, :220:29, :304:5, :321:5, :535:65, :766:39, :773:43, :780:45, :793:44, :1306:5, :1308:7, :1328:7, :1330:62, :1505:3, :1509:35
    if (_GEN_1476) begin	// lsu.scala:1596:22
      ldq_head <= 4'h0;	// lsu.scala:215:29
      ldq_tail <= 4'h0;	// lsu.scala:216:29
      if (reset)
        stq_tail <= 4'h0;	// lsu.scala:218:29
      else
        stq_tail <= stq_commit_head;	// lsu.scala:218:29, :219:29
    end
    else begin	// lsu.scala:1596:22
      if (commit_load_1)	// lsu.scala:1452:49
        ldq_head <= _GEN_624 + 4'h1;	// lsu.scala:215:29, :305:44, :1486:31, util.scala:203:14
      else if (commit_load)	// lsu.scala:1452:49
        ldq_head <= _GEN_623;	// lsu.scala:215:29, util.scala:203:14
      if (io_core_brupdate_b2_mispredict & ~io_core_exception) begin	// lsu.scala:669:22, :1435:40
        ldq_tail <= io_core_brupdate_b2_uop_ldq_idx;	// lsu.scala:216:29
        stq_tail <= io_core_brupdate_b2_uop_stq_idx;	// lsu.scala:218:29
      end
      else begin	// lsu.scala:1435:40
        if (dis_ld_val_1)	// lsu.scala:301:85
          ldq_tail <= _GEN_100;	// lsu.scala:216:29, util.scala:203:14
        else if (dis_ld_val)	// lsu.scala:301:85
          ldq_tail <= _GEN_95;	// lsu.scala:216:29, util.scala:203:14
        if (dis_st_val_1)	// lsu.scala:302:85
          stq_tail <= _GEN_101;	// lsu.scala:218:29, util.scala:203:14
        else if (dis_st_val)	// lsu.scala:302:85
          stq_tail <= _GEN_96;	// lsu.scala:218:29, util.scala:203:14
      end
    end
    if (_GEN_1474) begin	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
      hella_req_addr <= io_hellacache_req_bits_addr;	// lsu.scala:243:34
      hella_req_cmd <= 5'h0;	// lsu.scala:243:34
      hella_req_size <= 2'h3;	// lsu.scala:243:34
    end
    hella_req_signed <= ~_GEN_1474 & hella_req_signed;	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
    hella_req_phys <= _GEN_1474 | hella_req_phys;	// lsu.scala:243:34, :1527:34, :1529:37, :1530:19
    if (_GEN_1475)	// lsu.scala:244:34, :1527:34, :1533:38
      hella_data_data <= 64'h0;	// AMOALU.scala:26:13, lsu.scala:244:34, :249:20
    if (can_fire_load_incoming_0 | will_fire_load_retry_0 | _GEN_273
        | ~will_fire_hella_incoming_0) begin	// lsu.scala:245:34, :441:63, :535:65, :766:39, :773:43, :780:45, :794:44, :802:47
    end
    else	// lsu.scala:245:34, :766:39, :773:43, :780:45, :794:44, :802:47
      hella_paddr <= exe_tlb_paddr_0;	// Cat.scala:30:58, lsu.scala:245:34
    if (_GEN_1475) begin	// lsu.scala:244:34, :246:34, :1527:34, :1533:38
      hella_xcpt_ma_ld <= _dtlb_io_resp_0_ma_ld;	// lsu.scala:246:34, :249:20
      hella_xcpt_ma_st <= _dtlb_io_resp_0_ma_st;	// lsu.scala:246:34, :249:20
      hella_xcpt_pf_ld <= _dtlb_io_resp_0_pf_ld;	// lsu.scala:246:34, :249:20
      hella_xcpt_pf_st <= _dtlb_io_resp_0_pf_st;	// lsu.scala:246:34, :249:20
      hella_xcpt_ae_ld <= _dtlb_io_resp_0_ae_ld;	// lsu.scala:246:34, :249:20
      hella_xcpt_ae_st <= _dtlb_io_resp_0_ae_st;	// lsu.scala:246:34, :249:20
    end
    if (will_fire_load_wakeup_0) begin	// lsu.scala:535:65
      p1_block_load_mask_0 <= _GEN_208;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_1 <= _GEN_209;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_2 <= _GEN_210;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_3 <= _GEN_211;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_4 <= _GEN_212;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_5 <= _GEN_213;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_6 <= _GEN_214;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_7 <= _GEN_215;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_8 <= _GEN_216;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_9 <= _GEN_217;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_10 <= _GEN_218;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_11 <= _GEN_219;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_12 <= _GEN_220;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_13 <= _GEN_221;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_14 <= _GEN_222;	// lsu.scala:398:35, :570:49
      p1_block_load_mask_15 <= &ldq_wakeup_idx;	// lsu.scala:398:35, :430:31, :570:49
    end
    else if (can_fire_load_incoming_0) begin	// lsu.scala:441:63
      p1_block_load_mask_0 <= _GEN_223;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_1 <= _GEN_224;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_2 <= _GEN_225;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_3 <= _GEN_226;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_4 <= _GEN_227;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_5 <= _GEN_228;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_6 <= _GEN_229;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_7 <= _GEN_230;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_8 <= _GEN_231;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_9 <= _GEN_232;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_10 <= _GEN_233;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_11 <= _GEN_234;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_12 <= _GEN_235;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_13 <= _GEN_236;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_14 <= _GEN_237;	// lsu.scala:398:35, :572:52
      p1_block_load_mask_15 <= &io_core_exe_0_req_bits_uop_ldq_idx;	// lsu.scala:398:35, :572:52
    end
    else begin	// lsu.scala:441:63
      p1_block_load_mask_0 <= _GEN_239;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_1 <= _GEN_241;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_2 <= _GEN_243;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_3 <= _GEN_245;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_4 <= _GEN_247;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_5 <= _GEN_249;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_6 <= _GEN_251;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_7 <= _GEN_253;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_8 <= _GEN_255;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_9 <= _GEN_257;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_10 <= _GEN_259;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_11 <= _GEN_261;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_12 <= _GEN_263;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_13 <= _GEN_265;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_14 <= _GEN_267;	// lsu.scala:398:35, :573:43, :574:49
      p1_block_load_mask_15 <= _GEN_268;	// lsu.scala:398:35, :573:43, :574:49
    end
    p2_block_load_mask_0 <= p1_block_load_mask_0;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_1 <= p1_block_load_mask_1;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_2 <= p1_block_load_mask_2;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_3 <= p1_block_load_mask_3;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_4 <= p1_block_load_mask_4;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_5 <= p1_block_load_mask_5;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_6 <= p1_block_load_mask_6;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_7 <= p1_block_load_mask_7;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_8 <= p1_block_load_mask_8;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_9 <= p1_block_load_mask_9;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_10 <= p1_block_load_mask_10;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_11 <= p1_block_load_mask_11;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_12 <= p1_block_load_mask_12;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_13 <= p1_block_load_mask_13;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_14 <= p1_block_load_mask_14;	// lsu.scala:398:35, :399:35
    p2_block_load_mask_15 <= p1_block_load_mask_15;	// lsu.scala:398:35, :399:35
    _ldq_retry_idx_idx_T_10 =
      _ldq_retry_idx_T_14
        ? 5'h14
        : _ldq_retry_idx_T_17
            ? 5'h15
            : _ldq_retry_idx_T_20
                ? 5'h16
                : _ldq_retry_idx_T_23
                    ? 5'h17
                    : _ldq_retry_idx_T_26
                        ? 5'h18
                        : _ldq_retry_idx_T_29
                            ? 5'h19
                            : _ldq_retry_idx_T_32
                                ? 5'h1A
                                : _ldq_retry_idx_T_35
                                    ? 5'h1B
                                    : _ldq_retry_idx_T_38
                                        ? 5'h1C
                                        : _ldq_retry_idx_T_41
                                            ? 5'h1D
                                            : {4'hF, ~_ldq_retry_idx_T_44};	// Mux.scala:47:69, lsu.scala:305:44, :418:39
    ldq_retry_idx <=
      _ldq_retry_idx_T_2 & _temp_bits_T
        ? 4'h0
        : _ldq_retry_idx_T_5 & _temp_bits_T_2
            ? 4'h1
            : _ldq_retry_idx_T_8 & _temp_bits_T_4
                ? 4'h2
                : _ldq_retry_idx_T_11 & _temp_bits_T_6
                    ? 4'h3
                    : _ldq_retry_idx_T_14 & _temp_bits_T_8
                        ? 4'h4
                        : _ldq_retry_idx_T_17 & _temp_bits_T_10
                            ? 4'h5
                            : _ldq_retry_idx_T_20 & _temp_bits_T_12
                                ? 4'h6
                                : _ldq_retry_idx_T_23 & ~(ldq_head[3])
                                    ? 4'h7
                                    : _ldq_retry_idx_T_26 & _temp_bits_T_16
                                        ? 4'h8
                                        : _ldq_retry_idx_T_29 & _temp_bits_T_18
                                            ? 4'h9
                                            : _ldq_retry_idx_T_32 & _temp_bits_T_20
                                                ? 4'hA
                                                : _ldq_retry_idx_T_35 & _temp_bits_T_22
                                                    ? 4'hB
                                                    : _ldq_retry_idx_T_38
                                                      & _temp_bits_T_24
                                                        ? 4'hC
                                                        : _ldq_retry_idx_T_41
                                                          & _temp_bits_T_26
                                                            ? 4'hD
                                                            : _ldq_retry_idx_T_44
                                                              & _temp_bits_T_28
                                                                ? 4'hE
                                                                : ldq_15_bits_addr_valid
                                                                  & ldq_15_bits_addr_is_virtual
                                                                  & ~ldq_retry_idx_block_15
                                                                    ? 4'hF
                                                                    : _ldq_retry_idx_T_2
                                                                        ? 4'h0
                                                                        : _ldq_retry_idx_T_5
                                                                            ? 4'h1
                                                                            : _ldq_retry_idx_T_8
                                                                                ? 4'h2
                                                                                : _ldq_retry_idx_T_11
                                                                                    ? 4'h3
                                                                                    : _ldq_retry_idx_idx_T_10[3:0];	// Mux.scala:47:69, lsu.scala:210:16, :215:29, :305:44, :415:30, :417:36, :418:{39,42}, util.scala:351:{65,72}
    _stq_retry_idx_idx_T_10 =
      _stq_retry_idx_T_4
        ? 5'h14
        : _stq_retry_idx_T_5
            ? 5'h15
            : _stq_retry_idx_T_6
                ? 5'h16
                : _stq_retry_idx_T_7
                    ? 5'h17
                    : _stq_retry_idx_T_8
                        ? 5'h18
                        : _stq_retry_idx_T_9
                            ? 5'h19
                            : _stq_retry_idx_T_10
                                ? 5'h1A
                                : _stq_retry_idx_T_11
                                    ? 5'h1B
                                    : _stq_retry_idx_T_12
                                        ? 5'h1C
                                        : _stq_retry_idx_T_13
                                            ? 5'h1D
                                            : {4'hF, ~_stq_retry_idx_T_14};	// Mux.scala:47:69, lsu.scala:305:44, :424:18
    stq_retry_idx <=
      _stq_retry_idx_T & stq_commit_head == 4'h0
        ? 4'h0
        : _stq_retry_idx_T_1 & stq_commit_head < 4'h2
            ? 4'h1
            : _stq_retry_idx_T_2 & stq_commit_head < 4'h3
                ? 4'h2
                : _stq_retry_idx_T_3 & stq_commit_head < 4'h4
                    ? 4'h3
                    : _stq_retry_idx_T_4 & stq_commit_head < 4'h5
                        ? 4'h4
                        : _stq_retry_idx_T_5 & stq_commit_head < 4'h6
                            ? 4'h5
                            : _stq_retry_idx_T_6 & stq_commit_head < 4'h7
                                ? 4'h6
                                : _stq_retry_idx_T_7 & ~(stq_commit_head[3])
                                    ? 4'h7
                                    : _stq_retry_idx_T_8 & stq_commit_head < 4'h9
                                        ? 4'h8
                                        : _stq_retry_idx_T_9 & stq_commit_head < 4'hA
                                            ? 4'h9
                                            : _stq_retry_idx_T_10 & stq_commit_head < 4'hB
                                                ? 4'hA
                                                : _stq_retry_idx_T_11
                                                  & stq_commit_head[3:2] != 2'h3
                                                    ? 4'hB
                                                    : _stq_retry_idx_T_12
                                                      & stq_commit_head < 4'hD
                                                        ? 4'hC
                                                        : _stq_retry_idx_T_13
                                                          & stq_commit_head[3:1] != 3'h7
                                                            ? 4'hD
                                                            : _stq_retry_idx_T_14
                                                              & stq_commit_head != 4'hF
                                                                ? 4'hE
                                                                : stq_15_bits_addr_valid
                                                                  & stq_15_bits_addr_is_virtual
                                                                    ? 4'hF
                                                                    : _stq_retry_idx_T
                                                                        ? 4'h0
                                                                        : _stq_retry_idx_T_1
                                                                            ? 4'h1
                                                                            : _stq_retry_idx_T_2
                                                                                ? 4'h2
                                                                                : _stq_retry_idx_T_3
                                                                                    ? 4'h3
                                                                                    : _stq_retry_idx_idx_T_10[3:0];	// Mux.scala:47:69, lsu.scala:211:16, :219:29, :305:44, :422:30, :424:18, util.scala:351:{65,72}
    _ldq_wakeup_idx_idx_T_10 =
      _ldq_wakeup_idx_T_39
        ? 5'h14
        : _ldq_wakeup_idx_T_47
            ? 5'h15
            : _ldq_wakeup_idx_T_55
                ? 5'h16
                : _ldq_wakeup_idx_T_63
                    ? 5'h17
                    : _ldq_wakeup_idx_T_71
                        ? 5'h18
                        : _ldq_wakeup_idx_T_79
                            ? 5'h19
                            : _ldq_wakeup_idx_T_87
                                ? 5'h1A
                                : _ldq_wakeup_idx_T_95
                                    ? 5'h1B
                                    : _ldq_wakeup_idx_T_103
                                        ? 5'h1C
                                        : _ldq_wakeup_idx_T_111
                                            ? 5'h1D
                                            : {4'hF, ~_ldq_wakeup_idx_T_119};	// Mux.scala:47:69, lsu.scala:305:44, :433:71
    ldq_wakeup_idx <=
      _ldq_wakeup_idx_T_7 & _temp_bits_T
        ? 4'h0
        : _ldq_wakeup_idx_T_15 & _temp_bits_T_2
            ? 4'h1
            : _ldq_wakeup_idx_T_23 & _temp_bits_T_4
                ? 4'h2
                : _ldq_wakeup_idx_T_31 & _temp_bits_T_6
                    ? 4'h3
                    : _ldq_wakeup_idx_T_39 & _temp_bits_T_8
                        ? 4'h4
                        : _ldq_wakeup_idx_T_47 & _temp_bits_T_10
                            ? 4'h5
                            : _ldq_wakeup_idx_T_55 & _temp_bits_T_12
                                ? 4'h6
                                : _ldq_wakeup_idx_T_63 & ~(ldq_head[3])
                                    ? 4'h7
                                    : _ldq_wakeup_idx_T_71 & _temp_bits_T_16
                                        ? 4'h8
                                        : _ldq_wakeup_idx_T_79 & _temp_bits_T_18
                                            ? 4'h9
                                            : _ldq_wakeup_idx_T_87 & _temp_bits_T_20
                                                ? 4'hA
                                                : _ldq_wakeup_idx_T_95 & _temp_bits_T_22
                                                    ? 4'hB
                                                    : _ldq_wakeup_idx_T_103
                                                      & _temp_bits_T_24
                                                        ? 4'hC
                                                        : _ldq_wakeup_idx_T_111
                                                          & _temp_bits_T_26
                                                            ? 4'hD
                                                            : _ldq_wakeup_idx_T_119
                                                              & _temp_bits_T_28
                                                                ? 4'hE
                                                                : ldq_15_bits_addr_valid
                                                                  & ~ldq_15_bits_executed
                                                                  & ~ldq_15_bits_succeeded
                                                                  & ~ldq_15_bits_addr_is_virtual
                                                                  & ~ldq_retry_idx_block_15
                                                                    ? 4'hF
                                                                    : _ldq_wakeup_idx_T_7
                                                                        ? 4'h0
                                                                        : _ldq_wakeup_idx_T_15
                                                                            ? 4'h1
                                                                            : _ldq_wakeup_idx_T_23
                                                                                ? 4'h2
                                                                                : _ldq_wakeup_idx_T_31
                                                                                    ? 4'h3
                                                                                    : _ldq_wakeup_idx_idx_T_10[3:0];	// Mux.scala:47:69, lsu.scala:210:16, :215:29, :305:44, :417:36, :430:31, :433:{21,36,52,71,74}, util.scala:351:{65,72}
    can_fire_load_retry_REG <= _dtlb_io_miss_rdy;	// lsu.scala:249:20, :470:40
    can_fire_sta_retry_REG <= _dtlb_io_miss_rdy;	// lsu.scala:249:20, :482:41
    mem_xcpt_valids_0 <=
      (pf_ld_0 | pf_st_0 | ae_ld_0 | ~_will_fire_store_commit_0_T_2
       & _dtlb_io_resp_0_ae_st & _mem_xcpt_uops_WIRE_0_uses_stq | ma_ld_0 | ma_st_0)
      & ~io_core_exception
      & (io_core_brupdate_b1_mispredict_mask & exe_tlb_uop_0_br_mask) == 12'h0;	// lsu.scala:249:20, :538:31, :576:25, :597:24, :659:56, :660:87, :661:75, :662:75, :663:75, :664:75, :667:32, :668:80, :669:{22,41}, util.scala:118:{51,59}
    mem_xcpt_uops_0_br_mask <= exe_tlb_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:597:24, :671:32, util.scala:85:{25,27}
    if (_exe_tlb_uop_T_2) begin	// lsu.scala:599:53
      mem_xcpt_uops_0_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;	// lsu.scala:671:32
      mem_xcpt_uops_0_ldq_idx <= io_core_exe_0_req_bits_uop_ldq_idx;	// lsu.scala:671:32
      mem_xcpt_uops_0_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;	// lsu.scala:671:32
      mem_xcpt_uops_0_uses_ldq <= io_core_exe_0_req_bits_uop_uses_ldq;	// lsu.scala:671:32
      mem_xcpt_uops_0_uses_stq <= io_core_exe_0_req_bits_uop_uses_stq;	// lsu.scala:671:32
    end
    else if (will_fire_load_retry_0) begin	// lsu.scala:535:65
      mem_xcpt_uops_0_rob_idx <= _GEN_141;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_ldq_idx <= _GEN_143;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_stq_idx <= mem_ldq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_uses_ldq <= _GEN_165;	// lsu.scala:465:79, :671:32
      mem_xcpt_uops_0_uses_stq <= _GEN_167;	// lsu.scala:465:79, :671:32
    end
    else begin	// lsu.scala:535:65
      if (will_fire_sta_retry_0) begin	// lsu.scala:536:61
        mem_xcpt_uops_0_rob_idx <= mem_stq_retry_e_out_bits_uop_rob_idx;	// lsu.scala:478:79, :671:32
        mem_xcpt_uops_0_ldq_idx <= _GEN_198;	// lsu.scala:478:79, :671:32
        mem_xcpt_uops_0_stq_idx <= mem_stq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:478:79, :671:32
      end
      else begin	// lsu.scala:536:61
        mem_xcpt_uops_0_rob_idx <= 6'h0;	// lsu.scala:671:32
        mem_xcpt_uops_0_ldq_idx <= 4'h0;	// lsu.scala:671:32
        mem_xcpt_uops_0_stq_idx <= 4'h0;	// lsu.scala:671:32
      end
      mem_xcpt_uops_0_uses_ldq <= _exe_tlb_uop_T_4_uses_ldq;	// lsu.scala:602:24, :671:32
      mem_xcpt_uops_0_uses_stq <= _exe_tlb_uop_T_4_uses_stq;	// lsu.scala:602:24, :671:32
    end
    if (ma_ld_0)	// lsu.scala:659:56
      mem_xcpt_causes_0 <= 4'h4;	// lsu.scala:305:44, :672:32
    else if (ma_st_0)	// lsu.scala:660:87
      mem_xcpt_causes_0 <= 4'h6;	// lsu.scala:305:44, :672:32
    else if (pf_ld_0)	// lsu.scala:661:75
      mem_xcpt_causes_0 <= 4'hD;	// lsu.scala:305:44, :672:32
    else if (pf_st_0)	// lsu.scala:662:75
      mem_xcpt_causes_0 <= 4'hF;	// lsu.scala:305:44, :672:32
    else	// lsu.scala:662:75
      mem_xcpt_causes_0 <= {2'h1, ~ae_ld_0, 1'h1};	// lsu.scala:249:20, :663:75, :672:32, :676:8, :677:8, :1312:58
    if (_exe_tlb_vaddr_T_1)	// lsu.scala:608:53
      mem_xcpt_vaddrs_0 <= io_core_exe_0_req_bits_addr;	// lsu.scala:679:32
    else if (will_fire_sfence_0)	// lsu.scala:536:61
      mem_xcpt_vaddrs_0 <= _GEN_269;	// lsu.scala:610:24, :679:32
    else if (will_fire_load_retry_0)	// lsu.scala:535:65
      mem_xcpt_vaddrs_0 <= _GEN_191;	// lsu.scala:465:79, :679:32
    else if (will_fire_sta_retry_0)	// lsu.scala:536:61
      mem_xcpt_vaddrs_0 <= _GEN_200;	// lsu.scala:478:79, :679:32
    else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
      mem_xcpt_vaddrs_0 <= hella_req_addr;	// lsu.scala:243:34, :679:32
    else	// lsu.scala:535:65
      mem_xcpt_vaddrs_0 <= 40'h0;	// lsu.scala:679:32
    REG <= _GEN_207 | will_fire_load_retry_0 | will_fire_sta_retry_0;	// lsu.scala:535:65, :536:61, :567:93, :718:21, :719:33
    fired_load_incoming_REG <= can_fire_load_incoming_0 & _fired_std_incoming_T;	// lsu.scala:441:63, :894:{51,79}, util.scala:118:59
    fired_stad_incoming_REG <= will_fire_stad_incoming_0 & _fired_std_incoming_T;	// lsu.scala:534:63, :895:{51,79}, util.scala:118:59
    fired_sta_incoming_REG <= will_fire_sta_incoming_0 & _fired_std_incoming_T;	// lsu.scala:536:61, :896:{51,79}, util.scala:118:59
    fired_std_incoming_REG <= will_fire_std_incoming_0 & _fired_std_incoming_T;	// lsu.scala:536:61, :897:{51,79}, util.scala:118:59
    fired_stdf_incoming <=
      fp_stdata_fire
      & (io_core_brupdate_b1_mispredict_mask
         & io_core_fp_stdata_bits_uop_br_mask) == 12'h0;	// Decoupled.scala:40:37, lsu.scala:898:{37,62}, util.scala:118:{51,59}
    fired_sfence_0 <= will_fire_sfence_0;	// lsu.scala:536:61, :899:37
    fired_release_0 <= will_fire_release_0;	// lsu.scala:534:63, :900:37
    fired_load_retry_REG <=
      will_fire_load_retry_0 & (io_core_brupdate_b1_mispredict_mask & _GEN_132) == 12'h0;	// lsu.scala:465:79, :535:65, :901:{51,79}, util.scala:118:{51,59}
    fired_sta_retry_REG <= will_fire_sta_retry_0 & _mem_stq_retry_e_out_valid_T == 12'h0;	// lsu.scala:536:61, :902:{51,79}, util.scala:118:{51,59}
    fired_load_wakeup_REG <=
      will_fire_load_wakeup_0 & (io_core_brupdate_b1_mispredict_mask & _GEN_201) == 12'h0;	// lsu.scala:502:88, :535:65, :904:{51,79}, util.scala:118:{51,59}
    mem_incoming_uop_0_br_mask <=
      io_core_exe_0_req_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:908:37, util.scala:85:{25,27}
    mem_incoming_uop_0_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;	// lsu.scala:908:37
    mem_incoming_uop_0_ldq_idx <= io_core_exe_0_req_bits_uop_ldq_idx;	// lsu.scala:908:37
    mem_incoming_uop_0_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;	// lsu.scala:908:37
    mem_incoming_uop_0_pdst <= io_core_exe_0_req_bits_uop_pdst;	// lsu.scala:908:37
    mem_incoming_uop_0_fp_val <= io_core_exe_0_req_bits_uop_fp_val;	// lsu.scala:908:37
    mem_ldq_incoming_e_0_bits_uop_br_mask <=
      _GEN_102[io_core_exe_0_req_bits_uop_ldq_idx] & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:264:49, :909:37, util.scala:85:27, :89:21
    mem_ldq_incoming_e_0_bits_uop_stq_idx <= _GEN_103[io_core_exe_0_req_bits_uop_ldq_idx];	// lsu.scala:264:49, :909:37
    mem_ldq_incoming_e_0_bits_uop_mem_size <=
      _GEN_104[io_core_exe_0_req_bits_uop_ldq_idx];	// lsu.scala:264:49, :909:37
    mem_ldq_incoming_e_0_bits_st_dep_mask <= _GEN_107[io_core_exe_0_req_bits_uop_ldq_idx];	// lsu.scala:264:49, :909:37
    mem_stq_incoming_e_0_valid <=
      _GEN_2[io_core_exe_0_req_bits_uop_stq_idx]
      & (io_core_brupdate_b1_mispredict_mask
         & _GEN_28[io_core_exe_0_req_bits_uop_stq_idx]) == 12'h0;	// lsu.scala:224:42, :264:49, :910:37, util.scala:108:31, :118:{51,59}
    mem_stq_incoming_e_0_bits_uop_br_mask <=
      _GEN_28[io_core_exe_0_req_bits_uop_stq_idx] & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:224:42, :264:49, :910:37, util.scala:85:27, :89:21
    mem_stq_incoming_e_0_bits_uop_rob_idx <= _GEN_36[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_uop_stq_idx <= _GEN_38[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_uop_mem_size <= _GEN_55[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_uop_is_amo <= _GEN_61[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_addr_valid <= _GEN_87[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_addr_is_virtual <=
      _GEN_90[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_stq_incoming_e_0_bits_data_valid <= _GEN_91[io_core_exe_0_req_bits_uop_stq_idx];	// lsu.scala:224:42, :264:49, :910:37
    mem_ldq_wakeup_e_bits_uop_br_mask <= _GEN_201 & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:502:88, :911:37, util.scala:85:27, :89:21
    mem_ldq_wakeup_e_bits_uop_stq_idx <= mem_ldq_wakeup_e_out_bits_uop_stq_idx;	// lsu.scala:502:88, :911:37
    mem_ldq_wakeup_e_bits_uop_mem_size <= mem_ldq_wakeup_e_out_bits_uop_mem_size;	// lsu.scala:502:88, :911:37
    mem_ldq_wakeup_e_bits_st_dep_mask <= mem_ldq_wakeup_e_out_bits_st_dep_mask;	// lsu.scala:502:88, :911:37
    mem_ldq_retry_e_bits_uop_br_mask <= _GEN_132 & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:465:79, :912:37, util.scala:85:27, :89:21
    mem_ldq_retry_e_bits_uop_stq_idx <= mem_ldq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:465:79, :912:37
    mem_ldq_retry_e_bits_uop_mem_size <= mem_ldq_retry_e_out_bits_uop_mem_size;	// lsu.scala:465:79, :912:37
    mem_ldq_retry_e_bits_st_dep_mask <= _GEN_107[ldq_retry_idx];	// lsu.scala:264:49, :415:30, :465:79, :912:37
    mem_stq_retry_e_valid <= _GEN_196 & _mem_stq_retry_e_out_valid_T == 12'h0;	// lsu.scala:478:79, :913:37, util.scala:108:31, :118:{51,59}
    mem_stq_retry_e_bits_uop_br_mask <= _GEN_197 & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:478:79, :913:37, util.scala:85:27, :89:21
    mem_stq_retry_e_bits_uop_rob_idx <= mem_stq_retry_e_out_bits_uop_rob_idx;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_uop_stq_idx <= mem_stq_retry_e_out_bits_uop_stq_idx;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_uop_mem_size <= mem_stq_retry_e_out_bits_uop_mem_size;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_uop_is_amo <= mem_stq_retry_e_out_bits_uop_is_amo;	// lsu.scala:478:79, :913:37
    mem_stq_retry_e_bits_data_valid <= _GEN_91[stq_retry_idx];	// lsu.scala:224:42, :422:30, :478:79, :913:37
    mem_stdf_uop_br_mask <=
      io_core_fp_stdata_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:922:37, util.scala:85:{25,27}
    mem_stdf_uop_rob_idx <= io_core_fp_stdata_bits_uop_rob_idx;	// lsu.scala:922:37
    mem_stdf_uop_stq_idx <= io_core_fp_stdata_bits_uop_stq_idx;	// lsu.scala:922:37
    mem_tlb_miss_0 <= exe_tlb_miss_0;	// lsu.scala:708:58, :925:41
    mem_tlb_uncacheable_0 <= ~_dtlb_io_resp_0_cacheable;	// lsu.scala:249:20, :711:43, :926:41
    if (_GEN_275)	// lsu.scala:766:39, :768:30, :773:43
      mem_paddr_0 <= _GEN_270;	// lsu.scala:768:30, :927:41
    else if (will_fire_store_commit_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_89;	// lsu.scala:224:42, :927:41
    else if (will_fire_load_wakeup_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_202;	// lsu.scala:502:88, :927:41
    else if (will_fire_hella_incoming_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_270;	// lsu.scala:768:30, :927:41
    else if (will_fire_hella_wakeup_0)	// lsu.scala:535:65
      mem_paddr_0 <= _GEN_274;	// lsu.scala:822:39, :927:41
    else	// lsu.scala:535:65
      mem_paddr_0 <= 40'h0;	// lsu.scala:927:41
    if (fired_stad_incoming_REG | fired_sta_incoming_REG | fired_std_incoming_REG)	// lsu.scala:895:51, :896:51, :897:51, :940:35, :945:27, :947:41, :953:27, :955:41, :961:27, :963:35
      clr_bsy_rob_idx_0 <= mem_stq_incoming_e_0_bits_uop_rob_idx;	// lsu.scala:910:37, :931:28
    else if (fired_sfence_0)	// lsu.scala:899:37
      clr_bsy_rob_idx_0 <= mem_incoming_uop_0_rob_idx;	// lsu.scala:908:37, :931:28
    else if (fired_sta_retry_REG)	// lsu.scala:902:51
      clr_bsy_rob_idx_0 <= mem_stq_retry_e_bits_uop_rob_idx;	// lsu.scala:913:37, :931:28
    else	// lsu.scala:902:51
      clr_bsy_rob_idx_0 <= 6'h0;	// lsu.scala:931:28
    if (fired_stad_incoming_REG)	// lsu.scala:895:51
      clr_bsy_brmask_0 <=
        mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:910:37, :932:28, util.scala:85:{25,27}
    else if (fired_sta_incoming_REG)	// lsu.scala:896:51
      clr_bsy_brmask_0 <=
        mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:910:37, :932:28, util.scala:85:{25,27}
    else if (fired_std_incoming_REG)	// lsu.scala:897:51
      clr_bsy_brmask_0 <=
        mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:910:37, :932:28, util.scala:85:{25,27}
    else if (fired_sfence_0)	// lsu.scala:899:37
      clr_bsy_brmask_0 <= mem_incoming_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:908:37, :932:28, util.scala:85:{25,27}
    else if (fired_sta_retry_REG)	// lsu.scala:902:51
      clr_bsy_brmask_0 <=
        mem_stq_retry_e_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:913:37, :932:28, util.scala:85:{25,27}
    else	// lsu.scala:902:51
      clr_bsy_brmask_0 <= 12'h0;	// lsu.scala:932:28
    io_core_clr_bsy_0_valid_REG <= io_core_exception;	// lsu.scala:979:62
    io_core_clr_bsy_0_valid_REG_1 <= io_core_exception;	// lsu.scala:979:101
    io_core_clr_bsy_0_valid_REG_2 <= io_core_clr_bsy_0_valid_REG_1;	// lsu.scala:979:{93,101}
    if (fired_stdf_incoming) begin	// lsu.scala:898:37
      stdf_clr_bsy_rob_idx <= mem_stdf_uop_rob_idx;	// lsu.scala:922:37, :984:33
      stdf_clr_bsy_brmask <= mem_stdf_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:922:37, :985:33, util.scala:85:{25,27}
    end
    else begin	// lsu.scala:898:37
      stdf_clr_bsy_rob_idx <= 6'h0;	// lsu.scala:984:33
      stdf_clr_bsy_brmask <= 12'h0;	// lsu.scala:985:33
    end
    io_core_clr_bsy_1_valid_REG <= io_core_exception;	// lsu.scala:1004:67
    io_core_clr_bsy_1_valid_REG_1 <= io_core_exception;	// lsu.scala:1004:106
    io_core_clr_bsy_1_valid_REG_2 <= io_core_clr_bsy_1_valid_REG_1;	// lsu.scala:1004:{98,106}
    lcam_addr_REG <= exe_tlb_paddr_0;	// Cat.scala:30:58, lsu.scala:1026:45
    lcam_addr_REG_1 <= io_dmem_release_bits_address;	// lsu.scala:1027:67
    lcam_ldq_idx_REG <= ldq_wakeup_idx;	// lsu.scala:430:31, :1037:58
    lcam_ldq_idx_REG_1 <= ldq_retry_idx;	// lsu.scala:415:30, :1038:58
    lcam_stq_idx_REG <= stq_retry_idx;	// lsu.scala:422:30, :1042:58
    if (can_fire_load_incoming_0) begin	// lsu.scala:441:63
      s1_executing_loads_0 <= _GEN_223 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_1 <= _GEN_224 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_2 <= _GEN_225 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_3 <= _GEN_226 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_4 <= _GEN_227 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_5 <= _GEN_228 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_6 <= _GEN_229 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_7 <= _GEN_230 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_8 <= _GEN_231 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_9 <= _GEN_232 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_10 <= _GEN_233 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_11 <= _GEN_234 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_12 <= _GEN_235 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_13 <= _GEN_236 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_14 <= _GEN_237 & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
      s1_executing_loads_15 <= (&io_core_exe_0_req_bits_uop_ldq_idx) & dmem_req_fire_0;	// lsu.scala:572:52, :752:55, :771:47, :1056:35
    end
    else if (will_fire_load_retry_0) begin	// lsu.scala:535:65
      s1_executing_loads_0 <= _GEN_238 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_1 <= _GEN_240 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_2 <= _GEN_242 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_3 <= _GEN_244 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_4 <= _GEN_246 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_5 <= _GEN_248 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_6 <= _GEN_250 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_7 <= _GEN_252 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_8 <= _GEN_254 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_9 <= _GEN_256 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_10 <= _GEN_258 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_11 <= _GEN_260 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_12 <= _GEN_262 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_13 <= _GEN_264 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_14 <= _GEN_266 & dmem_req_fire_0;	// lsu.scala:574:49, :752:55, :778:41, :1056:35
      s1_executing_loads_15 <= (&ldq_retry_idx) & dmem_req_fire_0;	// lsu.scala:415:30, :574:49, :752:55, :778:41, :1056:35
    end
    else begin	// lsu.scala:535:65
      s1_executing_loads_0 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_208 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_1 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_209 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_2 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_210 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_3 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_211 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_4 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_212 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_5 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_213 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_6 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_214 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_7 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_215 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_8 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_216 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_9 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_217 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_10 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_218 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_11 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_219 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_12 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_220 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_13 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_221 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_14 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & _GEN_222 & dmem_req_fire_0;	// lsu.scala:535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
      s1_executing_loads_15 <=
        ~will_fire_store_commit_0 & will_fire_load_wakeup_0 & (&ldq_wakeup_idx)
        & dmem_req_fire_0;	// lsu.scala:430:31, :535:65, :570:49, :752:55, :780:45, :794:44, :1056:35
    end
    wb_forward_valid_0 <= mem_forward_valid_0;	// lsu.scala:1064:36, :1189:53
    if (fired_load_incoming_REG)	// lsu.scala:894:51
      wb_forward_ldq_idx_0 <= mem_incoming_uop_0_ldq_idx;	// lsu.scala:908:37, :1065:36
    else if (fired_load_wakeup_REG)	// lsu.scala:904:51
      wb_forward_ldq_idx_0 <= lcam_ldq_idx_REG;	// lsu.scala:1037:58, :1065:36
    else if (fired_load_retry_REG)	// lsu.scala:901:51
      wb_forward_ldq_idx_0 <= lcam_ldq_idx_REG_1;	// lsu.scala:1038:58, :1065:36
    else	// lsu.scala:901:51
      wb_forward_ldq_idx_0 <= 4'h0;	// lsu.scala:1065:36
    if (_lcam_addr_T_1)	// lsu.scala:1025:86
      wb_forward_ld_addr_0 <= _GEN_281;	// lsu.scala:1025:37, :1066:36
    else if (fired_release_0)	// lsu.scala:900:37
      wb_forward_ld_addr_0 <= _GEN_280;	// lsu.scala:1027:41, :1066:36
    else	// lsu.scala:900:37
      wb_forward_ld_addr_0 <= mem_paddr_0;	// lsu.scala:927:41, :1066:36
    wb_forward_stq_idx_0 <= _forwarding_age_logic_0_io_forwarding_idx;	// lsu.scala:1067:36, :1178:57
    older_nacked_REG <= nacking_loads_0;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_1 <= nacking_loads_1;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_1 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_2 <= nacking_loads_2;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_2 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_3 <= nacking_loads_3;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_3 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_4 <= nacking_loads_4;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_4 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_5 <= nacking_loads_5;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_5 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_6 <= nacking_loads_6;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_6 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_7 <= nacking_loads_7;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_7 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_8 <= nacking_loads_8;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_8 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_9 <= nacking_loads_9;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_9 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_10 <= nacking_loads_10;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_10 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_11 <= nacking_loads_11;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_11 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_12 <= nacking_loads_12;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_12 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_13 <= nacking_loads_13;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_13 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_14 <= nacking_loads_14;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_14 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    older_nacked_REG_15 <= nacking_loads_15;	// lsu.scala:1128:57, :1284:5, :1287:7
    io_dmem_s1_kill_0_REG_15 <= dmem_req_fire_0;	// lsu.scala:752:55, :1131:58
    io_dmem_s1_kill_0_REG_16 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_17 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_18 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_19 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_20 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_21 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_22 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_23 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_24 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_25 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_26 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_27 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_28 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_29 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_30 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_31 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_32 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_33 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_34 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_35 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_36 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_37 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_38 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_39 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_40 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_41 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_42 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_43 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_44 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_45 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_46 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_47 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_48 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_49 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_50 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_51 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_52 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_53 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_54 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_55 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_56 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_57 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_58 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_59 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_60 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    io_dmem_s1_kill_0_REG_61 <= dmem_req_fire_0;	// lsu.scala:752:55, :1153:56
    io_dmem_s1_kill_0_REG_62 <= dmem_req_fire_0;	// lsu.scala:752:55, :1159:56
    io_dmem_s1_kill_0_REG_63 <= dmem_req_fire_0;	// lsu.scala:752:55, :1165:56
    REG_1 <= io_core_exception;	// lsu.scala:1189:64
    REG_2 <=
      (ldst_addr_matches_0_0 | ldst_addr_matches_0_1 | ldst_addr_matches_0_2
       | ldst_addr_matches_0_3 | ldst_addr_matches_0_4 | ldst_addr_matches_0_5
       | ldst_addr_matches_0_6 | ldst_addr_matches_0_7 | ldst_addr_matches_0_8
       | ldst_addr_matches_0_9 | ldst_addr_matches_0_10 | ldst_addr_matches_0_11
       | ldst_addr_matches_0_12 | ldst_addr_matches_0_13 | ldst_addr_matches_0_14
       | ldst_addr_matches_0_15) & ~mem_forward_valid_0;	// lsu.scala:1148:72, :1150:9, :1189:53, :1199:{18,48,53,56}
    if (will_fire_store_commit_0 | ~can_fire_store_commit_0)	// lsu.scala:493:79, :535:65, :1205:{37,40}
      store_blocked_counter <= 4'h0;	// lsu.scala:1204:36
    else if (can_fire_store_commit_0 & ~will_fire_store_commit_0) begin	// lsu.scala:493:79, :535:65, :584:6, :1207:43
      if (&store_blocked_counter)	// lsu.scala:1204:36, :1208:58
        store_blocked_counter <= store_blocked_counter + 4'h1;	// lsu.scala:305:44, :1204:36, :1208:90
      else	// lsu.scala:1208:58
        store_blocked_counter <= 4'hF;	// lsu.scala:305:44, :1204:36
    end
    r_xcpt_uop_br_mask <= xcpt_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;	// lsu.scala:1236:25, :1243:21, util.scala:85:{25,27}
    if (use_mem_xcpt) begin	// lsu.scala:1241:115
      r_xcpt_uop_rob_idx <= mem_xcpt_uops_0_rob_idx;	// lsu.scala:671:32, :1236:25
      r_xcpt_cause <= {1'h0, mem_xcpt_causes_0};	// lsu.scala:249:20, :672:32, :708:86, :1236:25, :1250:28
    end
    else begin	// lsu.scala:1241:115
      r_xcpt_uop_rob_idx <= _GEN_140[l_idx];	// Mux.scala:47:69, lsu.scala:465:79, :1236:25, util.scala:363:52
      r_xcpt_cause <= 5'h10;	// Mux.scala:47:69, lsu.scala:1236:25
    end
    r_xcpt_badvaddr <= mem_xcpt_vaddrs_0;	// lsu.scala:679:32, :1236:25
    io_core_ld_miss_REG <= _io_core_spec_ld_wakeup_0_valid_output;	// lsu.scala:1260:69, :1380:37
    spec_ld_succeed_REG <= _io_core_spec_ld_wakeup_0_valid_output;	// lsu.scala:1260:69, :1382:13
    spec_ld_succeed_REG_1 <= mem_incoming_uop_0_ldq_idx;	// lsu.scala:908:37, :1384:56
    if (reset) begin
      hella_state <= 3'h0;	// lsu.scala:242:38
      live_store_mask <= 16'h0;	// lsu.scala:259:32
      clr_bsy_valid_0 <= 1'h0;	// lsu.scala:249:20, :708:86, :930:32
      stdf_clr_bsy_valid <= 1'h0;	// lsu.scala:249:20, :708:86, :983:37
      r_xcpt_valid <= 1'h0;	// lsu.scala:249:20, :708:86, :1235:29
    end
    else begin
      if (|hella_state) begin	// lsu.scala:242:38, :593:24
        automatic logic            _GEN_1510;	// lsu.scala:1540:50
        automatic logic [2:0]      _GEN_1511;	// lsu.scala:242:38, :1582:40, :1584:69, :1585:21
        automatic logic [7:0][2:0] _GEN_1512;	// lsu.scala:803:26, :820:26, :1288:28, :1533:38, :1539:34, :1550:{28,43}, :1552:17, :1553:{28,38}, :1555:63, :1560:40, :1562:69, :1576:42, :1579:76, :1582:40
        _GEN_1510 = will_fire_hella_incoming_0 & dmem_req_fire_0;	// lsu.scala:535:65, :752:55, :1540:50
        _GEN_1511 = _GEN_572 & _GEN_641 ? 3'h0 : hella_state;	// lsu.scala:242:38, :1288:54, :1562:35, :1582:40, :1584:69, :1585:21
        _GEN_1512 =
          {{_GEN_1511},
           {_GEN_1511},
           {will_fire_hella_wakeup_0 & dmem_req_fire_0 ? 3'h4 : hella_state},
           {_GEN_641 ? 3'h0 : _GEN_570 ? 3'h5 : hella_state},
           {3'h0},
           {{1'h1,
             |{hella_xcpt_ma_ld,
               hella_xcpt_ma_st,
               hella_xcpt_pf_ld,
               hella_xcpt_pf_st,
               hella_xcpt_ae_ld,
               hella_xcpt_ae_st},
             1'h0}},
           {io_hellacache_s1_kill ? (_GEN_1510 ? 3'h6 : 3'h0) : {2'h1, ~_GEN_1510}},
           {_GEN_1511}};	// lsu.scala:242:38, :246:34, :249:20, :535:65, :708:86, :752:55, :803:26, :820:26, :1287:7, :1288:28, :1312:58, :1533:38, :1539:34, :1540:{50,80}, :1541:21, :1543:21, :1545:85, :1546:19, :1548:19, :1550:{28,43}, :1552:17, :1553:{28,38}, :1555:{47,54,63}, :1556:19, :1558:19, :1560:40, :1562:{35,69}, :1563:21, :1572:76, :1573:21, :1576:42, :1579:{46,76}, :1580:19, :1582:40, :1584:69, :1585:21, util.scala:351:72
        hella_state <= _GEN_1512[hella_state];	// lsu.scala:242:38, :803:26, :820:26, :1288:28, :1533:38, :1539:34, :1550:{28,43}, :1552:17, :1553:{28,38}, :1555:63, :1560:40, :1562:69, :1576:42, :1579:76, :1582:40
      end
      else if (_GEN_1473)	// Decoupled.scala:40:37
        hella_state <= 3'h1;	// lsu.scala:242:38, :803:26
      live_store_mask <=
        ({16{dis_st_val_1}} & 16'h1 << _GEN_99 | _GEN_691)
        & ~{stq_15_valid & (|_GEN_620),
            stq_14_valid & (|_GEN_619),
            stq_13_valid & (|_GEN_618),
            stq_12_valid & (|_GEN_617),
            stq_11_valid & (|_GEN_616),
            stq_10_valid & (|_GEN_615),
            stq_9_valid & (|_GEN_614),
            stq_8_valid & (|_GEN_613),
            stq_7_valid & (|_GEN_612),
            stq_6_valid & (|_GEN_611),
            stq_5_valid & (|_GEN_610),
            stq_4_valid & (|_GEN_609),
            stq_3_valid & (|_GEN_608),
            stq_2_valid & (|_GEN_607),
            stq_1_valid & (|_GEN_606),
            stq_0_valid & (|_GEN_605)}
        & ~{_GEN_1476 & ~reset & _GEN_1508,
            _GEN_1476 & ~reset & _GEN_1506,
            _GEN_1476 & ~reset & _GEN_1504,
            _GEN_1476 & ~reset & _GEN_1502,
            _GEN_1476 & ~reset & _GEN_1500,
            _GEN_1476 & ~reset & _GEN_1498,
            _GEN_1476 & ~reset & _GEN_1496,
            _GEN_1476 & ~reset & _GEN_1494,
            _GEN_1476 & ~reset & _GEN_1492,
            _GEN_1476 & ~reset & _GEN_1490,
            _GEN_1476 & ~reset & _GEN_1488,
            _GEN_1476 & ~reset & _GEN_1486,
            _GEN_1476 & ~reset & _GEN_1484,
            _GEN_1476 & ~reset & _GEN_1482,
            _GEN_1476 & ~reset & _GEN_1480,
            _GEN_1476 & ~reset & _GEN_1478};	// lsu.scala:211:16, :259:32, :260:71, :302:85, :336:{31,72}, :338:21, :1401:25, :1404:5, :1408:7, :1596:22, :1597:3, :1602:5, :1622:38, :1623:9, :1647:{21,40,48}, :1648:{21,42}, util.scala:118:{51,59}
      if (fired_stad_incoming_REG)	// lsu.scala:895:51
        clr_bsy_valid_0 <=
          mem_stq_incoming_e_0_valid & ~mem_tlb_miss_0
          & ~mem_stq_incoming_e_0_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_incoming_e_0_bits_uop_br_mask) == 12'h0;	// lsu.scala:910:37, :925:41, :930:32, :942:29, :943:{29,68}, util.scala:118:{51,59}
      else if (fired_sta_incoming_REG)	// lsu.scala:896:51
        clr_bsy_valid_0 <=
          mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_data_valid
          & ~mem_tlb_miss_0 & ~mem_stq_incoming_e_0_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_incoming_e_0_bits_uop_br_mask) == 12'h0;	// lsu.scala:910:37, :925:41, :930:32, :950:29, :951:{29,69}, util.scala:118:{51,59}
      else if (fired_std_incoming_REG)	// lsu.scala:897:51
        clr_bsy_valid_0 <=
          mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_addr_valid
          & ~mem_stq_incoming_e_0_bits_addr_is_virtual
          & ~mem_stq_incoming_e_0_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_incoming_e_0_bits_uop_br_mask) == 12'h0;	// lsu.scala:910:37, :930:32, :958:29, :959:{29,74}, util.scala:118:{51,59}
      else	// lsu.scala:897:51
        clr_bsy_valid_0 <=
          fired_sfence_0 | fired_sta_retry_REG & mem_stq_retry_e_valid
          & mem_stq_retry_e_bits_data_valid & ~mem_tlb_miss_0
          & ~mem_stq_retry_e_bits_uop_is_amo
          & (io_core_brupdate_b1_mispredict_mask
             & mem_stq_retry_e_bits_uop_br_mask) == 12'h0;	// lsu.scala:899:37, :902:51, :913:37, :925:41, :930:32, :935:25, :963:35, :964:27, :967:38, :968:27, :970:29, :971:29, util.scala:118:{51,59}
      stdf_clr_bsy_valid <=
        fired_stdf_incoming & _GEN_2[mem_stdf_uop_stq_idx] & _GEN_87[mem_stdf_uop_stq_idx]
        & ~_GEN_90[mem_stdf_uop_stq_idx] & ~_GEN_61[mem_stdf_uop_stq_idx]
        & (io_core_brupdate_b1_mispredict_mask & mem_stdf_uop_br_mask) == 12'h0;	// lsu.scala:224:42, :898:37, :922:37, :983:37, :986:24, :989:30, :991:{26,62}, :993:29, :994:29, util.scala:118:{51,59}
      r_xcpt_valid <=
        (ld_xcpt_valid | mem_xcpt_valids_0) & ~io_core_exception
        & (io_core_brupdate_b1_mispredict_mask & xcpt_uop_br_mask) == 12'h0;	// lsu.scala:667:32, :669:22, :1235:29, :1238:44, :1243:21, :1245:34, :1246:39, util.scala:118:{51,59}
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:719];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [9:0] i = 10'h0; i < 10'h2D0; i += 10'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        ldq_0_valid = _RANDOM[10'h0][0];	// lsu.scala:210:16
        ldq_0_bits_uop_uopc = _RANDOM[10'h0][7:1];	// lsu.scala:210:16
        ldq_0_bits_uop_inst = {_RANDOM[10'h0][31:8], _RANDOM[10'h1][7:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_debug_inst = {_RANDOM[10'h1][31:8], _RANDOM[10'h2][7:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_is_rvc = _RANDOM[10'h2][8];	// lsu.scala:210:16
        ldq_0_bits_uop_debug_pc = {_RANDOM[10'h2][31:9], _RANDOM[10'h3][16:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_iq_type = _RANDOM[10'h3][19:17];	// lsu.scala:210:16
        ldq_0_bits_uop_fu_code = _RANDOM[10'h3][29:20];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_br_type = {_RANDOM[10'h3][31:30], _RANDOM[10'h4][1:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_op1_sel = _RANDOM[10'h4][3:2];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_op2_sel = _RANDOM[10'h4][6:4];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_imm_sel = _RANDOM[10'h4][9:7];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_op_fcn = _RANDOM[10'h4][13:10];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_fcn_dw = _RANDOM[10'h4][14];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_csr_cmd = _RANDOM[10'h4][17:15];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_is_load = _RANDOM[10'h4][18];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_is_sta = _RANDOM[10'h4][19];	// lsu.scala:210:16
        ldq_0_bits_uop_ctrl_is_std = _RANDOM[10'h4][20];	// lsu.scala:210:16
        ldq_0_bits_uop_iw_state = _RANDOM[10'h4][22:21];	// lsu.scala:210:16
        ldq_0_bits_uop_iw_p1_poisoned = _RANDOM[10'h4][23];	// lsu.scala:210:16
        ldq_0_bits_uop_iw_p2_poisoned = _RANDOM[10'h4][24];	// lsu.scala:210:16
        ldq_0_bits_uop_is_br = _RANDOM[10'h4][25];	// lsu.scala:210:16
        ldq_0_bits_uop_is_jalr = _RANDOM[10'h4][26];	// lsu.scala:210:16
        ldq_0_bits_uop_is_jal = _RANDOM[10'h4][27];	// lsu.scala:210:16
        ldq_0_bits_uop_is_sfb = _RANDOM[10'h4][28];	// lsu.scala:210:16
        ldq_0_bits_uop_br_mask = {_RANDOM[10'h4][31:29], _RANDOM[10'h5][8:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_br_tag = _RANDOM[10'h5][12:9];	// lsu.scala:210:16
        ldq_0_bits_uop_ftq_idx = _RANDOM[10'h5][17:13];	// lsu.scala:210:16
        ldq_0_bits_uop_edge_inst = _RANDOM[10'h5][18];	// lsu.scala:210:16
        ldq_0_bits_uop_pc_lob = _RANDOM[10'h5][24:19];	// lsu.scala:210:16
        ldq_0_bits_uop_taken = _RANDOM[10'h5][25];	// lsu.scala:210:16
        ldq_0_bits_uop_imm_packed = {_RANDOM[10'h5][31:26], _RANDOM[10'h6][13:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_csr_addr = _RANDOM[10'h6][25:14];	// lsu.scala:210:16
        ldq_0_bits_uop_rob_idx = _RANDOM[10'h6][31:26];	// lsu.scala:210:16
        ldq_0_bits_uop_ldq_idx = _RANDOM[10'h7][3:0];	// lsu.scala:210:16
        ldq_0_bits_uop_stq_idx = _RANDOM[10'h7][7:4];	// lsu.scala:210:16
        ldq_0_bits_uop_rxq_idx = _RANDOM[10'h7][9:8];	// lsu.scala:210:16
        ldq_0_bits_uop_pdst = _RANDOM[10'h7][16:10];	// lsu.scala:210:16
        ldq_0_bits_uop_prs1 = _RANDOM[10'h7][23:17];	// lsu.scala:210:16
        ldq_0_bits_uop_prs2 = _RANDOM[10'h7][30:24];	// lsu.scala:210:16
        ldq_0_bits_uop_prs3 = {_RANDOM[10'h7][31], _RANDOM[10'h8][5:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_ppred = _RANDOM[10'h8][10:6];	// lsu.scala:210:16
        ldq_0_bits_uop_prs1_busy = _RANDOM[10'h8][11];	// lsu.scala:210:16
        ldq_0_bits_uop_prs2_busy = _RANDOM[10'h8][12];	// lsu.scala:210:16
        ldq_0_bits_uop_prs3_busy = _RANDOM[10'h8][13];	// lsu.scala:210:16
        ldq_0_bits_uop_ppred_busy = _RANDOM[10'h8][14];	// lsu.scala:210:16
        ldq_0_bits_uop_stale_pdst = _RANDOM[10'h8][21:15];	// lsu.scala:210:16
        ldq_0_bits_uop_exception = _RANDOM[10'h8][22];	// lsu.scala:210:16
        ldq_0_bits_uop_exc_cause =
          {_RANDOM[10'h8][31:23], _RANDOM[10'h9], _RANDOM[10'hA][22:0]};	// lsu.scala:210:16
        ldq_0_bits_uop_bypassable = _RANDOM[10'hA][23];	// lsu.scala:210:16
        ldq_0_bits_uop_mem_cmd = _RANDOM[10'hA][28:24];	// lsu.scala:210:16
        ldq_0_bits_uop_mem_size = _RANDOM[10'hA][30:29];	// lsu.scala:210:16
        ldq_0_bits_uop_mem_signed = _RANDOM[10'hA][31];	// lsu.scala:210:16
        ldq_0_bits_uop_is_fence = _RANDOM[10'hB][0];	// lsu.scala:210:16
        ldq_0_bits_uop_is_fencei = _RANDOM[10'hB][1];	// lsu.scala:210:16
        ldq_0_bits_uop_is_amo = _RANDOM[10'hB][2];	// lsu.scala:210:16
        ldq_0_bits_uop_uses_ldq = _RANDOM[10'hB][3];	// lsu.scala:210:16
        ldq_0_bits_uop_uses_stq = _RANDOM[10'hB][4];	// lsu.scala:210:16
        ldq_0_bits_uop_is_sys_pc2epc = _RANDOM[10'hB][5];	// lsu.scala:210:16
        ldq_0_bits_uop_is_unique = _RANDOM[10'hB][6];	// lsu.scala:210:16
        ldq_0_bits_uop_flush_on_commit = _RANDOM[10'hB][7];	// lsu.scala:210:16
        ldq_0_bits_uop_ldst_is_rs1 = _RANDOM[10'hB][8];	// lsu.scala:210:16
        ldq_0_bits_uop_ldst = _RANDOM[10'hB][14:9];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs1 = _RANDOM[10'hB][20:15];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs2 = _RANDOM[10'hB][26:21];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs3 = {_RANDOM[10'hB][31:27], _RANDOM[10'hC][0]};	// lsu.scala:210:16
        ldq_0_bits_uop_ldst_val = _RANDOM[10'hC][1];	// lsu.scala:210:16
        ldq_0_bits_uop_dst_rtype = _RANDOM[10'hC][3:2];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs1_rtype = _RANDOM[10'hC][5:4];	// lsu.scala:210:16
        ldq_0_bits_uop_lrs2_rtype = _RANDOM[10'hC][7:6];	// lsu.scala:210:16
        ldq_0_bits_uop_frs3_en = _RANDOM[10'hC][8];	// lsu.scala:210:16
        ldq_0_bits_uop_fp_val = _RANDOM[10'hC][9];	// lsu.scala:210:16
        ldq_0_bits_uop_fp_single = _RANDOM[10'hC][10];	// lsu.scala:210:16
        ldq_0_bits_uop_xcpt_pf_if = _RANDOM[10'hC][11];	// lsu.scala:210:16
        ldq_0_bits_uop_xcpt_ae_if = _RANDOM[10'hC][12];	// lsu.scala:210:16
        ldq_0_bits_uop_xcpt_ma_if = _RANDOM[10'hC][13];	// lsu.scala:210:16
        ldq_0_bits_uop_bp_debug_if = _RANDOM[10'hC][14];	// lsu.scala:210:16
        ldq_0_bits_uop_bp_xcpt_if = _RANDOM[10'hC][15];	// lsu.scala:210:16
        ldq_0_bits_uop_debug_fsrc = _RANDOM[10'hC][17:16];	// lsu.scala:210:16
        ldq_0_bits_uop_debug_tsrc = _RANDOM[10'hC][19:18];	// lsu.scala:210:16
        ldq_0_bits_addr_valid = _RANDOM[10'hC][20];	// lsu.scala:210:16
        ldq_0_bits_addr_bits = {_RANDOM[10'hC][31:21], _RANDOM[10'hD][28:0]};	// lsu.scala:210:16
        ldq_0_bits_addr_is_virtual = _RANDOM[10'hD][29];	// lsu.scala:210:16
        ldq_0_bits_addr_is_uncacheable = _RANDOM[10'hD][30];	// lsu.scala:210:16
        ldq_0_bits_executed = _RANDOM[10'hD][31];	// lsu.scala:210:16
        ldq_0_bits_succeeded = _RANDOM[10'hE][0];	// lsu.scala:210:16
        ldq_0_bits_order_fail = _RANDOM[10'hE][1];	// lsu.scala:210:16
        ldq_0_bits_observed = _RANDOM[10'hE][2];	// lsu.scala:210:16
        ldq_0_bits_st_dep_mask = _RANDOM[10'hE][18:3];	// lsu.scala:210:16
        ldq_0_bits_youngest_stq_idx = _RANDOM[10'hE][22:19];	// lsu.scala:210:16
        ldq_0_bits_forward_std_val = _RANDOM[10'hE][23];	// lsu.scala:210:16
        ldq_0_bits_forward_stq_idx = _RANDOM[10'hE][27:24];	// lsu.scala:210:16
        ldq_1_valid = _RANDOM[10'h10][28];	// lsu.scala:210:16
        ldq_1_bits_uop_uopc = {_RANDOM[10'h10][31:29], _RANDOM[10'h11][3:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_inst = {_RANDOM[10'h11][31:4], _RANDOM[10'h12][3:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_debug_inst = {_RANDOM[10'h12][31:4], _RANDOM[10'h13][3:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_is_rvc = _RANDOM[10'h13][4];	// lsu.scala:210:16
        ldq_1_bits_uop_debug_pc = {_RANDOM[10'h13][31:5], _RANDOM[10'h14][12:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_iq_type = _RANDOM[10'h14][15:13];	// lsu.scala:210:16
        ldq_1_bits_uop_fu_code = _RANDOM[10'h14][25:16];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_br_type = _RANDOM[10'h14][29:26];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_op1_sel = _RANDOM[10'h14][31:30];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_op2_sel = _RANDOM[10'h15][2:0];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_imm_sel = _RANDOM[10'h15][5:3];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_op_fcn = _RANDOM[10'h15][9:6];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_fcn_dw = _RANDOM[10'h15][10];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_csr_cmd = _RANDOM[10'h15][13:11];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_is_load = _RANDOM[10'h15][14];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_is_sta = _RANDOM[10'h15][15];	// lsu.scala:210:16
        ldq_1_bits_uop_ctrl_is_std = _RANDOM[10'h15][16];	// lsu.scala:210:16
        ldq_1_bits_uop_iw_state = _RANDOM[10'h15][18:17];	// lsu.scala:210:16
        ldq_1_bits_uop_iw_p1_poisoned = _RANDOM[10'h15][19];	// lsu.scala:210:16
        ldq_1_bits_uop_iw_p2_poisoned = _RANDOM[10'h15][20];	// lsu.scala:210:16
        ldq_1_bits_uop_is_br = _RANDOM[10'h15][21];	// lsu.scala:210:16
        ldq_1_bits_uop_is_jalr = _RANDOM[10'h15][22];	// lsu.scala:210:16
        ldq_1_bits_uop_is_jal = _RANDOM[10'h15][23];	// lsu.scala:210:16
        ldq_1_bits_uop_is_sfb = _RANDOM[10'h15][24];	// lsu.scala:210:16
        ldq_1_bits_uop_br_mask = {_RANDOM[10'h15][31:25], _RANDOM[10'h16][4:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_br_tag = _RANDOM[10'h16][8:5];	// lsu.scala:210:16
        ldq_1_bits_uop_ftq_idx = _RANDOM[10'h16][13:9];	// lsu.scala:210:16
        ldq_1_bits_uop_edge_inst = _RANDOM[10'h16][14];	// lsu.scala:210:16
        ldq_1_bits_uop_pc_lob = _RANDOM[10'h16][20:15];	// lsu.scala:210:16
        ldq_1_bits_uop_taken = _RANDOM[10'h16][21];	// lsu.scala:210:16
        ldq_1_bits_uop_imm_packed = {_RANDOM[10'h16][31:22], _RANDOM[10'h17][9:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_csr_addr = _RANDOM[10'h17][21:10];	// lsu.scala:210:16
        ldq_1_bits_uop_rob_idx = _RANDOM[10'h17][27:22];	// lsu.scala:210:16
        ldq_1_bits_uop_ldq_idx = _RANDOM[10'h17][31:28];	// lsu.scala:210:16
        ldq_1_bits_uop_stq_idx = _RANDOM[10'h18][3:0];	// lsu.scala:210:16
        ldq_1_bits_uop_rxq_idx = _RANDOM[10'h18][5:4];	// lsu.scala:210:16
        ldq_1_bits_uop_pdst = _RANDOM[10'h18][12:6];	// lsu.scala:210:16
        ldq_1_bits_uop_prs1 = _RANDOM[10'h18][19:13];	// lsu.scala:210:16
        ldq_1_bits_uop_prs2 = _RANDOM[10'h18][26:20];	// lsu.scala:210:16
        ldq_1_bits_uop_prs3 = {_RANDOM[10'h18][31:27], _RANDOM[10'h19][1:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_ppred = _RANDOM[10'h19][6:2];	// lsu.scala:210:16
        ldq_1_bits_uop_prs1_busy = _RANDOM[10'h19][7];	// lsu.scala:210:16
        ldq_1_bits_uop_prs2_busy = _RANDOM[10'h19][8];	// lsu.scala:210:16
        ldq_1_bits_uop_prs3_busy = _RANDOM[10'h19][9];	// lsu.scala:210:16
        ldq_1_bits_uop_ppred_busy = _RANDOM[10'h19][10];	// lsu.scala:210:16
        ldq_1_bits_uop_stale_pdst = _RANDOM[10'h19][17:11];	// lsu.scala:210:16
        ldq_1_bits_uop_exception = _RANDOM[10'h19][18];	// lsu.scala:210:16
        ldq_1_bits_uop_exc_cause =
          {_RANDOM[10'h19][31:19], _RANDOM[10'h1A], _RANDOM[10'h1B][18:0]};	// lsu.scala:210:16
        ldq_1_bits_uop_bypassable = _RANDOM[10'h1B][19];	// lsu.scala:210:16
        ldq_1_bits_uop_mem_cmd = _RANDOM[10'h1B][24:20];	// lsu.scala:210:16
        ldq_1_bits_uop_mem_size = _RANDOM[10'h1B][26:25];	// lsu.scala:210:16
        ldq_1_bits_uop_mem_signed = _RANDOM[10'h1B][27];	// lsu.scala:210:16
        ldq_1_bits_uop_is_fence = _RANDOM[10'h1B][28];	// lsu.scala:210:16
        ldq_1_bits_uop_is_fencei = _RANDOM[10'h1B][29];	// lsu.scala:210:16
        ldq_1_bits_uop_is_amo = _RANDOM[10'h1B][30];	// lsu.scala:210:16
        ldq_1_bits_uop_uses_ldq = _RANDOM[10'h1B][31];	// lsu.scala:210:16
        ldq_1_bits_uop_uses_stq = _RANDOM[10'h1C][0];	// lsu.scala:210:16
        ldq_1_bits_uop_is_sys_pc2epc = _RANDOM[10'h1C][1];	// lsu.scala:210:16
        ldq_1_bits_uop_is_unique = _RANDOM[10'h1C][2];	// lsu.scala:210:16
        ldq_1_bits_uop_flush_on_commit = _RANDOM[10'h1C][3];	// lsu.scala:210:16
        ldq_1_bits_uop_ldst_is_rs1 = _RANDOM[10'h1C][4];	// lsu.scala:210:16
        ldq_1_bits_uop_ldst = _RANDOM[10'h1C][10:5];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs1 = _RANDOM[10'h1C][16:11];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs2 = _RANDOM[10'h1C][22:17];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs3 = _RANDOM[10'h1C][28:23];	// lsu.scala:210:16
        ldq_1_bits_uop_ldst_val = _RANDOM[10'h1C][29];	// lsu.scala:210:16
        ldq_1_bits_uop_dst_rtype = _RANDOM[10'h1C][31:30];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs1_rtype = _RANDOM[10'h1D][1:0];	// lsu.scala:210:16
        ldq_1_bits_uop_lrs2_rtype = _RANDOM[10'h1D][3:2];	// lsu.scala:210:16
        ldq_1_bits_uop_frs3_en = _RANDOM[10'h1D][4];	// lsu.scala:210:16
        ldq_1_bits_uop_fp_val = _RANDOM[10'h1D][5];	// lsu.scala:210:16
        ldq_1_bits_uop_fp_single = _RANDOM[10'h1D][6];	// lsu.scala:210:16
        ldq_1_bits_uop_xcpt_pf_if = _RANDOM[10'h1D][7];	// lsu.scala:210:16
        ldq_1_bits_uop_xcpt_ae_if = _RANDOM[10'h1D][8];	// lsu.scala:210:16
        ldq_1_bits_uop_xcpt_ma_if = _RANDOM[10'h1D][9];	// lsu.scala:210:16
        ldq_1_bits_uop_bp_debug_if = _RANDOM[10'h1D][10];	// lsu.scala:210:16
        ldq_1_bits_uop_bp_xcpt_if = _RANDOM[10'h1D][11];	// lsu.scala:210:16
        ldq_1_bits_uop_debug_fsrc = _RANDOM[10'h1D][13:12];	// lsu.scala:210:16
        ldq_1_bits_uop_debug_tsrc = _RANDOM[10'h1D][15:14];	// lsu.scala:210:16
        ldq_1_bits_addr_valid = _RANDOM[10'h1D][16];	// lsu.scala:210:16
        ldq_1_bits_addr_bits = {_RANDOM[10'h1D][31:17], _RANDOM[10'h1E][24:0]};	// lsu.scala:210:16
        ldq_1_bits_addr_is_virtual = _RANDOM[10'h1E][25];	// lsu.scala:210:16
        ldq_1_bits_addr_is_uncacheable = _RANDOM[10'h1E][26];	// lsu.scala:210:16
        ldq_1_bits_executed = _RANDOM[10'h1E][27];	// lsu.scala:210:16
        ldq_1_bits_succeeded = _RANDOM[10'h1E][28];	// lsu.scala:210:16
        ldq_1_bits_order_fail = _RANDOM[10'h1E][29];	// lsu.scala:210:16
        ldq_1_bits_observed = _RANDOM[10'h1E][30];	// lsu.scala:210:16
        ldq_1_bits_st_dep_mask = {_RANDOM[10'h1E][31], _RANDOM[10'h1F][14:0]};	// lsu.scala:210:16
        ldq_1_bits_youngest_stq_idx = _RANDOM[10'h1F][18:15];	// lsu.scala:210:16
        ldq_1_bits_forward_std_val = _RANDOM[10'h1F][19];	// lsu.scala:210:16
        ldq_1_bits_forward_stq_idx = _RANDOM[10'h1F][23:20];	// lsu.scala:210:16
        ldq_2_valid = _RANDOM[10'h21][24];	// lsu.scala:210:16
        ldq_2_bits_uop_uopc = _RANDOM[10'h21][31:25];	// lsu.scala:210:16
        ldq_2_bits_uop_inst = _RANDOM[10'h22];	// lsu.scala:210:16
        ldq_2_bits_uop_debug_inst = _RANDOM[10'h23];	// lsu.scala:210:16
        ldq_2_bits_uop_is_rvc = _RANDOM[10'h24][0];	// lsu.scala:210:16
        ldq_2_bits_uop_debug_pc = {_RANDOM[10'h24][31:1], _RANDOM[10'h25][8:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_iq_type = _RANDOM[10'h25][11:9];	// lsu.scala:210:16
        ldq_2_bits_uop_fu_code = _RANDOM[10'h25][21:12];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_br_type = _RANDOM[10'h25][25:22];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_op1_sel = _RANDOM[10'h25][27:26];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_op2_sel = _RANDOM[10'h25][30:28];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_imm_sel = {_RANDOM[10'h25][31], _RANDOM[10'h26][1:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_op_fcn = _RANDOM[10'h26][5:2];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_fcn_dw = _RANDOM[10'h26][6];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_csr_cmd = _RANDOM[10'h26][9:7];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_is_load = _RANDOM[10'h26][10];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_is_sta = _RANDOM[10'h26][11];	// lsu.scala:210:16
        ldq_2_bits_uop_ctrl_is_std = _RANDOM[10'h26][12];	// lsu.scala:210:16
        ldq_2_bits_uop_iw_state = _RANDOM[10'h26][14:13];	// lsu.scala:210:16
        ldq_2_bits_uop_iw_p1_poisoned = _RANDOM[10'h26][15];	// lsu.scala:210:16
        ldq_2_bits_uop_iw_p2_poisoned = _RANDOM[10'h26][16];	// lsu.scala:210:16
        ldq_2_bits_uop_is_br = _RANDOM[10'h26][17];	// lsu.scala:210:16
        ldq_2_bits_uop_is_jalr = _RANDOM[10'h26][18];	// lsu.scala:210:16
        ldq_2_bits_uop_is_jal = _RANDOM[10'h26][19];	// lsu.scala:210:16
        ldq_2_bits_uop_is_sfb = _RANDOM[10'h26][20];	// lsu.scala:210:16
        ldq_2_bits_uop_br_mask = {_RANDOM[10'h26][31:21], _RANDOM[10'h27][0]};	// lsu.scala:210:16
        ldq_2_bits_uop_br_tag = _RANDOM[10'h27][4:1];	// lsu.scala:210:16
        ldq_2_bits_uop_ftq_idx = _RANDOM[10'h27][9:5];	// lsu.scala:210:16
        ldq_2_bits_uop_edge_inst = _RANDOM[10'h27][10];	// lsu.scala:210:16
        ldq_2_bits_uop_pc_lob = _RANDOM[10'h27][16:11];	// lsu.scala:210:16
        ldq_2_bits_uop_taken = _RANDOM[10'h27][17];	// lsu.scala:210:16
        ldq_2_bits_uop_imm_packed = {_RANDOM[10'h27][31:18], _RANDOM[10'h28][5:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_csr_addr = _RANDOM[10'h28][17:6];	// lsu.scala:210:16
        ldq_2_bits_uop_rob_idx = _RANDOM[10'h28][23:18];	// lsu.scala:210:16
        ldq_2_bits_uop_ldq_idx = _RANDOM[10'h28][27:24];	// lsu.scala:210:16
        ldq_2_bits_uop_stq_idx = _RANDOM[10'h28][31:28];	// lsu.scala:210:16
        ldq_2_bits_uop_rxq_idx = _RANDOM[10'h29][1:0];	// lsu.scala:210:16
        ldq_2_bits_uop_pdst = _RANDOM[10'h29][8:2];	// lsu.scala:210:16
        ldq_2_bits_uop_prs1 = _RANDOM[10'h29][15:9];	// lsu.scala:210:16
        ldq_2_bits_uop_prs2 = _RANDOM[10'h29][22:16];	// lsu.scala:210:16
        ldq_2_bits_uop_prs3 = _RANDOM[10'h29][29:23];	// lsu.scala:210:16
        ldq_2_bits_uop_ppred = {_RANDOM[10'h29][31:30], _RANDOM[10'h2A][2:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_prs1_busy = _RANDOM[10'h2A][3];	// lsu.scala:210:16
        ldq_2_bits_uop_prs2_busy = _RANDOM[10'h2A][4];	// lsu.scala:210:16
        ldq_2_bits_uop_prs3_busy = _RANDOM[10'h2A][5];	// lsu.scala:210:16
        ldq_2_bits_uop_ppred_busy = _RANDOM[10'h2A][6];	// lsu.scala:210:16
        ldq_2_bits_uop_stale_pdst = _RANDOM[10'h2A][13:7];	// lsu.scala:210:16
        ldq_2_bits_uop_exception = _RANDOM[10'h2A][14];	// lsu.scala:210:16
        ldq_2_bits_uop_exc_cause =
          {_RANDOM[10'h2A][31:15], _RANDOM[10'h2B], _RANDOM[10'h2C][14:0]};	// lsu.scala:210:16
        ldq_2_bits_uop_bypassable = _RANDOM[10'h2C][15];	// lsu.scala:210:16
        ldq_2_bits_uop_mem_cmd = _RANDOM[10'h2C][20:16];	// lsu.scala:210:16
        ldq_2_bits_uop_mem_size = _RANDOM[10'h2C][22:21];	// lsu.scala:210:16
        ldq_2_bits_uop_mem_signed = _RANDOM[10'h2C][23];	// lsu.scala:210:16
        ldq_2_bits_uop_is_fence = _RANDOM[10'h2C][24];	// lsu.scala:210:16
        ldq_2_bits_uop_is_fencei = _RANDOM[10'h2C][25];	// lsu.scala:210:16
        ldq_2_bits_uop_is_amo = _RANDOM[10'h2C][26];	// lsu.scala:210:16
        ldq_2_bits_uop_uses_ldq = _RANDOM[10'h2C][27];	// lsu.scala:210:16
        ldq_2_bits_uop_uses_stq = _RANDOM[10'h2C][28];	// lsu.scala:210:16
        ldq_2_bits_uop_is_sys_pc2epc = _RANDOM[10'h2C][29];	// lsu.scala:210:16
        ldq_2_bits_uop_is_unique = _RANDOM[10'h2C][30];	// lsu.scala:210:16
        ldq_2_bits_uop_flush_on_commit = _RANDOM[10'h2C][31];	// lsu.scala:210:16
        ldq_2_bits_uop_ldst_is_rs1 = _RANDOM[10'h2D][0];	// lsu.scala:210:16
        ldq_2_bits_uop_ldst = _RANDOM[10'h2D][6:1];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs1 = _RANDOM[10'h2D][12:7];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs2 = _RANDOM[10'h2D][18:13];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs3 = _RANDOM[10'h2D][24:19];	// lsu.scala:210:16
        ldq_2_bits_uop_ldst_val = _RANDOM[10'h2D][25];	// lsu.scala:210:16
        ldq_2_bits_uop_dst_rtype = _RANDOM[10'h2D][27:26];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs1_rtype = _RANDOM[10'h2D][29:28];	// lsu.scala:210:16
        ldq_2_bits_uop_lrs2_rtype = _RANDOM[10'h2D][31:30];	// lsu.scala:210:16
        ldq_2_bits_uop_frs3_en = _RANDOM[10'h2E][0];	// lsu.scala:210:16
        ldq_2_bits_uop_fp_val = _RANDOM[10'h2E][1];	// lsu.scala:210:16
        ldq_2_bits_uop_fp_single = _RANDOM[10'h2E][2];	// lsu.scala:210:16
        ldq_2_bits_uop_xcpt_pf_if = _RANDOM[10'h2E][3];	// lsu.scala:210:16
        ldq_2_bits_uop_xcpt_ae_if = _RANDOM[10'h2E][4];	// lsu.scala:210:16
        ldq_2_bits_uop_xcpt_ma_if = _RANDOM[10'h2E][5];	// lsu.scala:210:16
        ldq_2_bits_uop_bp_debug_if = _RANDOM[10'h2E][6];	// lsu.scala:210:16
        ldq_2_bits_uop_bp_xcpt_if = _RANDOM[10'h2E][7];	// lsu.scala:210:16
        ldq_2_bits_uop_debug_fsrc = _RANDOM[10'h2E][9:8];	// lsu.scala:210:16
        ldq_2_bits_uop_debug_tsrc = _RANDOM[10'h2E][11:10];	// lsu.scala:210:16
        ldq_2_bits_addr_valid = _RANDOM[10'h2E][12];	// lsu.scala:210:16
        ldq_2_bits_addr_bits = {_RANDOM[10'h2E][31:13], _RANDOM[10'h2F][20:0]};	// lsu.scala:210:16
        ldq_2_bits_addr_is_virtual = _RANDOM[10'h2F][21];	// lsu.scala:210:16
        ldq_2_bits_addr_is_uncacheable = _RANDOM[10'h2F][22];	// lsu.scala:210:16
        ldq_2_bits_executed = _RANDOM[10'h2F][23];	// lsu.scala:210:16
        ldq_2_bits_succeeded = _RANDOM[10'h2F][24];	// lsu.scala:210:16
        ldq_2_bits_order_fail = _RANDOM[10'h2F][25];	// lsu.scala:210:16
        ldq_2_bits_observed = _RANDOM[10'h2F][26];	// lsu.scala:210:16
        ldq_2_bits_st_dep_mask = {_RANDOM[10'h2F][31:27], _RANDOM[10'h30][10:0]};	// lsu.scala:210:16
        ldq_2_bits_youngest_stq_idx = _RANDOM[10'h30][14:11];	// lsu.scala:210:16
        ldq_2_bits_forward_std_val = _RANDOM[10'h30][15];	// lsu.scala:210:16
        ldq_2_bits_forward_stq_idx = _RANDOM[10'h30][19:16];	// lsu.scala:210:16
        ldq_3_valid = _RANDOM[10'h32][20];	// lsu.scala:210:16
        ldq_3_bits_uop_uopc = _RANDOM[10'h32][27:21];	// lsu.scala:210:16
        ldq_3_bits_uop_inst = {_RANDOM[10'h32][31:28], _RANDOM[10'h33][27:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_debug_inst = {_RANDOM[10'h33][31:28], _RANDOM[10'h34][27:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_is_rvc = _RANDOM[10'h34][28];	// lsu.scala:210:16
        ldq_3_bits_uop_debug_pc =
          {_RANDOM[10'h34][31:29], _RANDOM[10'h35], _RANDOM[10'h36][4:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_iq_type = _RANDOM[10'h36][7:5];	// lsu.scala:210:16
        ldq_3_bits_uop_fu_code = _RANDOM[10'h36][17:8];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_br_type = _RANDOM[10'h36][21:18];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_op1_sel = _RANDOM[10'h36][23:22];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_op2_sel = _RANDOM[10'h36][26:24];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_imm_sel = _RANDOM[10'h36][29:27];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_op_fcn = {_RANDOM[10'h36][31:30], _RANDOM[10'h37][1:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_fcn_dw = _RANDOM[10'h37][2];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_csr_cmd = _RANDOM[10'h37][5:3];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_is_load = _RANDOM[10'h37][6];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_is_sta = _RANDOM[10'h37][7];	// lsu.scala:210:16
        ldq_3_bits_uop_ctrl_is_std = _RANDOM[10'h37][8];	// lsu.scala:210:16
        ldq_3_bits_uop_iw_state = _RANDOM[10'h37][10:9];	// lsu.scala:210:16
        ldq_3_bits_uop_iw_p1_poisoned = _RANDOM[10'h37][11];	// lsu.scala:210:16
        ldq_3_bits_uop_iw_p2_poisoned = _RANDOM[10'h37][12];	// lsu.scala:210:16
        ldq_3_bits_uop_is_br = _RANDOM[10'h37][13];	// lsu.scala:210:16
        ldq_3_bits_uop_is_jalr = _RANDOM[10'h37][14];	// lsu.scala:210:16
        ldq_3_bits_uop_is_jal = _RANDOM[10'h37][15];	// lsu.scala:210:16
        ldq_3_bits_uop_is_sfb = _RANDOM[10'h37][16];	// lsu.scala:210:16
        ldq_3_bits_uop_br_mask = _RANDOM[10'h37][28:17];	// lsu.scala:210:16
        ldq_3_bits_uop_br_tag = {_RANDOM[10'h37][31:29], _RANDOM[10'h38][0]};	// lsu.scala:210:16
        ldq_3_bits_uop_ftq_idx = _RANDOM[10'h38][5:1];	// lsu.scala:210:16
        ldq_3_bits_uop_edge_inst = _RANDOM[10'h38][6];	// lsu.scala:210:16
        ldq_3_bits_uop_pc_lob = _RANDOM[10'h38][12:7];	// lsu.scala:210:16
        ldq_3_bits_uop_taken = _RANDOM[10'h38][13];	// lsu.scala:210:16
        ldq_3_bits_uop_imm_packed = {_RANDOM[10'h38][31:14], _RANDOM[10'h39][1:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_csr_addr = _RANDOM[10'h39][13:2];	// lsu.scala:210:16
        ldq_3_bits_uop_rob_idx = _RANDOM[10'h39][19:14];	// lsu.scala:210:16
        ldq_3_bits_uop_ldq_idx = _RANDOM[10'h39][23:20];	// lsu.scala:210:16
        ldq_3_bits_uop_stq_idx = _RANDOM[10'h39][27:24];	// lsu.scala:210:16
        ldq_3_bits_uop_rxq_idx = _RANDOM[10'h39][29:28];	// lsu.scala:210:16
        ldq_3_bits_uop_pdst = {_RANDOM[10'h39][31:30], _RANDOM[10'h3A][4:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_prs1 = _RANDOM[10'h3A][11:5];	// lsu.scala:210:16
        ldq_3_bits_uop_prs2 = _RANDOM[10'h3A][18:12];	// lsu.scala:210:16
        ldq_3_bits_uop_prs3 = _RANDOM[10'h3A][25:19];	// lsu.scala:210:16
        ldq_3_bits_uop_ppred = _RANDOM[10'h3A][30:26];	// lsu.scala:210:16
        ldq_3_bits_uop_prs1_busy = _RANDOM[10'h3A][31];	// lsu.scala:210:16
        ldq_3_bits_uop_prs2_busy = _RANDOM[10'h3B][0];	// lsu.scala:210:16
        ldq_3_bits_uop_prs3_busy = _RANDOM[10'h3B][1];	// lsu.scala:210:16
        ldq_3_bits_uop_ppred_busy = _RANDOM[10'h3B][2];	// lsu.scala:210:16
        ldq_3_bits_uop_stale_pdst = _RANDOM[10'h3B][9:3];	// lsu.scala:210:16
        ldq_3_bits_uop_exception = _RANDOM[10'h3B][10];	// lsu.scala:210:16
        ldq_3_bits_uop_exc_cause =
          {_RANDOM[10'h3B][31:11], _RANDOM[10'h3C], _RANDOM[10'h3D][10:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_bypassable = _RANDOM[10'h3D][11];	// lsu.scala:210:16
        ldq_3_bits_uop_mem_cmd = _RANDOM[10'h3D][16:12];	// lsu.scala:210:16
        ldq_3_bits_uop_mem_size = _RANDOM[10'h3D][18:17];	// lsu.scala:210:16
        ldq_3_bits_uop_mem_signed = _RANDOM[10'h3D][19];	// lsu.scala:210:16
        ldq_3_bits_uop_is_fence = _RANDOM[10'h3D][20];	// lsu.scala:210:16
        ldq_3_bits_uop_is_fencei = _RANDOM[10'h3D][21];	// lsu.scala:210:16
        ldq_3_bits_uop_is_amo = _RANDOM[10'h3D][22];	// lsu.scala:210:16
        ldq_3_bits_uop_uses_ldq = _RANDOM[10'h3D][23];	// lsu.scala:210:16
        ldq_3_bits_uop_uses_stq = _RANDOM[10'h3D][24];	// lsu.scala:210:16
        ldq_3_bits_uop_is_sys_pc2epc = _RANDOM[10'h3D][25];	// lsu.scala:210:16
        ldq_3_bits_uop_is_unique = _RANDOM[10'h3D][26];	// lsu.scala:210:16
        ldq_3_bits_uop_flush_on_commit = _RANDOM[10'h3D][27];	// lsu.scala:210:16
        ldq_3_bits_uop_ldst_is_rs1 = _RANDOM[10'h3D][28];	// lsu.scala:210:16
        ldq_3_bits_uop_ldst = {_RANDOM[10'h3D][31:29], _RANDOM[10'h3E][2:0]};	// lsu.scala:210:16
        ldq_3_bits_uop_lrs1 = _RANDOM[10'h3E][8:3];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs2 = _RANDOM[10'h3E][14:9];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs3 = _RANDOM[10'h3E][20:15];	// lsu.scala:210:16
        ldq_3_bits_uop_ldst_val = _RANDOM[10'h3E][21];	// lsu.scala:210:16
        ldq_3_bits_uop_dst_rtype = _RANDOM[10'h3E][23:22];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs1_rtype = _RANDOM[10'h3E][25:24];	// lsu.scala:210:16
        ldq_3_bits_uop_lrs2_rtype = _RANDOM[10'h3E][27:26];	// lsu.scala:210:16
        ldq_3_bits_uop_frs3_en = _RANDOM[10'h3E][28];	// lsu.scala:210:16
        ldq_3_bits_uop_fp_val = _RANDOM[10'h3E][29];	// lsu.scala:210:16
        ldq_3_bits_uop_fp_single = _RANDOM[10'h3E][30];	// lsu.scala:210:16
        ldq_3_bits_uop_xcpt_pf_if = _RANDOM[10'h3E][31];	// lsu.scala:210:16
        ldq_3_bits_uop_xcpt_ae_if = _RANDOM[10'h3F][0];	// lsu.scala:210:16
        ldq_3_bits_uop_xcpt_ma_if = _RANDOM[10'h3F][1];	// lsu.scala:210:16
        ldq_3_bits_uop_bp_debug_if = _RANDOM[10'h3F][2];	// lsu.scala:210:16
        ldq_3_bits_uop_bp_xcpt_if = _RANDOM[10'h3F][3];	// lsu.scala:210:16
        ldq_3_bits_uop_debug_fsrc = _RANDOM[10'h3F][5:4];	// lsu.scala:210:16
        ldq_3_bits_uop_debug_tsrc = _RANDOM[10'h3F][7:6];	// lsu.scala:210:16
        ldq_3_bits_addr_valid = _RANDOM[10'h3F][8];	// lsu.scala:210:16
        ldq_3_bits_addr_bits = {_RANDOM[10'h3F][31:9], _RANDOM[10'h40][16:0]};	// lsu.scala:210:16
        ldq_3_bits_addr_is_virtual = _RANDOM[10'h40][17];	// lsu.scala:210:16
        ldq_3_bits_addr_is_uncacheable = _RANDOM[10'h40][18];	// lsu.scala:210:16
        ldq_3_bits_executed = _RANDOM[10'h40][19];	// lsu.scala:210:16
        ldq_3_bits_succeeded = _RANDOM[10'h40][20];	// lsu.scala:210:16
        ldq_3_bits_order_fail = _RANDOM[10'h40][21];	// lsu.scala:210:16
        ldq_3_bits_observed = _RANDOM[10'h40][22];	// lsu.scala:210:16
        ldq_3_bits_st_dep_mask = {_RANDOM[10'h40][31:23], _RANDOM[10'h41][6:0]};	// lsu.scala:210:16
        ldq_3_bits_youngest_stq_idx = _RANDOM[10'h41][10:7];	// lsu.scala:210:16
        ldq_3_bits_forward_std_val = _RANDOM[10'h41][11];	// lsu.scala:210:16
        ldq_3_bits_forward_stq_idx = _RANDOM[10'h41][15:12];	// lsu.scala:210:16
        ldq_4_valid = _RANDOM[10'h43][16];	// lsu.scala:210:16
        ldq_4_bits_uop_uopc = _RANDOM[10'h43][23:17];	// lsu.scala:210:16
        ldq_4_bits_uop_inst = {_RANDOM[10'h43][31:24], _RANDOM[10'h44][23:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_debug_inst = {_RANDOM[10'h44][31:24], _RANDOM[10'h45][23:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_is_rvc = _RANDOM[10'h45][24];	// lsu.scala:210:16
        ldq_4_bits_uop_debug_pc =
          {_RANDOM[10'h45][31:25], _RANDOM[10'h46], _RANDOM[10'h47][0]};	// lsu.scala:210:16
        ldq_4_bits_uop_iq_type = _RANDOM[10'h47][3:1];	// lsu.scala:210:16
        ldq_4_bits_uop_fu_code = _RANDOM[10'h47][13:4];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_br_type = _RANDOM[10'h47][17:14];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_op1_sel = _RANDOM[10'h47][19:18];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_op2_sel = _RANDOM[10'h47][22:20];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_imm_sel = _RANDOM[10'h47][25:23];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_op_fcn = _RANDOM[10'h47][29:26];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_fcn_dw = _RANDOM[10'h47][30];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h47][31], _RANDOM[10'h48][1:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_is_load = _RANDOM[10'h48][2];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_is_sta = _RANDOM[10'h48][3];	// lsu.scala:210:16
        ldq_4_bits_uop_ctrl_is_std = _RANDOM[10'h48][4];	// lsu.scala:210:16
        ldq_4_bits_uop_iw_state = _RANDOM[10'h48][6:5];	// lsu.scala:210:16
        ldq_4_bits_uop_iw_p1_poisoned = _RANDOM[10'h48][7];	// lsu.scala:210:16
        ldq_4_bits_uop_iw_p2_poisoned = _RANDOM[10'h48][8];	// lsu.scala:210:16
        ldq_4_bits_uop_is_br = _RANDOM[10'h48][9];	// lsu.scala:210:16
        ldq_4_bits_uop_is_jalr = _RANDOM[10'h48][10];	// lsu.scala:210:16
        ldq_4_bits_uop_is_jal = _RANDOM[10'h48][11];	// lsu.scala:210:16
        ldq_4_bits_uop_is_sfb = _RANDOM[10'h48][12];	// lsu.scala:210:16
        ldq_4_bits_uop_br_mask = _RANDOM[10'h48][24:13];	// lsu.scala:210:16
        ldq_4_bits_uop_br_tag = _RANDOM[10'h48][28:25];	// lsu.scala:210:16
        ldq_4_bits_uop_ftq_idx = {_RANDOM[10'h48][31:29], _RANDOM[10'h49][1:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_edge_inst = _RANDOM[10'h49][2];	// lsu.scala:210:16
        ldq_4_bits_uop_pc_lob = _RANDOM[10'h49][8:3];	// lsu.scala:210:16
        ldq_4_bits_uop_taken = _RANDOM[10'h49][9];	// lsu.scala:210:16
        ldq_4_bits_uop_imm_packed = _RANDOM[10'h49][29:10];	// lsu.scala:210:16
        ldq_4_bits_uop_csr_addr = {_RANDOM[10'h49][31:30], _RANDOM[10'h4A][9:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_rob_idx = _RANDOM[10'h4A][15:10];	// lsu.scala:210:16
        ldq_4_bits_uop_ldq_idx = _RANDOM[10'h4A][19:16];	// lsu.scala:210:16
        ldq_4_bits_uop_stq_idx = _RANDOM[10'h4A][23:20];	// lsu.scala:210:16
        ldq_4_bits_uop_rxq_idx = _RANDOM[10'h4A][25:24];	// lsu.scala:210:16
        ldq_4_bits_uop_pdst = {_RANDOM[10'h4A][31:26], _RANDOM[10'h4B][0]};	// lsu.scala:210:16
        ldq_4_bits_uop_prs1 = _RANDOM[10'h4B][7:1];	// lsu.scala:210:16
        ldq_4_bits_uop_prs2 = _RANDOM[10'h4B][14:8];	// lsu.scala:210:16
        ldq_4_bits_uop_prs3 = _RANDOM[10'h4B][21:15];	// lsu.scala:210:16
        ldq_4_bits_uop_ppred = _RANDOM[10'h4B][26:22];	// lsu.scala:210:16
        ldq_4_bits_uop_prs1_busy = _RANDOM[10'h4B][27];	// lsu.scala:210:16
        ldq_4_bits_uop_prs2_busy = _RANDOM[10'h4B][28];	// lsu.scala:210:16
        ldq_4_bits_uop_prs3_busy = _RANDOM[10'h4B][29];	// lsu.scala:210:16
        ldq_4_bits_uop_ppred_busy = _RANDOM[10'h4B][30];	// lsu.scala:210:16
        ldq_4_bits_uop_stale_pdst = {_RANDOM[10'h4B][31], _RANDOM[10'h4C][5:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_exception = _RANDOM[10'h4C][6];	// lsu.scala:210:16
        ldq_4_bits_uop_exc_cause =
          {_RANDOM[10'h4C][31:7], _RANDOM[10'h4D], _RANDOM[10'h4E][6:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_bypassable = _RANDOM[10'h4E][7];	// lsu.scala:210:16
        ldq_4_bits_uop_mem_cmd = _RANDOM[10'h4E][12:8];	// lsu.scala:210:16
        ldq_4_bits_uop_mem_size = _RANDOM[10'h4E][14:13];	// lsu.scala:210:16
        ldq_4_bits_uop_mem_signed = _RANDOM[10'h4E][15];	// lsu.scala:210:16
        ldq_4_bits_uop_is_fence = _RANDOM[10'h4E][16];	// lsu.scala:210:16
        ldq_4_bits_uop_is_fencei = _RANDOM[10'h4E][17];	// lsu.scala:210:16
        ldq_4_bits_uop_is_amo = _RANDOM[10'h4E][18];	// lsu.scala:210:16
        ldq_4_bits_uop_uses_ldq = _RANDOM[10'h4E][19];	// lsu.scala:210:16
        ldq_4_bits_uop_uses_stq = _RANDOM[10'h4E][20];	// lsu.scala:210:16
        ldq_4_bits_uop_is_sys_pc2epc = _RANDOM[10'h4E][21];	// lsu.scala:210:16
        ldq_4_bits_uop_is_unique = _RANDOM[10'h4E][22];	// lsu.scala:210:16
        ldq_4_bits_uop_flush_on_commit = _RANDOM[10'h4E][23];	// lsu.scala:210:16
        ldq_4_bits_uop_ldst_is_rs1 = _RANDOM[10'h4E][24];	// lsu.scala:210:16
        ldq_4_bits_uop_ldst = _RANDOM[10'h4E][30:25];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs1 = {_RANDOM[10'h4E][31], _RANDOM[10'h4F][4:0]};	// lsu.scala:210:16
        ldq_4_bits_uop_lrs2 = _RANDOM[10'h4F][10:5];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs3 = _RANDOM[10'h4F][16:11];	// lsu.scala:210:16
        ldq_4_bits_uop_ldst_val = _RANDOM[10'h4F][17];	// lsu.scala:210:16
        ldq_4_bits_uop_dst_rtype = _RANDOM[10'h4F][19:18];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs1_rtype = _RANDOM[10'h4F][21:20];	// lsu.scala:210:16
        ldq_4_bits_uop_lrs2_rtype = _RANDOM[10'h4F][23:22];	// lsu.scala:210:16
        ldq_4_bits_uop_frs3_en = _RANDOM[10'h4F][24];	// lsu.scala:210:16
        ldq_4_bits_uop_fp_val = _RANDOM[10'h4F][25];	// lsu.scala:210:16
        ldq_4_bits_uop_fp_single = _RANDOM[10'h4F][26];	// lsu.scala:210:16
        ldq_4_bits_uop_xcpt_pf_if = _RANDOM[10'h4F][27];	// lsu.scala:210:16
        ldq_4_bits_uop_xcpt_ae_if = _RANDOM[10'h4F][28];	// lsu.scala:210:16
        ldq_4_bits_uop_xcpt_ma_if = _RANDOM[10'h4F][29];	// lsu.scala:210:16
        ldq_4_bits_uop_bp_debug_if = _RANDOM[10'h4F][30];	// lsu.scala:210:16
        ldq_4_bits_uop_bp_xcpt_if = _RANDOM[10'h4F][31];	// lsu.scala:210:16
        ldq_4_bits_uop_debug_fsrc = _RANDOM[10'h50][1:0];	// lsu.scala:210:16
        ldq_4_bits_uop_debug_tsrc = _RANDOM[10'h50][3:2];	// lsu.scala:210:16
        ldq_4_bits_addr_valid = _RANDOM[10'h50][4];	// lsu.scala:210:16
        ldq_4_bits_addr_bits = {_RANDOM[10'h50][31:5], _RANDOM[10'h51][12:0]};	// lsu.scala:210:16
        ldq_4_bits_addr_is_virtual = _RANDOM[10'h51][13];	// lsu.scala:210:16
        ldq_4_bits_addr_is_uncacheable = _RANDOM[10'h51][14];	// lsu.scala:210:16
        ldq_4_bits_executed = _RANDOM[10'h51][15];	// lsu.scala:210:16
        ldq_4_bits_succeeded = _RANDOM[10'h51][16];	// lsu.scala:210:16
        ldq_4_bits_order_fail = _RANDOM[10'h51][17];	// lsu.scala:210:16
        ldq_4_bits_observed = _RANDOM[10'h51][18];	// lsu.scala:210:16
        ldq_4_bits_st_dep_mask = {_RANDOM[10'h51][31:19], _RANDOM[10'h52][2:0]};	// lsu.scala:210:16
        ldq_4_bits_youngest_stq_idx = _RANDOM[10'h52][6:3];	// lsu.scala:210:16
        ldq_4_bits_forward_std_val = _RANDOM[10'h52][7];	// lsu.scala:210:16
        ldq_4_bits_forward_stq_idx = _RANDOM[10'h52][11:8];	// lsu.scala:210:16
        ldq_5_valid = _RANDOM[10'h54][12];	// lsu.scala:210:16
        ldq_5_bits_uop_uopc = _RANDOM[10'h54][19:13];	// lsu.scala:210:16
        ldq_5_bits_uop_inst = {_RANDOM[10'h54][31:20], _RANDOM[10'h55][19:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_debug_inst = {_RANDOM[10'h55][31:20], _RANDOM[10'h56][19:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_is_rvc = _RANDOM[10'h56][20];	// lsu.scala:210:16
        ldq_5_bits_uop_debug_pc = {_RANDOM[10'h56][31:21], _RANDOM[10'h57][28:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_iq_type = _RANDOM[10'h57][31:29];	// lsu.scala:210:16
        ldq_5_bits_uop_fu_code = _RANDOM[10'h58][9:0];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_br_type = _RANDOM[10'h58][13:10];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_op1_sel = _RANDOM[10'h58][15:14];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_op2_sel = _RANDOM[10'h58][18:16];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_imm_sel = _RANDOM[10'h58][21:19];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_op_fcn = _RANDOM[10'h58][25:22];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_fcn_dw = _RANDOM[10'h58][26];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_csr_cmd = _RANDOM[10'h58][29:27];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_is_load = _RANDOM[10'h58][30];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_is_sta = _RANDOM[10'h58][31];	// lsu.scala:210:16
        ldq_5_bits_uop_ctrl_is_std = _RANDOM[10'h59][0];	// lsu.scala:210:16
        ldq_5_bits_uop_iw_state = _RANDOM[10'h59][2:1];	// lsu.scala:210:16
        ldq_5_bits_uop_iw_p1_poisoned = _RANDOM[10'h59][3];	// lsu.scala:210:16
        ldq_5_bits_uop_iw_p2_poisoned = _RANDOM[10'h59][4];	// lsu.scala:210:16
        ldq_5_bits_uop_is_br = _RANDOM[10'h59][5];	// lsu.scala:210:16
        ldq_5_bits_uop_is_jalr = _RANDOM[10'h59][6];	// lsu.scala:210:16
        ldq_5_bits_uop_is_jal = _RANDOM[10'h59][7];	// lsu.scala:210:16
        ldq_5_bits_uop_is_sfb = _RANDOM[10'h59][8];	// lsu.scala:210:16
        ldq_5_bits_uop_br_mask = _RANDOM[10'h59][20:9];	// lsu.scala:210:16
        ldq_5_bits_uop_br_tag = _RANDOM[10'h59][24:21];	// lsu.scala:210:16
        ldq_5_bits_uop_ftq_idx = _RANDOM[10'h59][29:25];	// lsu.scala:210:16
        ldq_5_bits_uop_edge_inst = _RANDOM[10'h59][30];	// lsu.scala:210:16
        ldq_5_bits_uop_pc_lob = {_RANDOM[10'h59][31], _RANDOM[10'h5A][4:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_taken = _RANDOM[10'h5A][5];	// lsu.scala:210:16
        ldq_5_bits_uop_imm_packed = _RANDOM[10'h5A][25:6];	// lsu.scala:210:16
        ldq_5_bits_uop_csr_addr = {_RANDOM[10'h5A][31:26], _RANDOM[10'h5B][5:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_rob_idx = _RANDOM[10'h5B][11:6];	// lsu.scala:210:16
        ldq_5_bits_uop_ldq_idx = _RANDOM[10'h5B][15:12];	// lsu.scala:210:16
        ldq_5_bits_uop_stq_idx = _RANDOM[10'h5B][19:16];	// lsu.scala:210:16
        ldq_5_bits_uop_rxq_idx = _RANDOM[10'h5B][21:20];	// lsu.scala:210:16
        ldq_5_bits_uop_pdst = _RANDOM[10'h5B][28:22];	// lsu.scala:210:16
        ldq_5_bits_uop_prs1 = {_RANDOM[10'h5B][31:29], _RANDOM[10'h5C][3:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_prs2 = _RANDOM[10'h5C][10:4];	// lsu.scala:210:16
        ldq_5_bits_uop_prs3 = _RANDOM[10'h5C][17:11];	// lsu.scala:210:16
        ldq_5_bits_uop_ppred = _RANDOM[10'h5C][22:18];	// lsu.scala:210:16
        ldq_5_bits_uop_prs1_busy = _RANDOM[10'h5C][23];	// lsu.scala:210:16
        ldq_5_bits_uop_prs2_busy = _RANDOM[10'h5C][24];	// lsu.scala:210:16
        ldq_5_bits_uop_prs3_busy = _RANDOM[10'h5C][25];	// lsu.scala:210:16
        ldq_5_bits_uop_ppred_busy = _RANDOM[10'h5C][26];	// lsu.scala:210:16
        ldq_5_bits_uop_stale_pdst = {_RANDOM[10'h5C][31:27], _RANDOM[10'h5D][1:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_exception = _RANDOM[10'h5D][2];	// lsu.scala:210:16
        ldq_5_bits_uop_exc_cause =
          {_RANDOM[10'h5D][31:3], _RANDOM[10'h5E], _RANDOM[10'h5F][2:0]};	// lsu.scala:210:16
        ldq_5_bits_uop_bypassable = _RANDOM[10'h5F][3];	// lsu.scala:210:16
        ldq_5_bits_uop_mem_cmd = _RANDOM[10'h5F][8:4];	// lsu.scala:210:16
        ldq_5_bits_uop_mem_size = _RANDOM[10'h5F][10:9];	// lsu.scala:210:16
        ldq_5_bits_uop_mem_signed = _RANDOM[10'h5F][11];	// lsu.scala:210:16
        ldq_5_bits_uop_is_fence = _RANDOM[10'h5F][12];	// lsu.scala:210:16
        ldq_5_bits_uop_is_fencei = _RANDOM[10'h5F][13];	// lsu.scala:210:16
        ldq_5_bits_uop_is_amo = _RANDOM[10'h5F][14];	// lsu.scala:210:16
        ldq_5_bits_uop_uses_ldq = _RANDOM[10'h5F][15];	// lsu.scala:210:16
        ldq_5_bits_uop_uses_stq = _RANDOM[10'h5F][16];	// lsu.scala:210:16
        ldq_5_bits_uop_is_sys_pc2epc = _RANDOM[10'h5F][17];	// lsu.scala:210:16
        ldq_5_bits_uop_is_unique = _RANDOM[10'h5F][18];	// lsu.scala:210:16
        ldq_5_bits_uop_flush_on_commit = _RANDOM[10'h5F][19];	// lsu.scala:210:16
        ldq_5_bits_uop_ldst_is_rs1 = _RANDOM[10'h5F][20];	// lsu.scala:210:16
        ldq_5_bits_uop_ldst = _RANDOM[10'h5F][26:21];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs1 = {_RANDOM[10'h5F][31:27], _RANDOM[10'h60][0]};	// lsu.scala:210:16
        ldq_5_bits_uop_lrs2 = _RANDOM[10'h60][6:1];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs3 = _RANDOM[10'h60][12:7];	// lsu.scala:210:16
        ldq_5_bits_uop_ldst_val = _RANDOM[10'h60][13];	// lsu.scala:210:16
        ldq_5_bits_uop_dst_rtype = _RANDOM[10'h60][15:14];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs1_rtype = _RANDOM[10'h60][17:16];	// lsu.scala:210:16
        ldq_5_bits_uop_lrs2_rtype = _RANDOM[10'h60][19:18];	// lsu.scala:210:16
        ldq_5_bits_uop_frs3_en = _RANDOM[10'h60][20];	// lsu.scala:210:16
        ldq_5_bits_uop_fp_val = _RANDOM[10'h60][21];	// lsu.scala:210:16
        ldq_5_bits_uop_fp_single = _RANDOM[10'h60][22];	// lsu.scala:210:16
        ldq_5_bits_uop_xcpt_pf_if = _RANDOM[10'h60][23];	// lsu.scala:210:16
        ldq_5_bits_uop_xcpt_ae_if = _RANDOM[10'h60][24];	// lsu.scala:210:16
        ldq_5_bits_uop_xcpt_ma_if = _RANDOM[10'h60][25];	// lsu.scala:210:16
        ldq_5_bits_uop_bp_debug_if = _RANDOM[10'h60][26];	// lsu.scala:210:16
        ldq_5_bits_uop_bp_xcpt_if = _RANDOM[10'h60][27];	// lsu.scala:210:16
        ldq_5_bits_uop_debug_fsrc = _RANDOM[10'h60][29:28];	// lsu.scala:210:16
        ldq_5_bits_uop_debug_tsrc = _RANDOM[10'h60][31:30];	// lsu.scala:210:16
        ldq_5_bits_addr_valid = _RANDOM[10'h61][0];	// lsu.scala:210:16
        ldq_5_bits_addr_bits = {_RANDOM[10'h61][31:1], _RANDOM[10'h62][8:0]};	// lsu.scala:210:16
        ldq_5_bits_addr_is_virtual = _RANDOM[10'h62][9];	// lsu.scala:210:16
        ldq_5_bits_addr_is_uncacheable = _RANDOM[10'h62][10];	// lsu.scala:210:16
        ldq_5_bits_executed = _RANDOM[10'h62][11];	// lsu.scala:210:16
        ldq_5_bits_succeeded = _RANDOM[10'h62][12];	// lsu.scala:210:16
        ldq_5_bits_order_fail = _RANDOM[10'h62][13];	// lsu.scala:210:16
        ldq_5_bits_observed = _RANDOM[10'h62][14];	// lsu.scala:210:16
        ldq_5_bits_st_dep_mask = _RANDOM[10'h62][30:15];	// lsu.scala:210:16
        ldq_5_bits_youngest_stq_idx = {_RANDOM[10'h62][31], _RANDOM[10'h63][2:0]};	// lsu.scala:210:16
        ldq_5_bits_forward_std_val = _RANDOM[10'h63][3];	// lsu.scala:210:16
        ldq_5_bits_forward_stq_idx = _RANDOM[10'h63][7:4];	// lsu.scala:210:16
        ldq_6_valid = _RANDOM[10'h65][8];	// lsu.scala:210:16
        ldq_6_bits_uop_uopc = _RANDOM[10'h65][15:9];	// lsu.scala:210:16
        ldq_6_bits_uop_inst = {_RANDOM[10'h65][31:16], _RANDOM[10'h66][15:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_debug_inst = {_RANDOM[10'h66][31:16], _RANDOM[10'h67][15:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_is_rvc = _RANDOM[10'h67][16];	// lsu.scala:210:16
        ldq_6_bits_uop_debug_pc = {_RANDOM[10'h67][31:17], _RANDOM[10'h68][24:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_iq_type = _RANDOM[10'h68][27:25];	// lsu.scala:210:16
        ldq_6_bits_uop_fu_code = {_RANDOM[10'h68][31:28], _RANDOM[10'h69][5:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_br_type = _RANDOM[10'h69][9:6];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_op1_sel = _RANDOM[10'h69][11:10];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_op2_sel = _RANDOM[10'h69][14:12];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_imm_sel = _RANDOM[10'h69][17:15];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_op_fcn = _RANDOM[10'h69][21:18];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_fcn_dw = _RANDOM[10'h69][22];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_csr_cmd = _RANDOM[10'h69][25:23];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_is_load = _RANDOM[10'h69][26];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_is_sta = _RANDOM[10'h69][27];	// lsu.scala:210:16
        ldq_6_bits_uop_ctrl_is_std = _RANDOM[10'h69][28];	// lsu.scala:210:16
        ldq_6_bits_uop_iw_state = _RANDOM[10'h69][30:29];	// lsu.scala:210:16
        ldq_6_bits_uop_iw_p1_poisoned = _RANDOM[10'h69][31];	// lsu.scala:210:16
        ldq_6_bits_uop_iw_p2_poisoned = _RANDOM[10'h6A][0];	// lsu.scala:210:16
        ldq_6_bits_uop_is_br = _RANDOM[10'h6A][1];	// lsu.scala:210:16
        ldq_6_bits_uop_is_jalr = _RANDOM[10'h6A][2];	// lsu.scala:210:16
        ldq_6_bits_uop_is_jal = _RANDOM[10'h6A][3];	// lsu.scala:210:16
        ldq_6_bits_uop_is_sfb = _RANDOM[10'h6A][4];	// lsu.scala:210:16
        ldq_6_bits_uop_br_mask = _RANDOM[10'h6A][16:5];	// lsu.scala:210:16
        ldq_6_bits_uop_br_tag = _RANDOM[10'h6A][20:17];	// lsu.scala:210:16
        ldq_6_bits_uop_ftq_idx = _RANDOM[10'h6A][25:21];	// lsu.scala:210:16
        ldq_6_bits_uop_edge_inst = _RANDOM[10'h6A][26];	// lsu.scala:210:16
        ldq_6_bits_uop_pc_lob = {_RANDOM[10'h6A][31:27], _RANDOM[10'h6B][0]};	// lsu.scala:210:16
        ldq_6_bits_uop_taken = _RANDOM[10'h6B][1];	// lsu.scala:210:16
        ldq_6_bits_uop_imm_packed = _RANDOM[10'h6B][21:2];	// lsu.scala:210:16
        ldq_6_bits_uop_csr_addr = {_RANDOM[10'h6B][31:22], _RANDOM[10'h6C][1:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_rob_idx = _RANDOM[10'h6C][7:2];	// lsu.scala:210:16
        ldq_6_bits_uop_ldq_idx = _RANDOM[10'h6C][11:8];	// lsu.scala:210:16
        ldq_6_bits_uop_stq_idx = _RANDOM[10'h6C][15:12];	// lsu.scala:210:16
        ldq_6_bits_uop_rxq_idx = _RANDOM[10'h6C][17:16];	// lsu.scala:210:16
        ldq_6_bits_uop_pdst = _RANDOM[10'h6C][24:18];	// lsu.scala:210:16
        ldq_6_bits_uop_prs1 = _RANDOM[10'h6C][31:25];	// lsu.scala:210:16
        ldq_6_bits_uop_prs2 = _RANDOM[10'h6D][6:0];	// lsu.scala:210:16
        ldq_6_bits_uop_prs3 = _RANDOM[10'h6D][13:7];	// lsu.scala:210:16
        ldq_6_bits_uop_ppred = _RANDOM[10'h6D][18:14];	// lsu.scala:210:16
        ldq_6_bits_uop_prs1_busy = _RANDOM[10'h6D][19];	// lsu.scala:210:16
        ldq_6_bits_uop_prs2_busy = _RANDOM[10'h6D][20];	// lsu.scala:210:16
        ldq_6_bits_uop_prs3_busy = _RANDOM[10'h6D][21];	// lsu.scala:210:16
        ldq_6_bits_uop_ppred_busy = _RANDOM[10'h6D][22];	// lsu.scala:210:16
        ldq_6_bits_uop_stale_pdst = _RANDOM[10'h6D][29:23];	// lsu.scala:210:16
        ldq_6_bits_uop_exception = _RANDOM[10'h6D][30];	// lsu.scala:210:16
        ldq_6_bits_uop_exc_cause =
          {_RANDOM[10'h6D][31], _RANDOM[10'h6E], _RANDOM[10'h6F][30:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_bypassable = _RANDOM[10'h6F][31];	// lsu.scala:210:16
        ldq_6_bits_uop_mem_cmd = _RANDOM[10'h70][4:0];	// lsu.scala:210:16
        ldq_6_bits_uop_mem_size = _RANDOM[10'h70][6:5];	// lsu.scala:210:16
        ldq_6_bits_uop_mem_signed = _RANDOM[10'h70][7];	// lsu.scala:210:16
        ldq_6_bits_uop_is_fence = _RANDOM[10'h70][8];	// lsu.scala:210:16
        ldq_6_bits_uop_is_fencei = _RANDOM[10'h70][9];	// lsu.scala:210:16
        ldq_6_bits_uop_is_amo = _RANDOM[10'h70][10];	// lsu.scala:210:16
        ldq_6_bits_uop_uses_ldq = _RANDOM[10'h70][11];	// lsu.scala:210:16
        ldq_6_bits_uop_uses_stq = _RANDOM[10'h70][12];	// lsu.scala:210:16
        ldq_6_bits_uop_is_sys_pc2epc = _RANDOM[10'h70][13];	// lsu.scala:210:16
        ldq_6_bits_uop_is_unique = _RANDOM[10'h70][14];	// lsu.scala:210:16
        ldq_6_bits_uop_flush_on_commit = _RANDOM[10'h70][15];	// lsu.scala:210:16
        ldq_6_bits_uop_ldst_is_rs1 = _RANDOM[10'h70][16];	// lsu.scala:210:16
        ldq_6_bits_uop_ldst = _RANDOM[10'h70][22:17];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs1 = _RANDOM[10'h70][28:23];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs2 = {_RANDOM[10'h70][31:29], _RANDOM[10'h71][2:0]};	// lsu.scala:210:16
        ldq_6_bits_uop_lrs3 = _RANDOM[10'h71][8:3];	// lsu.scala:210:16
        ldq_6_bits_uop_ldst_val = _RANDOM[10'h71][9];	// lsu.scala:210:16
        ldq_6_bits_uop_dst_rtype = _RANDOM[10'h71][11:10];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs1_rtype = _RANDOM[10'h71][13:12];	// lsu.scala:210:16
        ldq_6_bits_uop_lrs2_rtype = _RANDOM[10'h71][15:14];	// lsu.scala:210:16
        ldq_6_bits_uop_frs3_en = _RANDOM[10'h71][16];	// lsu.scala:210:16
        ldq_6_bits_uop_fp_val = _RANDOM[10'h71][17];	// lsu.scala:210:16
        ldq_6_bits_uop_fp_single = _RANDOM[10'h71][18];	// lsu.scala:210:16
        ldq_6_bits_uop_xcpt_pf_if = _RANDOM[10'h71][19];	// lsu.scala:210:16
        ldq_6_bits_uop_xcpt_ae_if = _RANDOM[10'h71][20];	// lsu.scala:210:16
        ldq_6_bits_uop_xcpt_ma_if = _RANDOM[10'h71][21];	// lsu.scala:210:16
        ldq_6_bits_uop_bp_debug_if = _RANDOM[10'h71][22];	// lsu.scala:210:16
        ldq_6_bits_uop_bp_xcpt_if = _RANDOM[10'h71][23];	// lsu.scala:210:16
        ldq_6_bits_uop_debug_fsrc = _RANDOM[10'h71][25:24];	// lsu.scala:210:16
        ldq_6_bits_uop_debug_tsrc = _RANDOM[10'h71][27:26];	// lsu.scala:210:16
        ldq_6_bits_addr_valid = _RANDOM[10'h71][28];	// lsu.scala:210:16
        ldq_6_bits_addr_bits =
          {_RANDOM[10'h71][31:29], _RANDOM[10'h72], _RANDOM[10'h73][4:0]};	// lsu.scala:210:16
        ldq_6_bits_addr_is_virtual = _RANDOM[10'h73][5];	// lsu.scala:210:16
        ldq_6_bits_addr_is_uncacheable = _RANDOM[10'h73][6];	// lsu.scala:210:16
        ldq_6_bits_executed = _RANDOM[10'h73][7];	// lsu.scala:210:16
        ldq_6_bits_succeeded = _RANDOM[10'h73][8];	// lsu.scala:210:16
        ldq_6_bits_order_fail = _RANDOM[10'h73][9];	// lsu.scala:210:16
        ldq_6_bits_observed = _RANDOM[10'h73][10];	// lsu.scala:210:16
        ldq_6_bits_st_dep_mask = _RANDOM[10'h73][26:11];	// lsu.scala:210:16
        ldq_6_bits_youngest_stq_idx = _RANDOM[10'h73][30:27];	// lsu.scala:210:16
        ldq_6_bits_forward_std_val = _RANDOM[10'h73][31];	// lsu.scala:210:16
        ldq_6_bits_forward_stq_idx = _RANDOM[10'h74][3:0];	// lsu.scala:210:16
        ldq_7_valid = _RANDOM[10'h76][4];	// lsu.scala:210:16
        ldq_7_bits_uop_uopc = _RANDOM[10'h76][11:5];	// lsu.scala:210:16
        ldq_7_bits_uop_inst = {_RANDOM[10'h76][31:12], _RANDOM[10'h77][11:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_debug_inst = {_RANDOM[10'h77][31:12], _RANDOM[10'h78][11:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_is_rvc = _RANDOM[10'h78][12];	// lsu.scala:210:16
        ldq_7_bits_uop_debug_pc = {_RANDOM[10'h78][31:13], _RANDOM[10'h79][20:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_iq_type = _RANDOM[10'h79][23:21];	// lsu.scala:210:16
        ldq_7_bits_uop_fu_code = {_RANDOM[10'h79][31:24], _RANDOM[10'h7A][1:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_br_type = _RANDOM[10'h7A][5:2];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_op1_sel = _RANDOM[10'h7A][7:6];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_op2_sel = _RANDOM[10'h7A][10:8];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_imm_sel = _RANDOM[10'h7A][13:11];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_op_fcn = _RANDOM[10'h7A][17:14];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_fcn_dw = _RANDOM[10'h7A][18];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_csr_cmd = _RANDOM[10'h7A][21:19];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_is_load = _RANDOM[10'h7A][22];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_is_sta = _RANDOM[10'h7A][23];	// lsu.scala:210:16
        ldq_7_bits_uop_ctrl_is_std = _RANDOM[10'h7A][24];	// lsu.scala:210:16
        ldq_7_bits_uop_iw_state = _RANDOM[10'h7A][26:25];	// lsu.scala:210:16
        ldq_7_bits_uop_iw_p1_poisoned = _RANDOM[10'h7A][27];	// lsu.scala:210:16
        ldq_7_bits_uop_iw_p2_poisoned = _RANDOM[10'h7A][28];	// lsu.scala:210:16
        ldq_7_bits_uop_is_br = _RANDOM[10'h7A][29];	// lsu.scala:210:16
        ldq_7_bits_uop_is_jalr = _RANDOM[10'h7A][30];	// lsu.scala:210:16
        ldq_7_bits_uop_is_jal = _RANDOM[10'h7A][31];	// lsu.scala:210:16
        ldq_7_bits_uop_is_sfb = _RANDOM[10'h7B][0];	// lsu.scala:210:16
        ldq_7_bits_uop_br_mask = _RANDOM[10'h7B][12:1];	// lsu.scala:210:16
        ldq_7_bits_uop_br_tag = _RANDOM[10'h7B][16:13];	// lsu.scala:210:16
        ldq_7_bits_uop_ftq_idx = _RANDOM[10'h7B][21:17];	// lsu.scala:210:16
        ldq_7_bits_uop_edge_inst = _RANDOM[10'h7B][22];	// lsu.scala:210:16
        ldq_7_bits_uop_pc_lob = _RANDOM[10'h7B][28:23];	// lsu.scala:210:16
        ldq_7_bits_uop_taken = _RANDOM[10'h7B][29];	// lsu.scala:210:16
        ldq_7_bits_uop_imm_packed = {_RANDOM[10'h7B][31:30], _RANDOM[10'h7C][17:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_csr_addr = _RANDOM[10'h7C][29:18];	// lsu.scala:210:16
        ldq_7_bits_uop_rob_idx = {_RANDOM[10'h7C][31:30], _RANDOM[10'h7D][3:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_ldq_idx = _RANDOM[10'h7D][7:4];	// lsu.scala:210:16
        ldq_7_bits_uop_stq_idx = _RANDOM[10'h7D][11:8];	// lsu.scala:210:16
        ldq_7_bits_uop_rxq_idx = _RANDOM[10'h7D][13:12];	// lsu.scala:210:16
        ldq_7_bits_uop_pdst = _RANDOM[10'h7D][20:14];	// lsu.scala:210:16
        ldq_7_bits_uop_prs1 = _RANDOM[10'h7D][27:21];	// lsu.scala:210:16
        ldq_7_bits_uop_prs2 = {_RANDOM[10'h7D][31:28], _RANDOM[10'h7E][2:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_prs3 = _RANDOM[10'h7E][9:3];	// lsu.scala:210:16
        ldq_7_bits_uop_ppred = _RANDOM[10'h7E][14:10];	// lsu.scala:210:16
        ldq_7_bits_uop_prs1_busy = _RANDOM[10'h7E][15];	// lsu.scala:210:16
        ldq_7_bits_uop_prs2_busy = _RANDOM[10'h7E][16];	// lsu.scala:210:16
        ldq_7_bits_uop_prs3_busy = _RANDOM[10'h7E][17];	// lsu.scala:210:16
        ldq_7_bits_uop_ppred_busy = _RANDOM[10'h7E][18];	// lsu.scala:210:16
        ldq_7_bits_uop_stale_pdst = _RANDOM[10'h7E][25:19];	// lsu.scala:210:16
        ldq_7_bits_uop_exception = _RANDOM[10'h7E][26];	// lsu.scala:210:16
        ldq_7_bits_uop_exc_cause =
          {_RANDOM[10'h7E][31:27], _RANDOM[10'h7F], _RANDOM[10'h80][26:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_bypassable = _RANDOM[10'h80][27];	// lsu.scala:210:16
        ldq_7_bits_uop_mem_cmd = {_RANDOM[10'h80][31:28], _RANDOM[10'h81][0]};	// lsu.scala:210:16
        ldq_7_bits_uop_mem_size = _RANDOM[10'h81][2:1];	// lsu.scala:210:16
        ldq_7_bits_uop_mem_signed = _RANDOM[10'h81][3];	// lsu.scala:210:16
        ldq_7_bits_uop_is_fence = _RANDOM[10'h81][4];	// lsu.scala:210:16
        ldq_7_bits_uop_is_fencei = _RANDOM[10'h81][5];	// lsu.scala:210:16
        ldq_7_bits_uop_is_amo = _RANDOM[10'h81][6];	// lsu.scala:210:16
        ldq_7_bits_uop_uses_ldq = _RANDOM[10'h81][7];	// lsu.scala:210:16
        ldq_7_bits_uop_uses_stq = _RANDOM[10'h81][8];	// lsu.scala:210:16
        ldq_7_bits_uop_is_sys_pc2epc = _RANDOM[10'h81][9];	// lsu.scala:210:16
        ldq_7_bits_uop_is_unique = _RANDOM[10'h81][10];	// lsu.scala:210:16
        ldq_7_bits_uop_flush_on_commit = _RANDOM[10'h81][11];	// lsu.scala:210:16
        ldq_7_bits_uop_ldst_is_rs1 = _RANDOM[10'h81][12];	// lsu.scala:210:16
        ldq_7_bits_uop_ldst = _RANDOM[10'h81][18:13];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs1 = _RANDOM[10'h81][24:19];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs2 = _RANDOM[10'h81][30:25];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs3 = {_RANDOM[10'h81][31], _RANDOM[10'h82][4:0]};	// lsu.scala:210:16
        ldq_7_bits_uop_ldst_val = _RANDOM[10'h82][5];	// lsu.scala:210:16
        ldq_7_bits_uop_dst_rtype = _RANDOM[10'h82][7:6];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs1_rtype = _RANDOM[10'h82][9:8];	// lsu.scala:210:16
        ldq_7_bits_uop_lrs2_rtype = _RANDOM[10'h82][11:10];	// lsu.scala:210:16
        ldq_7_bits_uop_frs3_en = _RANDOM[10'h82][12];	// lsu.scala:210:16
        ldq_7_bits_uop_fp_val = _RANDOM[10'h82][13];	// lsu.scala:210:16
        ldq_7_bits_uop_fp_single = _RANDOM[10'h82][14];	// lsu.scala:210:16
        ldq_7_bits_uop_xcpt_pf_if = _RANDOM[10'h82][15];	// lsu.scala:210:16
        ldq_7_bits_uop_xcpt_ae_if = _RANDOM[10'h82][16];	// lsu.scala:210:16
        ldq_7_bits_uop_xcpt_ma_if = _RANDOM[10'h82][17];	// lsu.scala:210:16
        ldq_7_bits_uop_bp_debug_if = _RANDOM[10'h82][18];	// lsu.scala:210:16
        ldq_7_bits_uop_bp_xcpt_if = _RANDOM[10'h82][19];	// lsu.scala:210:16
        ldq_7_bits_uop_debug_fsrc = _RANDOM[10'h82][21:20];	// lsu.scala:210:16
        ldq_7_bits_uop_debug_tsrc = _RANDOM[10'h82][23:22];	// lsu.scala:210:16
        ldq_7_bits_addr_valid = _RANDOM[10'h82][24];	// lsu.scala:210:16
        ldq_7_bits_addr_bits =
          {_RANDOM[10'h82][31:25], _RANDOM[10'h83], _RANDOM[10'h84][0]};	// lsu.scala:210:16
        ldq_7_bits_addr_is_virtual = _RANDOM[10'h84][1];	// lsu.scala:210:16
        ldq_7_bits_addr_is_uncacheable = _RANDOM[10'h84][2];	// lsu.scala:210:16
        ldq_7_bits_executed = _RANDOM[10'h84][3];	// lsu.scala:210:16
        ldq_7_bits_succeeded = _RANDOM[10'h84][4];	// lsu.scala:210:16
        ldq_7_bits_order_fail = _RANDOM[10'h84][5];	// lsu.scala:210:16
        ldq_7_bits_observed = _RANDOM[10'h84][6];	// lsu.scala:210:16
        ldq_7_bits_st_dep_mask = _RANDOM[10'h84][22:7];	// lsu.scala:210:16
        ldq_7_bits_youngest_stq_idx = _RANDOM[10'h84][26:23];	// lsu.scala:210:16
        ldq_7_bits_forward_std_val = _RANDOM[10'h84][27];	// lsu.scala:210:16
        ldq_7_bits_forward_stq_idx = _RANDOM[10'h84][31:28];	// lsu.scala:210:16
        ldq_8_valid = _RANDOM[10'h87][0];	// lsu.scala:210:16
        ldq_8_bits_uop_uopc = _RANDOM[10'h87][7:1];	// lsu.scala:210:16
        ldq_8_bits_uop_inst = {_RANDOM[10'h87][31:8], _RANDOM[10'h88][7:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_debug_inst = {_RANDOM[10'h88][31:8], _RANDOM[10'h89][7:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_is_rvc = _RANDOM[10'h89][8];	// lsu.scala:210:16
        ldq_8_bits_uop_debug_pc = {_RANDOM[10'h89][31:9], _RANDOM[10'h8A][16:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_iq_type = _RANDOM[10'h8A][19:17];	// lsu.scala:210:16
        ldq_8_bits_uop_fu_code = _RANDOM[10'h8A][29:20];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_br_type = {_RANDOM[10'h8A][31:30], _RANDOM[10'h8B][1:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_op1_sel = _RANDOM[10'h8B][3:2];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_op2_sel = _RANDOM[10'h8B][6:4];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_imm_sel = _RANDOM[10'h8B][9:7];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_op_fcn = _RANDOM[10'h8B][13:10];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_fcn_dw = _RANDOM[10'h8B][14];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_csr_cmd = _RANDOM[10'h8B][17:15];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_is_load = _RANDOM[10'h8B][18];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_is_sta = _RANDOM[10'h8B][19];	// lsu.scala:210:16
        ldq_8_bits_uop_ctrl_is_std = _RANDOM[10'h8B][20];	// lsu.scala:210:16
        ldq_8_bits_uop_iw_state = _RANDOM[10'h8B][22:21];	// lsu.scala:210:16
        ldq_8_bits_uop_iw_p1_poisoned = _RANDOM[10'h8B][23];	// lsu.scala:210:16
        ldq_8_bits_uop_iw_p2_poisoned = _RANDOM[10'h8B][24];	// lsu.scala:210:16
        ldq_8_bits_uop_is_br = _RANDOM[10'h8B][25];	// lsu.scala:210:16
        ldq_8_bits_uop_is_jalr = _RANDOM[10'h8B][26];	// lsu.scala:210:16
        ldq_8_bits_uop_is_jal = _RANDOM[10'h8B][27];	// lsu.scala:210:16
        ldq_8_bits_uop_is_sfb = _RANDOM[10'h8B][28];	// lsu.scala:210:16
        ldq_8_bits_uop_br_mask = {_RANDOM[10'h8B][31:29], _RANDOM[10'h8C][8:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_br_tag = _RANDOM[10'h8C][12:9];	// lsu.scala:210:16
        ldq_8_bits_uop_ftq_idx = _RANDOM[10'h8C][17:13];	// lsu.scala:210:16
        ldq_8_bits_uop_edge_inst = _RANDOM[10'h8C][18];	// lsu.scala:210:16
        ldq_8_bits_uop_pc_lob = _RANDOM[10'h8C][24:19];	// lsu.scala:210:16
        ldq_8_bits_uop_taken = _RANDOM[10'h8C][25];	// lsu.scala:210:16
        ldq_8_bits_uop_imm_packed = {_RANDOM[10'h8C][31:26], _RANDOM[10'h8D][13:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_csr_addr = _RANDOM[10'h8D][25:14];	// lsu.scala:210:16
        ldq_8_bits_uop_rob_idx = _RANDOM[10'h8D][31:26];	// lsu.scala:210:16
        ldq_8_bits_uop_ldq_idx = _RANDOM[10'h8E][3:0];	// lsu.scala:210:16
        ldq_8_bits_uop_stq_idx = _RANDOM[10'h8E][7:4];	// lsu.scala:210:16
        ldq_8_bits_uop_rxq_idx = _RANDOM[10'h8E][9:8];	// lsu.scala:210:16
        ldq_8_bits_uop_pdst = _RANDOM[10'h8E][16:10];	// lsu.scala:210:16
        ldq_8_bits_uop_prs1 = _RANDOM[10'h8E][23:17];	// lsu.scala:210:16
        ldq_8_bits_uop_prs2 = _RANDOM[10'h8E][30:24];	// lsu.scala:210:16
        ldq_8_bits_uop_prs3 = {_RANDOM[10'h8E][31], _RANDOM[10'h8F][5:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_ppred = _RANDOM[10'h8F][10:6];	// lsu.scala:210:16
        ldq_8_bits_uop_prs1_busy = _RANDOM[10'h8F][11];	// lsu.scala:210:16
        ldq_8_bits_uop_prs2_busy = _RANDOM[10'h8F][12];	// lsu.scala:210:16
        ldq_8_bits_uop_prs3_busy = _RANDOM[10'h8F][13];	// lsu.scala:210:16
        ldq_8_bits_uop_ppred_busy = _RANDOM[10'h8F][14];	// lsu.scala:210:16
        ldq_8_bits_uop_stale_pdst = _RANDOM[10'h8F][21:15];	// lsu.scala:210:16
        ldq_8_bits_uop_exception = _RANDOM[10'h8F][22];	// lsu.scala:210:16
        ldq_8_bits_uop_exc_cause =
          {_RANDOM[10'h8F][31:23], _RANDOM[10'h90], _RANDOM[10'h91][22:0]};	// lsu.scala:210:16
        ldq_8_bits_uop_bypassable = _RANDOM[10'h91][23];	// lsu.scala:210:16
        ldq_8_bits_uop_mem_cmd = _RANDOM[10'h91][28:24];	// lsu.scala:210:16
        ldq_8_bits_uop_mem_size = _RANDOM[10'h91][30:29];	// lsu.scala:210:16
        ldq_8_bits_uop_mem_signed = _RANDOM[10'h91][31];	// lsu.scala:210:16
        ldq_8_bits_uop_is_fence = _RANDOM[10'h92][0];	// lsu.scala:210:16
        ldq_8_bits_uop_is_fencei = _RANDOM[10'h92][1];	// lsu.scala:210:16
        ldq_8_bits_uop_is_amo = _RANDOM[10'h92][2];	// lsu.scala:210:16
        ldq_8_bits_uop_uses_ldq = _RANDOM[10'h92][3];	// lsu.scala:210:16
        ldq_8_bits_uop_uses_stq = _RANDOM[10'h92][4];	// lsu.scala:210:16
        ldq_8_bits_uop_is_sys_pc2epc = _RANDOM[10'h92][5];	// lsu.scala:210:16
        ldq_8_bits_uop_is_unique = _RANDOM[10'h92][6];	// lsu.scala:210:16
        ldq_8_bits_uop_flush_on_commit = _RANDOM[10'h92][7];	// lsu.scala:210:16
        ldq_8_bits_uop_ldst_is_rs1 = _RANDOM[10'h92][8];	// lsu.scala:210:16
        ldq_8_bits_uop_ldst = _RANDOM[10'h92][14:9];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs1 = _RANDOM[10'h92][20:15];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs2 = _RANDOM[10'h92][26:21];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs3 = {_RANDOM[10'h92][31:27], _RANDOM[10'h93][0]};	// lsu.scala:210:16
        ldq_8_bits_uop_ldst_val = _RANDOM[10'h93][1];	// lsu.scala:210:16
        ldq_8_bits_uop_dst_rtype = _RANDOM[10'h93][3:2];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs1_rtype = _RANDOM[10'h93][5:4];	// lsu.scala:210:16
        ldq_8_bits_uop_lrs2_rtype = _RANDOM[10'h93][7:6];	// lsu.scala:210:16
        ldq_8_bits_uop_frs3_en = _RANDOM[10'h93][8];	// lsu.scala:210:16
        ldq_8_bits_uop_fp_val = _RANDOM[10'h93][9];	// lsu.scala:210:16
        ldq_8_bits_uop_fp_single = _RANDOM[10'h93][10];	// lsu.scala:210:16
        ldq_8_bits_uop_xcpt_pf_if = _RANDOM[10'h93][11];	// lsu.scala:210:16
        ldq_8_bits_uop_xcpt_ae_if = _RANDOM[10'h93][12];	// lsu.scala:210:16
        ldq_8_bits_uop_xcpt_ma_if = _RANDOM[10'h93][13];	// lsu.scala:210:16
        ldq_8_bits_uop_bp_debug_if = _RANDOM[10'h93][14];	// lsu.scala:210:16
        ldq_8_bits_uop_bp_xcpt_if = _RANDOM[10'h93][15];	// lsu.scala:210:16
        ldq_8_bits_uop_debug_fsrc = _RANDOM[10'h93][17:16];	// lsu.scala:210:16
        ldq_8_bits_uop_debug_tsrc = _RANDOM[10'h93][19:18];	// lsu.scala:210:16
        ldq_8_bits_addr_valid = _RANDOM[10'h93][20];	// lsu.scala:210:16
        ldq_8_bits_addr_bits = {_RANDOM[10'h93][31:21], _RANDOM[10'h94][28:0]};	// lsu.scala:210:16
        ldq_8_bits_addr_is_virtual = _RANDOM[10'h94][29];	// lsu.scala:210:16
        ldq_8_bits_addr_is_uncacheable = _RANDOM[10'h94][30];	// lsu.scala:210:16
        ldq_8_bits_executed = _RANDOM[10'h94][31];	// lsu.scala:210:16
        ldq_8_bits_succeeded = _RANDOM[10'h95][0];	// lsu.scala:210:16
        ldq_8_bits_order_fail = _RANDOM[10'h95][1];	// lsu.scala:210:16
        ldq_8_bits_observed = _RANDOM[10'h95][2];	// lsu.scala:210:16
        ldq_8_bits_st_dep_mask = _RANDOM[10'h95][18:3];	// lsu.scala:210:16
        ldq_8_bits_youngest_stq_idx = _RANDOM[10'h95][22:19];	// lsu.scala:210:16
        ldq_8_bits_forward_std_val = _RANDOM[10'h95][23];	// lsu.scala:210:16
        ldq_8_bits_forward_stq_idx = _RANDOM[10'h95][27:24];	// lsu.scala:210:16
        ldq_9_valid = _RANDOM[10'h97][28];	// lsu.scala:210:16
        ldq_9_bits_uop_uopc = {_RANDOM[10'h97][31:29], _RANDOM[10'h98][3:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_inst = {_RANDOM[10'h98][31:4], _RANDOM[10'h99][3:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_debug_inst = {_RANDOM[10'h99][31:4], _RANDOM[10'h9A][3:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_is_rvc = _RANDOM[10'h9A][4];	// lsu.scala:210:16
        ldq_9_bits_uop_debug_pc = {_RANDOM[10'h9A][31:5], _RANDOM[10'h9B][12:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_iq_type = _RANDOM[10'h9B][15:13];	// lsu.scala:210:16
        ldq_9_bits_uop_fu_code = _RANDOM[10'h9B][25:16];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_br_type = _RANDOM[10'h9B][29:26];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_op1_sel = _RANDOM[10'h9B][31:30];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_op2_sel = _RANDOM[10'h9C][2:0];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_imm_sel = _RANDOM[10'h9C][5:3];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_op_fcn = _RANDOM[10'h9C][9:6];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_fcn_dw = _RANDOM[10'h9C][10];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_csr_cmd = _RANDOM[10'h9C][13:11];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_is_load = _RANDOM[10'h9C][14];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_is_sta = _RANDOM[10'h9C][15];	// lsu.scala:210:16
        ldq_9_bits_uop_ctrl_is_std = _RANDOM[10'h9C][16];	// lsu.scala:210:16
        ldq_9_bits_uop_iw_state = _RANDOM[10'h9C][18:17];	// lsu.scala:210:16
        ldq_9_bits_uop_iw_p1_poisoned = _RANDOM[10'h9C][19];	// lsu.scala:210:16
        ldq_9_bits_uop_iw_p2_poisoned = _RANDOM[10'h9C][20];	// lsu.scala:210:16
        ldq_9_bits_uop_is_br = _RANDOM[10'h9C][21];	// lsu.scala:210:16
        ldq_9_bits_uop_is_jalr = _RANDOM[10'h9C][22];	// lsu.scala:210:16
        ldq_9_bits_uop_is_jal = _RANDOM[10'h9C][23];	// lsu.scala:210:16
        ldq_9_bits_uop_is_sfb = _RANDOM[10'h9C][24];	// lsu.scala:210:16
        ldq_9_bits_uop_br_mask = {_RANDOM[10'h9C][31:25], _RANDOM[10'h9D][4:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_br_tag = _RANDOM[10'h9D][8:5];	// lsu.scala:210:16
        ldq_9_bits_uop_ftq_idx = _RANDOM[10'h9D][13:9];	// lsu.scala:210:16
        ldq_9_bits_uop_edge_inst = _RANDOM[10'h9D][14];	// lsu.scala:210:16
        ldq_9_bits_uop_pc_lob = _RANDOM[10'h9D][20:15];	// lsu.scala:210:16
        ldq_9_bits_uop_taken = _RANDOM[10'h9D][21];	// lsu.scala:210:16
        ldq_9_bits_uop_imm_packed = {_RANDOM[10'h9D][31:22], _RANDOM[10'h9E][9:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_csr_addr = _RANDOM[10'h9E][21:10];	// lsu.scala:210:16
        ldq_9_bits_uop_rob_idx = _RANDOM[10'h9E][27:22];	// lsu.scala:210:16
        ldq_9_bits_uop_ldq_idx = _RANDOM[10'h9E][31:28];	// lsu.scala:210:16
        ldq_9_bits_uop_stq_idx = _RANDOM[10'h9F][3:0];	// lsu.scala:210:16
        ldq_9_bits_uop_rxq_idx = _RANDOM[10'h9F][5:4];	// lsu.scala:210:16
        ldq_9_bits_uop_pdst = _RANDOM[10'h9F][12:6];	// lsu.scala:210:16
        ldq_9_bits_uop_prs1 = _RANDOM[10'h9F][19:13];	// lsu.scala:210:16
        ldq_9_bits_uop_prs2 = _RANDOM[10'h9F][26:20];	// lsu.scala:210:16
        ldq_9_bits_uop_prs3 = {_RANDOM[10'h9F][31:27], _RANDOM[10'hA0][1:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_ppred = _RANDOM[10'hA0][6:2];	// lsu.scala:210:16
        ldq_9_bits_uop_prs1_busy = _RANDOM[10'hA0][7];	// lsu.scala:210:16
        ldq_9_bits_uop_prs2_busy = _RANDOM[10'hA0][8];	// lsu.scala:210:16
        ldq_9_bits_uop_prs3_busy = _RANDOM[10'hA0][9];	// lsu.scala:210:16
        ldq_9_bits_uop_ppred_busy = _RANDOM[10'hA0][10];	// lsu.scala:210:16
        ldq_9_bits_uop_stale_pdst = _RANDOM[10'hA0][17:11];	// lsu.scala:210:16
        ldq_9_bits_uop_exception = _RANDOM[10'hA0][18];	// lsu.scala:210:16
        ldq_9_bits_uop_exc_cause =
          {_RANDOM[10'hA0][31:19], _RANDOM[10'hA1], _RANDOM[10'hA2][18:0]};	// lsu.scala:210:16
        ldq_9_bits_uop_bypassable = _RANDOM[10'hA2][19];	// lsu.scala:210:16
        ldq_9_bits_uop_mem_cmd = _RANDOM[10'hA2][24:20];	// lsu.scala:210:16
        ldq_9_bits_uop_mem_size = _RANDOM[10'hA2][26:25];	// lsu.scala:210:16
        ldq_9_bits_uop_mem_signed = _RANDOM[10'hA2][27];	// lsu.scala:210:16
        ldq_9_bits_uop_is_fence = _RANDOM[10'hA2][28];	// lsu.scala:210:16
        ldq_9_bits_uop_is_fencei = _RANDOM[10'hA2][29];	// lsu.scala:210:16
        ldq_9_bits_uop_is_amo = _RANDOM[10'hA2][30];	// lsu.scala:210:16
        ldq_9_bits_uop_uses_ldq = _RANDOM[10'hA2][31];	// lsu.scala:210:16
        ldq_9_bits_uop_uses_stq = _RANDOM[10'hA3][0];	// lsu.scala:210:16
        ldq_9_bits_uop_is_sys_pc2epc = _RANDOM[10'hA3][1];	// lsu.scala:210:16
        ldq_9_bits_uop_is_unique = _RANDOM[10'hA3][2];	// lsu.scala:210:16
        ldq_9_bits_uop_flush_on_commit = _RANDOM[10'hA3][3];	// lsu.scala:210:16
        ldq_9_bits_uop_ldst_is_rs1 = _RANDOM[10'hA3][4];	// lsu.scala:210:16
        ldq_9_bits_uop_ldst = _RANDOM[10'hA3][10:5];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs1 = _RANDOM[10'hA3][16:11];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs2 = _RANDOM[10'hA3][22:17];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs3 = _RANDOM[10'hA3][28:23];	// lsu.scala:210:16
        ldq_9_bits_uop_ldst_val = _RANDOM[10'hA3][29];	// lsu.scala:210:16
        ldq_9_bits_uop_dst_rtype = _RANDOM[10'hA3][31:30];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs1_rtype = _RANDOM[10'hA4][1:0];	// lsu.scala:210:16
        ldq_9_bits_uop_lrs2_rtype = _RANDOM[10'hA4][3:2];	// lsu.scala:210:16
        ldq_9_bits_uop_frs3_en = _RANDOM[10'hA4][4];	// lsu.scala:210:16
        ldq_9_bits_uop_fp_val = _RANDOM[10'hA4][5];	// lsu.scala:210:16
        ldq_9_bits_uop_fp_single = _RANDOM[10'hA4][6];	// lsu.scala:210:16
        ldq_9_bits_uop_xcpt_pf_if = _RANDOM[10'hA4][7];	// lsu.scala:210:16
        ldq_9_bits_uop_xcpt_ae_if = _RANDOM[10'hA4][8];	// lsu.scala:210:16
        ldq_9_bits_uop_xcpt_ma_if = _RANDOM[10'hA4][9];	// lsu.scala:210:16
        ldq_9_bits_uop_bp_debug_if = _RANDOM[10'hA4][10];	// lsu.scala:210:16
        ldq_9_bits_uop_bp_xcpt_if = _RANDOM[10'hA4][11];	// lsu.scala:210:16
        ldq_9_bits_uop_debug_fsrc = _RANDOM[10'hA4][13:12];	// lsu.scala:210:16
        ldq_9_bits_uop_debug_tsrc = _RANDOM[10'hA4][15:14];	// lsu.scala:210:16
        ldq_9_bits_addr_valid = _RANDOM[10'hA4][16];	// lsu.scala:210:16
        ldq_9_bits_addr_bits = {_RANDOM[10'hA4][31:17], _RANDOM[10'hA5][24:0]};	// lsu.scala:210:16
        ldq_9_bits_addr_is_virtual = _RANDOM[10'hA5][25];	// lsu.scala:210:16
        ldq_9_bits_addr_is_uncacheable = _RANDOM[10'hA5][26];	// lsu.scala:210:16
        ldq_9_bits_executed = _RANDOM[10'hA5][27];	// lsu.scala:210:16
        ldq_9_bits_succeeded = _RANDOM[10'hA5][28];	// lsu.scala:210:16
        ldq_9_bits_order_fail = _RANDOM[10'hA5][29];	// lsu.scala:210:16
        ldq_9_bits_observed = _RANDOM[10'hA5][30];	// lsu.scala:210:16
        ldq_9_bits_st_dep_mask = {_RANDOM[10'hA5][31], _RANDOM[10'hA6][14:0]};	// lsu.scala:210:16
        ldq_9_bits_youngest_stq_idx = _RANDOM[10'hA6][18:15];	// lsu.scala:210:16
        ldq_9_bits_forward_std_val = _RANDOM[10'hA6][19];	// lsu.scala:210:16
        ldq_9_bits_forward_stq_idx = _RANDOM[10'hA6][23:20];	// lsu.scala:210:16
        ldq_10_valid = _RANDOM[10'hA8][24];	// lsu.scala:210:16
        ldq_10_bits_uop_uopc = _RANDOM[10'hA8][31:25];	// lsu.scala:210:16
        ldq_10_bits_uop_inst = _RANDOM[10'hA9];	// lsu.scala:210:16
        ldq_10_bits_uop_debug_inst = _RANDOM[10'hAA];	// lsu.scala:210:16
        ldq_10_bits_uop_is_rvc = _RANDOM[10'hAB][0];	// lsu.scala:210:16
        ldq_10_bits_uop_debug_pc = {_RANDOM[10'hAB][31:1], _RANDOM[10'hAC][8:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_iq_type = _RANDOM[10'hAC][11:9];	// lsu.scala:210:16
        ldq_10_bits_uop_fu_code = _RANDOM[10'hAC][21:12];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_br_type = _RANDOM[10'hAC][25:22];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_op1_sel = _RANDOM[10'hAC][27:26];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_op2_sel = _RANDOM[10'hAC][30:28];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_imm_sel = {_RANDOM[10'hAC][31], _RANDOM[10'hAD][1:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_op_fcn = _RANDOM[10'hAD][5:2];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_fcn_dw = _RANDOM[10'hAD][6];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_csr_cmd = _RANDOM[10'hAD][9:7];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_is_load = _RANDOM[10'hAD][10];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_is_sta = _RANDOM[10'hAD][11];	// lsu.scala:210:16
        ldq_10_bits_uop_ctrl_is_std = _RANDOM[10'hAD][12];	// lsu.scala:210:16
        ldq_10_bits_uop_iw_state = _RANDOM[10'hAD][14:13];	// lsu.scala:210:16
        ldq_10_bits_uop_iw_p1_poisoned = _RANDOM[10'hAD][15];	// lsu.scala:210:16
        ldq_10_bits_uop_iw_p2_poisoned = _RANDOM[10'hAD][16];	// lsu.scala:210:16
        ldq_10_bits_uop_is_br = _RANDOM[10'hAD][17];	// lsu.scala:210:16
        ldq_10_bits_uop_is_jalr = _RANDOM[10'hAD][18];	// lsu.scala:210:16
        ldq_10_bits_uop_is_jal = _RANDOM[10'hAD][19];	// lsu.scala:210:16
        ldq_10_bits_uop_is_sfb = _RANDOM[10'hAD][20];	// lsu.scala:210:16
        ldq_10_bits_uop_br_mask = {_RANDOM[10'hAD][31:21], _RANDOM[10'hAE][0]};	// lsu.scala:210:16
        ldq_10_bits_uop_br_tag = _RANDOM[10'hAE][4:1];	// lsu.scala:210:16
        ldq_10_bits_uop_ftq_idx = _RANDOM[10'hAE][9:5];	// lsu.scala:210:16
        ldq_10_bits_uop_edge_inst = _RANDOM[10'hAE][10];	// lsu.scala:210:16
        ldq_10_bits_uop_pc_lob = _RANDOM[10'hAE][16:11];	// lsu.scala:210:16
        ldq_10_bits_uop_taken = _RANDOM[10'hAE][17];	// lsu.scala:210:16
        ldq_10_bits_uop_imm_packed = {_RANDOM[10'hAE][31:18], _RANDOM[10'hAF][5:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_csr_addr = _RANDOM[10'hAF][17:6];	// lsu.scala:210:16
        ldq_10_bits_uop_rob_idx = _RANDOM[10'hAF][23:18];	// lsu.scala:210:16
        ldq_10_bits_uop_ldq_idx = _RANDOM[10'hAF][27:24];	// lsu.scala:210:16
        ldq_10_bits_uop_stq_idx = _RANDOM[10'hAF][31:28];	// lsu.scala:210:16
        ldq_10_bits_uop_rxq_idx = _RANDOM[10'hB0][1:0];	// lsu.scala:210:16
        ldq_10_bits_uop_pdst = _RANDOM[10'hB0][8:2];	// lsu.scala:210:16
        ldq_10_bits_uop_prs1 = _RANDOM[10'hB0][15:9];	// lsu.scala:210:16
        ldq_10_bits_uop_prs2 = _RANDOM[10'hB0][22:16];	// lsu.scala:210:16
        ldq_10_bits_uop_prs3 = _RANDOM[10'hB0][29:23];	// lsu.scala:210:16
        ldq_10_bits_uop_ppred = {_RANDOM[10'hB0][31:30], _RANDOM[10'hB1][2:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_prs1_busy = _RANDOM[10'hB1][3];	// lsu.scala:210:16
        ldq_10_bits_uop_prs2_busy = _RANDOM[10'hB1][4];	// lsu.scala:210:16
        ldq_10_bits_uop_prs3_busy = _RANDOM[10'hB1][5];	// lsu.scala:210:16
        ldq_10_bits_uop_ppred_busy = _RANDOM[10'hB1][6];	// lsu.scala:210:16
        ldq_10_bits_uop_stale_pdst = _RANDOM[10'hB1][13:7];	// lsu.scala:210:16
        ldq_10_bits_uop_exception = _RANDOM[10'hB1][14];	// lsu.scala:210:16
        ldq_10_bits_uop_exc_cause =
          {_RANDOM[10'hB1][31:15], _RANDOM[10'hB2], _RANDOM[10'hB3][14:0]};	// lsu.scala:210:16
        ldq_10_bits_uop_bypassable = _RANDOM[10'hB3][15];	// lsu.scala:210:16
        ldq_10_bits_uop_mem_cmd = _RANDOM[10'hB3][20:16];	// lsu.scala:210:16
        ldq_10_bits_uop_mem_size = _RANDOM[10'hB3][22:21];	// lsu.scala:210:16
        ldq_10_bits_uop_mem_signed = _RANDOM[10'hB3][23];	// lsu.scala:210:16
        ldq_10_bits_uop_is_fence = _RANDOM[10'hB3][24];	// lsu.scala:210:16
        ldq_10_bits_uop_is_fencei = _RANDOM[10'hB3][25];	// lsu.scala:210:16
        ldq_10_bits_uop_is_amo = _RANDOM[10'hB3][26];	// lsu.scala:210:16
        ldq_10_bits_uop_uses_ldq = _RANDOM[10'hB3][27];	// lsu.scala:210:16
        ldq_10_bits_uop_uses_stq = _RANDOM[10'hB3][28];	// lsu.scala:210:16
        ldq_10_bits_uop_is_sys_pc2epc = _RANDOM[10'hB3][29];	// lsu.scala:210:16
        ldq_10_bits_uop_is_unique = _RANDOM[10'hB3][30];	// lsu.scala:210:16
        ldq_10_bits_uop_flush_on_commit = _RANDOM[10'hB3][31];	// lsu.scala:210:16
        ldq_10_bits_uop_ldst_is_rs1 = _RANDOM[10'hB4][0];	// lsu.scala:210:16
        ldq_10_bits_uop_ldst = _RANDOM[10'hB4][6:1];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs1 = _RANDOM[10'hB4][12:7];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs2 = _RANDOM[10'hB4][18:13];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs3 = _RANDOM[10'hB4][24:19];	// lsu.scala:210:16
        ldq_10_bits_uop_ldst_val = _RANDOM[10'hB4][25];	// lsu.scala:210:16
        ldq_10_bits_uop_dst_rtype = _RANDOM[10'hB4][27:26];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs1_rtype = _RANDOM[10'hB4][29:28];	// lsu.scala:210:16
        ldq_10_bits_uop_lrs2_rtype = _RANDOM[10'hB4][31:30];	// lsu.scala:210:16
        ldq_10_bits_uop_frs3_en = _RANDOM[10'hB5][0];	// lsu.scala:210:16
        ldq_10_bits_uop_fp_val = _RANDOM[10'hB5][1];	// lsu.scala:210:16
        ldq_10_bits_uop_fp_single = _RANDOM[10'hB5][2];	// lsu.scala:210:16
        ldq_10_bits_uop_xcpt_pf_if = _RANDOM[10'hB5][3];	// lsu.scala:210:16
        ldq_10_bits_uop_xcpt_ae_if = _RANDOM[10'hB5][4];	// lsu.scala:210:16
        ldq_10_bits_uop_xcpt_ma_if = _RANDOM[10'hB5][5];	// lsu.scala:210:16
        ldq_10_bits_uop_bp_debug_if = _RANDOM[10'hB5][6];	// lsu.scala:210:16
        ldq_10_bits_uop_bp_xcpt_if = _RANDOM[10'hB5][7];	// lsu.scala:210:16
        ldq_10_bits_uop_debug_fsrc = _RANDOM[10'hB5][9:8];	// lsu.scala:210:16
        ldq_10_bits_uop_debug_tsrc = _RANDOM[10'hB5][11:10];	// lsu.scala:210:16
        ldq_10_bits_addr_valid = _RANDOM[10'hB5][12];	// lsu.scala:210:16
        ldq_10_bits_addr_bits = {_RANDOM[10'hB5][31:13], _RANDOM[10'hB6][20:0]};	// lsu.scala:210:16
        ldq_10_bits_addr_is_virtual = _RANDOM[10'hB6][21];	// lsu.scala:210:16
        ldq_10_bits_addr_is_uncacheable = _RANDOM[10'hB6][22];	// lsu.scala:210:16
        ldq_10_bits_executed = _RANDOM[10'hB6][23];	// lsu.scala:210:16
        ldq_10_bits_succeeded = _RANDOM[10'hB6][24];	// lsu.scala:210:16
        ldq_10_bits_order_fail = _RANDOM[10'hB6][25];	// lsu.scala:210:16
        ldq_10_bits_observed = _RANDOM[10'hB6][26];	// lsu.scala:210:16
        ldq_10_bits_st_dep_mask = {_RANDOM[10'hB6][31:27], _RANDOM[10'hB7][10:0]};	// lsu.scala:210:16
        ldq_10_bits_youngest_stq_idx = _RANDOM[10'hB7][14:11];	// lsu.scala:210:16
        ldq_10_bits_forward_std_val = _RANDOM[10'hB7][15];	// lsu.scala:210:16
        ldq_10_bits_forward_stq_idx = _RANDOM[10'hB7][19:16];	// lsu.scala:210:16
        ldq_11_valid = _RANDOM[10'hB9][20];	// lsu.scala:210:16
        ldq_11_bits_uop_uopc = _RANDOM[10'hB9][27:21];	// lsu.scala:210:16
        ldq_11_bits_uop_inst = {_RANDOM[10'hB9][31:28], _RANDOM[10'hBA][27:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_debug_inst = {_RANDOM[10'hBA][31:28], _RANDOM[10'hBB][27:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_is_rvc = _RANDOM[10'hBB][28];	// lsu.scala:210:16
        ldq_11_bits_uop_debug_pc =
          {_RANDOM[10'hBB][31:29], _RANDOM[10'hBC], _RANDOM[10'hBD][4:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_iq_type = _RANDOM[10'hBD][7:5];	// lsu.scala:210:16
        ldq_11_bits_uop_fu_code = _RANDOM[10'hBD][17:8];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_br_type = _RANDOM[10'hBD][21:18];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_op1_sel = _RANDOM[10'hBD][23:22];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_op2_sel = _RANDOM[10'hBD][26:24];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_imm_sel = _RANDOM[10'hBD][29:27];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_op_fcn = {_RANDOM[10'hBD][31:30], _RANDOM[10'hBE][1:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_fcn_dw = _RANDOM[10'hBE][2];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_csr_cmd = _RANDOM[10'hBE][5:3];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_is_load = _RANDOM[10'hBE][6];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_is_sta = _RANDOM[10'hBE][7];	// lsu.scala:210:16
        ldq_11_bits_uop_ctrl_is_std = _RANDOM[10'hBE][8];	// lsu.scala:210:16
        ldq_11_bits_uop_iw_state = _RANDOM[10'hBE][10:9];	// lsu.scala:210:16
        ldq_11_bits_uop_iw_p1_poisoned = _RANDOM[10'hBE][11];	// lsu.scala:210:16
        ldq_11_bits_uop_iw_p2_poisoned = _RANDOM[10'hBE][12];	// lsu.scala:210:16
        ldq_11_bits_uop_is_br = _RANDOM[10'hBE][13];	// lsu.scala:210:16
        ldq_11_bits_uop_is_jalr = _RANDOM[10'hBE][14];	// lsu.scala:210:16
        ldq_11_bits_uop_is_jal = _RANDOM[10'hBE][15];	// lsu.scala:210:16
        ldq_11_bits_uop_is_sfb = _RANDOM[10'hBE][16];	// lsu.scala:210:16
        ldq_11_bits_uop_br_mask = _RANDOM[10'hBE][28:17];	// lsu.scala:210:16
        ldq_11_bits_uop_br_tag = {_RANDOM[10'hBE][31:29], _RANDOM[10'hBF][0]};	// lsu.scala:210:16
        ldq_11_bits_uop_ftq_idx = _RANDOM[10'hBF][5:1];	// lsu.scala:210:16
        ldq_11_bits_uop_edge_inst = _RANDOM[10'hBF][6];	// lsu.scala:210:16
        ldq_11_bits_uop_pc_lob = _RANDOM[10'hBF][12:7];	// lsu.scala:210:16
        ldq_11_bits_uop_taken = _RANDOM[10'hBF][13];	// lsu.scala:210:16
        ldq_11_bits_uop_imm_packed = {_RANDOM[10'hBF][31:14], _RANDOM[10'hC0][1:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_csr_addr = _RANDOM[10'hC0][13:2];	// lsu.scala:210:16
        ldq_11_bits_uop_rob_idx = _RANDOM[10'hC0][19:14];	// lsu.scala:210:16
        ldq_11_bits_uop_ldq_idx = _RANDOM[10'hC0][23:20];	// lsu.scala:210:16
        ldq_11_bits_uop_stq_idx = _RANDOM[10'hC0][27:24];	// lsu.scala:210:16
        ldq_11_bits_uop_rxq_idx = _RANDOM[10'hC0][29:28];	// lsu.scala:210:16
        ldq_11_bits_uop_pdst = {_RANDOM[10'hC0][31:30], _RANDOM[10'hC1][4:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_prs1 = _RANDOM[10'hC1][11:5];	// lsu.scala:210:16
        ldq_11_bits_uop_prs2 = _RANDOM[10'hC1][18:12];	// lsu.scala:210:16
        ldq_11_bits_uop_prs3 = _RANDOM[10'hC1][25:19];	// lsu.scala:210:16
        ldq_11_bits_uop_ppred = _RANDOM[10'hC1][30:26];	// lsu.scala:210:16
        ldq_11_bits_uop_prs1_busy = _RANDOM[10'hC1][31];	// lsu.scala:210:16
        ldq_11_bits_uop_prs2_busy = _RANDOM[10'hC2][0];	// lsu.scala:210:16
        ldq_11_bits_uop_prs3_busy = _RANDOM[10'hC2][1];	// lsu.scala:210:16
        ldq_11_bits_uop_ppred_busy = _RANDOM[10'hC2][2];	// lsu.scala:210:16
        ldq_11_bits_uop_stale_pdst = _RANDOM[10'hC2][9:3];	// lsu.scala:210:16
        ldq_11_bits_uop_exception = _RANDOM[10'hC2][10];	// lsu.scala:210:16
        ldq_11_bits_uop_exc_cause =
          {_RANDOM[10'hC2][31:11], _RANDOM[10'hC3], _RANDOM[10'hC4][10:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_bypassable = _RANDOM[10'hC4][11];	// lsu.scala:210:16
        ldq_11_bits_uop_mem_cmd = _RANDOM[10'hC4][16:12];	// lsu.scala:210:16
        ldq_11_bits_uop_mem_size = _RANDOM[10'hC4][18:17];	// lsu.scala:210:16
        ldq_11_bits_uop_mem_signed = _RANDOM[10'hC4][19];	// lsu.scala:210:16
        ldq_11_bits_uop_is_fence = _RANDOM[10'hC4][20];	// lsu.scala:210:16
        ldq_11_bits_uop_is_fencei = _RANDOM[10'hC4][21];	// lsu.scala:210:16
        ldq_11_bits_uop_is_amo = _RANDOM[10'hC4][22];	// lsu.scala:210:16
        ldq_11_bits_uop_uses_ldq = _RANDOM[10'hC4][23];	// lsu.scala:210:16
        ldq_11_bits_uop_uses_stq = _RANDOM[10'hC4][24];	// lsu.scala:210:16
        ldq_11_bits_uop_is_sys_pc2epc = _RANDOM[10'hC4][25];	// lsu.scala:210:16
        ldq_11_bits_uop_is_unique = _RANDOM[10'hC4][26];	// lsu.scala:210:16
        ldq_11_bits_uop_flush_on_commit = _RANDOM[10'hC4][27];	// lsu.scala:210:16
        ldq_11_bits_uop_ldst_is_rs1 = _RANDOM[10'hC4][28];	// lsu.scala:210:16
        ldq_11_bits_uop_ldst = {_RANDOM[10'hC4][31:29], _RANDOM[10'hC5][2:0]};	// lsu.scala:210:16
        ldq_11_bits_uop_lrs1 = _RANDOM[10'hC5][8:3];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs2 = _RANDOM[10'hC5][14:9];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs3 = _RANDOM[10'hC5][20:15];	// lsu.scala:210:16
        ldq_11_bits_uop_ldst_val = _RANDOM[10'hC5][21];	// lsu.scala:210:16
        ldq_11_bits_uop_dst_rtype = _RANDOM[10'hC5][23:22];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs1_rtype = _RANDOM[10'hC5][25:24];	// lsu.scala:210:16
        ldq_11_bits_uop_lrs2_rtype = _RANDOM[10'hC5][27:26];	// lsu.scala:210:16
        ldq_11_bits_uop_frs3_en = _RANDOM[10'hC5][28];	// lsu.scala:210:16
        ldq_11_bits_uop_fp_val = _RANDOM[10'hC5][29];	// lsu.scala:210:16
        ldq_11_bits_uop_fp_single = _RANDOM[10'hC5][30];	// lsu.scala:210:16
        ldq_11_bits_uop_xcpt_pf_if = _RANDOM[10'hC5][31];	// lsu.scala:210:16
        ldq_11_bits_uop_xcpt_ae_if = _RANDOM[10'hC6][0];	// lsu.scala:210:16
        ldq_11_bits_uop_xcpt_ma_if = _RANDOM[10'hC6][1];	// lsu.scala:210:16
        ldq_11_bits_uop_bp_debug_if = _RANDOM[10'hC6][2];	// lsu.scala:210:16
        ldq_11_bits_uop_bp_xcpt_if = _RANDOM[10'hC6][3];	// lsu.scala:210:16
        ldq_11_bits_uop_debug_fsrc = _RANDOM[10'hC6][5:4];	// lsu.scala:210:16
        ldq_11_bits_uop_debug_tsrc = _RANDOM[10'hC6][7:6];	// lsu.scala:210:16
        ldq_11_bits_addr_valid = _RANDOM[10'hC6][8];	// lsu.scala:210:16
        ldq_11_bits_addr_bits = {_RANDOM[10'hC6][31:9], _RANDOM[10'hC7][16:0]};	// lsu.scala:210:16
        ldq_11_bits_addr_is_virtual = _RANDOM[10'hC7][17];	// lsu.scala:210:16
        ldq_11_bits_addr_is_uncacheable = _RANDOM[10'hC7][18];	// lsu.scala:210:16
        ldq_11_bits_executed = _RANDOM[10'hC7][19];	// lsu.scala:210:16
        ldq_11_bits_succeeded = _RANDOM[10'hC7][20];	// lsu.scala:210:16
        ldq_11_bits_order_fail = _RANDOM[10'hC7][21];	// lsu.scala:210:16
        ldq_11_bits_observed = _RANDOM[10'hC7][22];	// lsu.scala:210:16
        ldq_11_bits_st_dep_mask = {_RANDOM[10'hC7][31:23], _RANDOM[10'hC8][6:0]};	// lsu.scala:210:16
        ldq_11_bits_youngest_stq_idx = _RANDOM[10'hC8][10:7];	// lsu.scala:210:16
        ldq_11_bits_forward_std_val = _RANDOM[10'hC8][11];	// lsu.scala:210:16
        ldq_11_bits_forward_stq_idx = _RANDOM[10'hC8][15:12];	// lsu.scala:210:16
        ldq_12_valid = _RANDOM[10'hCA][16];	// lsu.scala:210:16
        ldq_12_bits_uop_uopc = _RANDOM[10'hCA][23:17];	// lsu.scala:210:16
        ldq_12_bits_uop_inst = {_RANDOM[10'hCA][31:24], _RANDOM[10'hCB][23:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_debug_inst = {_RANDOM[10'hCB][31:24], _RANDOM[10'hCC][23:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_is_rvc = _RANDOM[10'hCC][24];	// lsu.scala:210:16
        ldq_12_bits_uop_debug_pc =
          {_RANDOM[10'hCC][31:25], _RANDOM[10'hCD], _RANDOM[10'hCE][0]};	// lsu.scala:210:16
        ldq_12_bits_uop_iq_type = _RANDOM[10'hCE][3:1];	// lsu.scala:210:16
        ldq_12_bits_uop_fu_code = _RANDOM[10'hCE][13:4];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_br_type = _RANDOM[10'hCE][17:14];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_op1_sel = _RANDOM[10'hCE][19:18];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_op2_sel = _RANDOM[10'hCE][22:20];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_imm_sel = _RANDOM[10'hCE][25:23];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_op_fcn = _RANDOM[10'hCE][29:26];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_fcn_dw = _RANDOM[10'hCE][30];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_csr_cmd = {_RANDOM[10'hCE][31], _RANDOM[10'hCF][1:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_is_load = _RANDOM[10'hCF][2];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_is_sta = _RANDOM[10'hCF][3];	// lsu.scala:210:16
        ldq_12_bits_uop_ctrl_is_std = _RANDOM[10'hCF][4];	// lsu.scala:210:16
        ldq_12_bits_uop_iw_state = _RANDOM[10'hCF][6:5];	// lsu.scala:210:16
        ldq_12_bits_uop_iw_p1_poisoned = _RANDOM[10'hCF][7];	// lsu.scala:210:16
        ldq_12_bits_uop_iw_p2_poisoned = _RANDOM[10'hCF][8];	// lsu.scala:210:16
        ldq_12_bits_uop_is_br = _RANDOM[10'hCF][9];	// lsu.scala:210:16
        ldq_12_bits_uop_is_jalr = _RANDOM[10'hCF][10];	// lsu.scala:210:16
        ldq_12_bits_uop_is_jal = _RANDOM[10'hCF][11];	// lsu.scala:210:16
        ldq_12_bits_uop_is_sfb = _RANDOM[10'hCF][12];	// lsu.scala:210:16
        ldq_12_bits_uop_br_mask = _RANDOM[10'hCF][24:13];	// lsu.scala:210:16
        ldq_12_bits_uop_br_tag = _RANDOM[10'hCF][28:25];	// lsu.scala:210:16
        ldq_12_bits_uop_ftq_idx = {_RANDOM[10'hCF][31:29], _RANDOM[10'hD0][1:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_edge_inst = _RANDOM[10'hD0][2];	// lsu.scala:210:16
        ldq_12_bits_uop_pc_lob = _RANDOM[10'hD0][8:3];	// lsu.scala:210:16
        ldq_12_bits_uop_taken = _RANDOM[10'hD0][9];	// lsu.scala:210:16
        ldq_12_bits_uop_imm_packed = _RANDOM[10'hD0][29:10];	// lsu.scala:210:16
        ldq_12_bits_uop_csr_addr = {_RANDOM[10'hD0][31:30], _RANDOM[10'hD1][9:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_rob_idx = _RANDOM[10'hD1][15:10];	// lsu.scala:210:16
        ldq_12_bits_uop_ldq_idx = _RANDOM[10'hD1][19:16];	// lsu.scala:210:16
        ldq_12_bits_uop_stq_idx = _RANDOM[10'hD1][23:20];	// lsu.scala:210:16
        ldq_12_bits_uop_rxq_idx = _RANDOM[10'hD1][25:24];	// lsu.scala:210:16
        ldq_12_bits_uop_pdst = {_RANDOM[10'hD1][31:26], _RANDOM[10'hD2][0]};	// lsu.scala:210:16
        ldq_12_bits_uop_prs1 = _RANDOM[10'hD2][7:1];	// lsu.scala:210:16
        ldq_12_bits_uop_prs2 = _RANDOM[10'hD2][14:8];	// lsu.scala:210:16
        ldq_12_bits_uop_prs3 = _RANDOM[10'hD2][21:15];	// lsu.scala:210:16
        ldq_12_bits_uop_ppred = _RANDOM[10'hD2][26:22];	// lsu.scala:210:16
        ldq_12_bits_uop_prs1_busy = _RANDOM[10'hD2][27];	// lsu.scala:210:16
        ldq_12_bits_uop_prs2_busy = _RANDOM[10'hD2][28];	// lsu.scala:210:16
        ldq_12_bits_uop_prs3_busy = _RANDOM[10'hD2][29];	// lsu.scala:210:16
        ldq_12_bits_uop_ppred_busy = _RANDOM[10'hD2][30];	// lsu.scala:210:16
        ldq_12_bits_uop_stale_pdst = {_RANDOM[10'hD2][31], _RANDOM[10'hD3][5:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_exception = _RANDOM[10'hD3][6];	// lsu.scala:210:16
        ldq_12_bits_uop_exc_cause =
          {_RANDOM[10'hD3][31:7], _RANDOM[10'hD4], _RANDOM[10'hD5][6:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_bypassable = _RANDOM[10'hD5][7];	// lsu.scala:210:16
        ldq_12_bits_uop_mem_cmd = _RANDOM[10'hD5][12:8];	// lsu.scala:210:16
        ldq_12_bits_uop_mem_size = _RANDOM[10'hD5][14:13];	// lsu.scala:210:16
        ldq_12_bits_uop_mem_signed = _RANDOM[10'hD5][15];	// lsu.scala:210:16
        ldq_12_bits_uop_is_fence = _RANDOM[10'hD5][16];	// lsu.scala:210:16
        ldq_12_bits_uop_is_fencei = _RANDOM[10'hD5][17];	// lsu.scala:210:16
        ldq_12_bits_uop_is_amo = _RANDOM[10'hD5][18];	// lsu.scala:210:16
        ldq_12_bits_uop_uses_ldq = _RANDOM[10'hD5][19];	// lsu.scala:210:16
        ldq_12_bits_uop_uses_stq = _RANDOM[10'hD5][20];	// lsu.scala:210:16
        ldq_12_bits_uop_is_sys_pc2epc = _RANDOM[10'hD5][21];	// lsu.scala:210:16
        ldq_12_bits_uop_is_unique = _RANDOM[10'hD5][22];	// lsu.scala:210:16
        ldq_12_bits_uop_flush_on_commit = _RANDOM[10'hD5][23];	// lsu.scala:210:16
        ldq_12_bits_uop_ldst_is_rs1 = _RANDOM[10'hD5][24];	// lsu.scala:210:16
        ldq_12_bits_uop_ldst = _RANDOM[10'hD5][30:25];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs1 = {_RANDOM[10'hD5][31], _RANDOM[10'hD6][4:0]};	// lsu.scala:210:16
        ldq_12_bits_uop_lrs2 = _RANDOM[10'hD6][10:5];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs3 = _RANDOM[10'hD6][16:11];	// lsu.scala:210:16
        ldq_12_bits_uop_ldst_val = _RANDOM[10'hD6][17];	// lsu.scala:210:16
        ldq_12_bits_uop_dst_rtype = _RANDOM[10'hD6][19:18];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs1_rtype = _RANDOM[10'hD6][21:20];	// lsu.scala:210:16
        ldq_12_bits_uop_lrs2_rtype = _RANDOM[10'hD6][23:22];	// lsu.scala:210:16
        ldq_12_bits_uop_frs3_en = _RANDOM[10'hD6][24];	// lsu.scala:210:16
        ldq_12_bits_uop_fp_val = _RANDOM[10'hD6][25];	// lsu.scala:210:16
        ldq_12_bits_uop_fp_single = _RANDOM[10'hD6][26];	// lsu.scala:210:16
        ldq_12_bits_uop_xcpt_pf_if = _RANDOM[10'hD6][27];	// lsu.scala:210:16
        ldq_12_bits_uop_xcpt_ae_if = _RANDOM[10'hD6][28];	// lsu.scala:210:16
        ldq_12_bits_uop_xcpt_ma_if = _RANDOM[10'hD6][29];	// lsu.scala:210:16
        ldq_12_bits_uop_bp_debug_if = _RANDOM[10'hD6][30];	// lsu.scala:210:16
        ldq_12_bits_uop_bp_xcpt_if = _RANDOM[10'hD6][31];	// lsu.scala:210:16
        ldq_12_bits_uop_debug_fsrc = _RANDOM[10'hD7][1:0];	// lsu.scala:210:16
        ldq_12_bits_uop_debug_tsrc = _RANDOM[10'hD7][3:2];	// lsu.scala:210:16
        ldq_12_bits_addr_valid = _RANDOM[10'hD7][4];	// lsu.scala:210:16
        ldq_12_bits_addr_bits = {_RANDOM[10'hD7][31:5], _RANDOM[10'hD8][12:0]};	// lsu.scala:210:16
        ldq_12_bits_addr_is_virtual = _RANDOM[10'hD8][13];	// lsu.scala:210:16
        ldq_12_bits_addr_is_uncacheable = _RANDOM[10'hD8][14];	// lsu.scala:210:16
        ldq_12_bits_executed = _RANDOM[10'hD8][15];	// lsu.scala:210:16
        ldq_12_bits_succeeded = _RANDOM[10'hD8][16];	// lsu.scala:210:16
        ldq_12_bits_order_fail = _RANDOM[10'hD8][17];	// lsu.scala:210:16
        ldq_12_bits_observed = _RANDOM[10'hD8][18];	// lsu.scala:210:16
        ldq_12_bits_st_dep_mask = {_RANDOM[10'hD8][31:19], _RANDOM[10'hD9][2:0]};	// lsu.scala:210:16
        ldq_12_bits_youngest_stq_idx = _RANDOM[10'hD9][6:3];	// lsu.scala:210:16
        ldq_12_bits_forward_std_val = _RANDOM[10'hD9][7];	// lsu.scala:210:16
        ldq_12_bits_forward_stq_idx = _RANDOM[10'hD9][11:8];	// lsu.scala:210:16
        ldq_13_valid = _RANDOM[10'hDB][12];	// lsu.scala:210:16
        ldq_13_bits_uop_uopc = _RANDOM[10'hDB][19:13];	// lsu.scala:210:16
        ldq_13_bits_uop_inst = {_RANDOM[10'hDB][31:20], _RANDOM[10'hDC][19:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_debug_inst = {_RANDOM[10'hDC][31:20], _RANDOM[10'hDD][19:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_is_rvc = _RANDOM[10'hDD][20];	// lsu.scala:210:16
        ldq_13_bits_uop_debug_pc = {_RANDOM[10'hDD][31:21], _RANDOM[10'hDE][28:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_iq_type = _RANDOM[10'hDE][31:29];	// lsu.scala:210:16
        ldq_13_bits_uop_fu_code = _RANDOM[10'hDF][9:0];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_br_type = _RANDOM[10'hDF][13:10];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_op1_sel = _RANDOM[10'hDF][15:14];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_op2_sel = _RANDOM[10'hDF][18:16];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_imm_sel = _RANDOM[10'hDF][21:19];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_op_fcn = _RANDOM[10'hDF][25:22];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_fcn_dw = _RANDOM[10'hDF][26];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_csr_cmd = _RANDOM[10'hDF][29:27];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_is_load = _RANDOM[10'hDF][30];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_is_sta = _RANDOM[10'hDF][31];	// lsu.scala:210:16
        ldq_13_bits_uop_ctrl_is_std = _RANDOM[10'hE0][0];	// lsu.scala:210:16
        ldq_13_bits_uop_iw_state = _RANDOM[10'hE0][2:1];	// lsu.scala:210:16
        ldq_13_bits_uop_iw_p1_poisoned = _RANDOM[10'hE0][3];	// lsu.scala:210:16
        ldq_13_bits_uop_iw_p2_poisoned = _RANDOM[10'hE0][4];	// lsu.scala:210:16
        ldq_13_bits_uop_is_br = _RANDOM[10'hE0][5];	// lsu.scala:210:16
        ldq_13_bits_uop_is_jalr = _RANDOM[10'hE0][6];	// lsu.scala:210:16
        ldq_13_bits_uop_is_jal = _RANDOM[10'hE0][7];	// lsu.scala:210:16
        ldq_13_bits_uop_is_sfb = _RANDOM[10'hE0][8];	// lsu.scala:210:16
        ldq_13_bits_uop_br_mask = _RANDOM[10'hE0][20:9];	// lsu.scala:210:16
        ldq_13_bits_uop_br_tag = _RANDOM[10'hE0][24:21];	// lsu.scala:210:16
        ldq_13_bits_uop_ftq_idx = _RANDOM[10'hE0][29:25];	// lsu.scala:210:16
        ldq_13_bits_uop_edge_inst = _RANDOM[10'hE0][30];	// lsu.scala:210:16
        ldq_13_bits_uop_pc_lob = {_RANDOM[10'hE0][31], _RANDOM[10'hE1][4:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_taken = _RANDOM[10'hE1][5];	// lsu.scala:210:16
        ldq_13_bits_uop_imm_packed = _RANDOM[10'hE1][25:6];	// lsu.scala:210:16
        ldq_13_bits_uop_csr_addr = {_RANDOM[10'hE1][31:26], _RANDOM[10'hE2][5:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_rob_idx = _RANDOM[10'hE2][11:6];	// lsu.scala:210:16
        ldq_13_bits_uop_ldq_idx = _RANDOM[10'hE2][15:12];	// lsu.scala:210:16
        ldq_13_bits_uop_stq_idx = _RANDOM[10'hE2][19:16];	// lsu.scala:210:16
        ldq_13_bits_uop_rxq_idx = _RANDOM[10'hE2][21:20];	// lsu.scala:210:16
        ldq_13_bits_uop_pdst = _RANDOM[10'hE2][28:22];	// lsu.scala:210:16
        ldq_13_bits_uop_prs1 = {_RANDOM[10'hE2][31:29], _RANDOM[10'hE3][3:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_prs2 = _RANDOM[10'hE3][10:4];	// lsu.scala:210:16
        ldq_13_bits_uop_prs3 = _RANDOM[10'hE3][17:11];	// lsu.scala:210:16
        ldq_13_bits_uop_ppred = _RANDOM[10'hE3][22:18];	// lsu.scala:210:16
        ldq_13_bits_uop_prs1_busy = _RANDOM[10'hE3][23];	// lsu.scala:210:16
        ldq_13_bits_uop_prs2_busy = _RANDOM[10'hE3][24];	// lsu.scala:210:16
        ldq_13_bits_uop_prs3_busy = _RANDOM[10'hE3][25];	// lsu.scala:210:16
        ldq_13_bits_uop_ppred_busy = _RANDOM[10'hE3][26];	// lsu.scala:210:16
        ldq_13_bits_uop_stale_pdst = {_RANDOM[10'hE3][31:27], _RANDOM[10'hE4][1:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_exception = _RANDOM[10'hE4][2];	// lsu.scala:210:16
        ldq_13_bits_uop_exc_cause =
          {_RANDOM[10'hE4][31:3], _RANDOM[10'hE5], _RANDOM[10'hE6][2:0]};	// lsu.scala:210:16
        ldq_13_bits_uop_bypassable = _RANDOM[10'hE6][3];	// lsu.scala:210:16
        ldq_13_bits_uop_mem_cmd = _RANDOM[10'hE6][8:4];	// lsu.scala:210:16
        ldq_13_bits_uop_mem_size = _RANDOM[10'hE6][10:9];	// lsu.scala:210:16
        ldq_13_bits_uop_mem_signed = _RANDOM[10'hE6][11];	// lsu.scala:210:16
        ldq_13_bits_uop_is_fence = _RANDOM[10'hE6][12];	// lsu.scala:210:16
        ldq_13_bits_uop_is_fencei = _RANDOM[10'hE6][13];	// lsu.scala:210:16
        ldq_13_bits_uop_is_amo = _RANDOM[10'hE6][14];	// lsu.scala:210:16
        ldq_13_bits_uop_uses_ldq = _RANDOM[10'hE6][15];	// lsu.scala:210:16
        ldq_13_bits_uop_uses_stq = _RANDOM[10'hE6][16];	// lsu.scala:210:16
        ldq_13_bits_uop_is_sys_pc2epc = _RANDOM[10'hE6][17];	// lsu.scala:210:16
        ldq_13_bits_uop_is_unique = _RANDOM[10'hE6][18];	// lsu.scala:210:16
        ldq_13_bits_uop_flush_on_commit = _RANDOM[10'hE6][19];	// lsu.scala:210:16
        ldq_13_bits_uop_ldst_is_rs1 = _RANDOM[10'hE6][20];	// lsu.scala:210:16
        ldq_13_bits_uop_ldst = _RANDOM[10'hE6][26:21];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs1 = {_RANDOM[10'hE6][31:27], _RANDOM[10'hE7][0]};	// lsu.scala:210:16
        ldq_13_bits_uop_lrs2 = _RANDOM[10'hE7][6:1];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs3 = _RANDOM[10'hE7][12:7];	// lsu.scala:210:16
        ldq_13_bits_uop_ldst_val = _RANDOM[10'hE7][13];	// lsu.scala:210:16
        ldq_13_bits_uop_dst_rtype = _RANDOM[10'hE7][15:14];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs1_rtype = _RANDOM[10'hE7][17:16];	// lsu.scala:210:16
        ldq_13_bits_uop_lrs2_rtype = _RANDOM[10'hE7][19:18];	// lsu.scala:210:16
        ldq_13_bits_uop_frs3_en = _RANDOM[10'hE7][20];	// lsu.scala:210:16
        ldq_13_bits_uop_fp_val = _RANDOM[10'hE7][21];	// lsu.scala:210:16
        ldq_13_bits_uop_fp_single = _RANDOM[10'hE7][22];	// lsu.scala:210:16
        ldq_13_bits_uop_xcpt_pf_if = _RANDOM[10'hE7][23];	// lsu.scala:210:16
        ldq_13_bits_uop_xcpt_ae_if = _RANDOM[10'hE7][24];	// lsu.scala:210:16
        ldq_13_bits_uop_xcpt_ma_if = _RANDOM[10'hE7][25];	// lsu.scala:210:16
        ldq_13_bits_uop_bp_debug_if = _RANDOM[10'hE7][26];	// lsu.scala:210:16
        ldq_13_bits_uop_bp_xcpt_if = _RANDOM[10'hE7][27];	// lsu.scala:210:16
        ldq_13_bits_uop_debug_fsrc = _RANDOM[10'hE7][29:28];	// lsu.scala:210:16
        ldq_13_bits_uop_debug_tsrc = _RANDOM[10'hE7][31:30];	// lsu.scala:210:16
        ldq_13_bits_addr_valid = _RANDOM[10'hE8][0];	// lsu.scala:210:16
        ldq_13_bits_addr_bits = {_RANDOM[10'hE8][31:1], _RANDOM[10'hE9][8:0]};	// lsu.scala:210:16
        ldq_13_bits_addr_is_virtual = _RANDOM[10'hE9][9];	// lsu.scala:210:16
        ldq_13_bits_addr_is_uncacheable = _RANDOM[10'hE9][10];	// lsu.scala:210:16
        ldq_13_bits_executed = _RANDOM[10'hE9][11];	// lsu.scala:210:16
        ldq_13_bits_succeeded = _RANDOM[10'hE9][12];	// lsu.scala:210:16
        ldq_13_bits_order_fail = _RANDOM[10'hE9][13];	// lsu.scala:210:16
        ldq_13_bits_observed = _RANDOM[10'hE9][14];	// lsu.scala:210:16
        ldq_13_bits_st_dep_mask = _RANDOM[10'hE9][30:15];	// lsu.scala:210:16
        ldq_13_bits_youngest_stq_idx = {_RANDOM[10'hE9][31], _RANDOM[10'hEA][2:0]};	// lsu.scala:210:16
        ldq_13_bits_forward_std_val = _RANDOM[10'hEA][3];	// lsu.scala:210:16
        ldq_13_bits_forward_stq_idx = _RANDOM[10'hEA][7:4];	// lsu.scala:210:16
        ldq_14_valid = _RANDOM[10'hEC][8];	// lsu.scala:210:16
        ldq_14_bits_uop_uopc = _RANDOM[10'hEC][15:9];	// lsu.scala:210:16
        ldq_14_bits_uop_inst = {_RANDOM[10'hEC][31:16], _RANDOM[10'hED][15:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_debug_inst = {_RANDOM[10'hED][31:16], _RANDOM[10'hEE][15:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_is_rvc = _RANDOM[10'hEE][16];	// lsu.scala:210:16
        ldq_14_bits_uop_debug_pc = {_RANDOM[10'hEE][31:17], _RANDOM[10'hEF][24:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_iq_type = _RANDOM[10'hEF][27:25];	// lsu.scala:210:16
        ldq_14_bits_uop_fu_code = {_RANDOM[10'hEF][31:28], _RANDOM[10'hF0][5:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_br_type = _RANDOM[10'hF0][9:6];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_op1_sel = _RANDOM[10'hF0][11:10];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_op2_sel = _RANDOM[10'hF0][14:12];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_imm_sel = _RANDOM[10'hF0][17:15];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_op_fcn = _RANDOM[10'hF0][21:18];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_fcn_dw = _RANDOM[10'hF0][22];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_csr_cmd = _RANDOM[10'hF0][25:23];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_is_load = _RANDOM[10'hF0][26];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_is_sta = _RANDOM[10'hF0][27];	// lsu.scala:210:16
        ldq_14_bits_uop_ctrl_is_std = _RANDOM[10'hF0][28];	// lsu.scala:210:16
        ldq_14_bits_uop_iw_state = _RANDOM[10'hF0][30:29];	// lsu.scala:210:16
        ldq_14_bits_uop_iw_p1_poisoned = _RANDOM[10'hF0][31];	// lsu.scala:210:16
        ldq_14_bits_uop_iw_p2_poisoned = _RANDOM[10'hF1][0];	// lsu.scala:210:16
        ldq_14_bits_uop_is_br = _RANDOM[10'hF1][1];	// lsu.scala:210:16
        ldq_14_bits_uop_is_jalr = _RANDOM[10'hF1][2];	// lsu.scala:210:16
        ldq_14_bits_uop_is_jal = _RANDOM[10'hF1][3];	// lsu.scala:210:16
        ldq_14_bits_uop_is_sfb = _RANDOM[10'hF1][4];	// lsu.scala:210:16
        ldq_14_bits_uop_br_mask = _RANDOM[10'hF1][16:5];	// lsu.scala:210:16
        ldq_14_bits_uop_br_tag = _RANDOM[10'hF1][20:17];	// lsu.scala:210:16
        ldq_14_bits_uop_ftq_idx = _RANDOM[10'hF1][25:21];	// lsu.scala:210:16
        ldq_14_bits_uop_edge_inst = _RANDOM[10'hF1][26];	// lsu.scala:210:16
        ldq_14_bits_uop_pc_lob = {_RANDOM[10'hF1][31:27], _RANDOM[10'hF2][0]};	// lsu.scala:210:16
        ldq_14_bits_uop_taken = _RANDOM[10'hF2][1];	// lsu.scala:210:16
        ldq_14_bits_uop_imm_packed = _RANDOM[10'hF2][21:2];	// lsu.scala:210:16
        ldq_14_bits_uop_csr_addr = {_RANDOM[10'hF2][31:22], _RANDOM[10'hF3][1:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_rob_idx = _RANDOM[10'hF3][7:2];	// lsu.scala:210:16
        ldq_14_bits_uop_ldq_idx = _RANDOM[10'hF3][11:8];	// lsu.scala:210:16
        ldq_14_bits_uop_stq_idx = _RANDOM[10'hF3][15:12];	// lsu.scala:210:16
        ldq_14_bits_uop_rxq_idx = _RANDOM[10'hF3][17:16];	// lsu.scala:210:16
        ldq_14_bits_uop_pdst = _RANDOM[10'hF3][24:18];	// lsu.scala:210:16
        ldq_14_bits_uop_prs1 = _RANDOM[10'hF3][31:25];	// lsu.scala:210:16
        ldq_14_bits_uop_prs2 = _RANDOM[10'hF4][6:0];	// lsu.scala:210:16
        ldq_14_bits_uop_prs3 = _RANDOM[10'hF4][13:7];	// lsu.scala:210:16
        ldq_14_bits_uop_ppred = _RANDOM[10'hF4][18:14];	// lsu.scala:210:16
        ldq_14_bits_uop_prs1_busy = _RANDOM[10'hF4][19];	// lsu.scala:210:16
        ldq_14_bits_uop_prs2_busy = _RANDOM[10'hF4][20];	// lsu.scala:210:16
        ldq_14_bits_uop_prs3_busy = _RANDOM[10'hF4][21];	// lsu.scala:210:16
        ldq_14_bits_uop_ppred_busy = _RANDOM[10'hF4][22];	// lsu.scala:210:16
        ldq_14_bits_uop_stale_pdst = _RANDOM[10'hF4][29:23];	// lsu.scala:210:16
        ldq_14_bits_uop_exception = _RANDOM[10'hF4][30];	// lsu.scala:210:16
        ldq_14_bits_uop_exc_cause =
          {_RANDOM[10'hF4][31], _RANDOM[10'hF5], _RANDOM[10'hF6][30:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_bypassable = _RANDOM[10'hF6][31];	// lsu.scala:210:16
        ldq_14_bits_uop_mem_cmd = _RANDOM[10'hF7][4:0];	// lsu.scala:210:16
        ldq_14_bits_uop_mem_size = _RANDOM[10'hF7][6:5];	// lsu.scala:210:16
        ldq_14_bits_uop_mem_signed = _RANDOM[10'hF7][7];	// lsu.scala:210:16
        ldq_14_bits_uop_is_fence = _RANDOM[10'hF7][8];	// lsu.scala:210:16
        ldq_14_bits_uop_is_fencei = _RANDOM[10'hF7][9];	// lsu.scala:210:16
        ldq_14_bits_uop_is_amo = _RANDOM[10'hF7][10];	// lsu.scala:210:16
        ldq_14_bits_uop_uses_ldq = _RANDOM[10'hF7][11];	// lsu.scala:210:16
        ldq_14_bits_uop_uses_stq = _RANDOM[10'hF7][12];	// lsu.scala:210:16
        ldq_14_bits_uop_is_sys_pc2epc = _RANDOM[10'hF7][13];	// lsu.scala:210:16
        ldq_14_bits_uop_is_unique = _RANDOM[10'hF7][14];	// lsu.scala:210:16
        ldq_14_bits_uop_flush_on_commit = _RANDOM[10'hF7][15];	// lsu.scala:210:16
        ldq_14_bits_uop_ldst_is_rs1 = _RANDOM[10'hF7][16];	// lsu.scala:210:16
        ldq_14_bits_uop_ldst = _RANDOM[10'hF7][22:17];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs1 = _RANDOM[10'hF7][28:23];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs2 = {_RANDOM[10'hF7][31:29], _RANDOM[10'hF8][2:0]};	// lsu.scala:210:16
        ldq_14_bits_uop_lrs3 = _RANDOM[10'hF8][8:3];	// lsu.scala:210:16
        ldq_14_bits_uop_ldst_val = _RANDOM[10'hF8][9];	// lsu.scala:210:16
        ldq_14_bits_uop_dst_rtype = _RANDOM[10'hF8][11:10];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs1_rtype = _RANDOM[10'hF8][13:12];	// lsu.scala:210:16
        ldq_14_bits_uop_lrs2_rtype = _RANDOM[10'hF8][15:14];	// lsu.scala:210:16
        ldq_14_bits_uop_frs3_en = _RANDOM[10'hF8][16];	// lsu.scala:210:16
        ldq_14_bits_uop_fp_val = _RANDOM[10'hF8][17];	// lsu.scala:210:16
        ldq_14_bits_uop_fp_single = _RANDOM[10'hF8][18];	// lsu.scala:210:16
        ldq_14_bits_uop_xcpt_pf_if = _RANDOM[10'hF8][19];	// lsu.scala:210:16
        ldq_14_bits_uop_xcpt_ae_if = _RANDOM[10'hF8][20];	// lsu.scala:210:16
        ldq_14_bits_uop_xcpt_ma_if = _RANDOM[10'hF8][21];	// lsu.scala:210:16
        ldq_14_bits_uop_bp_debug_if = _RANDOM[10'hF8][22];	// lsu.scala:210:16
        ldq_14_bits_uop_bp_xcpt_if = _RANDOM[10'hF8][23];	// lsu.scala:210:16
        ldq_14_bits_uop_debug_fsrc = _RANDOM[10'hF8][25:24];	// lsu.scala:210:16
        ldq_14_bits_uop_debug_tsrc = _RANDOM[10'hF8][27:26];	// lsu.scala:210:16
        ldq_14_bits_addr_valid = _RANDOM[10'hF8][28];	// lsu.scala:210:16
        ldq_14_bits_addr_bits =
          {_RANDOM[10'hF8][31:29], _RANDOM[10'hF9], _RANDOM[10'hFA][4:0]};	// lsu.scala:210:16
        ldq_14_bits_addr_is_virtual = _RANDOM[10'hFA][5];	// lsu.scala:210:16
        ldq_14_bits_addr_is_uncacheable = _RANDOM[10'hFA][6];	// lsu.scala:210:16
        ldq_14_bits_executed = _RANDOM[10'hFA][7];	// lsu.scala:210:16
        ldq_14_bits_succeeded = _RANDOM[10'hFA][8];	// lsu.scala:210:16
        ldq_14_bits_order_fail = _RANDOM[10'hFA][9];	// lsu.scala:210:16
        ldq_14_bits_observed = _RANDOM[10'hFA][10];	// lsu.scala:210:16
        ldq_14_bits_st_dep_mask = _RANDOM[10'hFA][26:11];	// lsu.scala:210:16
        ldq_14_bits_youngest_stq_idx = _RANDOM[10'hFA][30:27];	// lsu.scala:210:16
        ldq_14_bits_forward_std_val = _RANDOM[10'hFA][31];	// lsu.scala:210:16
        ldq_14_bits_forward_stq_idx = _RANDOM[10'hFB][3:0];	// lsu.scala:210:16
        ldq_15_valid = _RANDOM[10'hFD][4];	// lsu.scala:210:16
        ldq_15_bits_uop_uopc = _RANDOM[10'hFD][11:5];	// lsu.scala:210:16
        ldq_15_bits_uop_inst = {_RANDOM[10'hFD][31:12], _RANDOM[10'hFE][11:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_debug_inst = {_RANDOM[10'hFE][31:12], _RANDOM[10'hFF][11:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_is_rvc = _RANDOM[10'hFF][12];	// lsu.scala:210:16
        ldq_15_bits_uop_debug_pc = {_RANDOM[10'hFF][31:13], _RANDOM[10'h100][20:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_iq_type = _RANDOM[10'h100][23:21];	// lsu.scala:210:16
        ldq_15_bits_uop_fu_code = {_RANDOM[10'h100][31:24], _RANDOM[10'h101][1:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_br_type = _RANDOM[10'h101][5:2];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_op1_sel = _RANDOM[10'h101][7:6];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_op2_sel = _RANDOM[10'h101][10:8];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_imm_sel = _RANDOM[10'h101][13:11];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_op_fcn = _RANDOM[10'h101][17:14];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_fcn_dw = _RANDOM[10'h101][18];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_csr_cmd = _RANDOM[10'h101][21:19];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_is_load = _RANDOM[10'h101][22];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_is_sta = _RANDOM[10'h101][23];	// lsu.scala:210:16
        ldq_15_bits_uop_ctrl_is_std = _RANDOM[10'h101][24];	// lsu.scala:210:16
        ldq_15_bits_uop_iw_state = _RANDOM[10'h101][26:25];	// lsu.scala:210:16
        ldq_15_bits_uop_iw_p1_poisoned = _RANDOM[10'h101][27];	// lsu.scala:210:16
        ldq_15_bits_uop_iw_p2_poisoned = _RANDOM[10'h101][28];	// lsu.scala:210:16
        ldq_15_bits_uop_is_br = _RANDOM[10'h101][29];	// lsu.scala:210:16
        ldq_15_bits_uop_is_jalr = _RANDOM[10'h101][30];	// lsu.scala:210:16
        ldq_15_bits_uop_is_jal = _RANDOM[10'h101][31];	// lsu.scala:210:16
        ldq_15_bits_uop_is_sfb = _RANDOM[10'h102][0];	// lsu.scala:210:16
        ldq_15_bits_uop_br_mask = _RANDOM[10'h102][12:1];	// lsu.scala:210:16
        ldq_15_bits_uop_br_tag = _RANDOM[10'h102][16:13];	// lsu.scala:210:16
        ldq_15_bits_uop_ftq_idx = _RANDOM[10'h102][21:17];	// lsu.scala:210:16
        ldq_15_bits_uop_edge_inst = _RANDOM[10'h102][22];	// lsu.scala:210:16
        ldq_15_bits_uop_pc_lob = _RANDOM[10'h102][28:23];	// lsu.scala:210:16
        ldq_15_bits_uop_taken = _RANDOM[10'h102][29];	// lsu.scala:210:16
        ldq_15_bits_uop_imm_packed = {_RANDOM[10'h102][31:30], _RANDOM[10'h103][17:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_csr_addr = _RANDOM[10'h103][29:18];	// lsu.scala:210:16
        ldq_15_bits_uop_rob_idx = {_RANDOM[10'h103][31:30], _RANDOM[10'h104][3:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_ldq_idx = _RANDOM[10'h104][7:4];	// lsu.scala:210:16
        ldq_15_bits_uop_stq_idx = _RANDOM[10'h104][11:8];	// lsu.scala:210:16
        ldq_15_bits_uop_rxq_idx = _RANDOM[10'h104][13:12];	// lsu.scala:210:16
        ldq_15_bits_uop_pdst = _RANDOM[10'h104][20:14];	// lsu.scala:210:16
        ldq_15_bits_uop_prs1 = _RANDOM[10'h104][27:21];	// lsu.scala:210:16
        ldq_15_bits_uop_prs2 = {_RANDOM[10'h104][31:28], _RANDOM[10'h105][2:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_prs3 = _RANDOM[10'h105][9:3];	// lsu.scala:210:16
        ldq_15_bits_uop_ppred = _RANDOM[10'h105][14:10];	// lsu.scala:210:16
        ldq_15_bits_uop_prs1_busy = _RANDOM[10'h105][15];	// lsu.scala:210:16
        ldq_15_bits_uop_prs2_busy = _RANDOM[10'h105][16];	// lsu.scala:210:16
        ldq_15_bits_uop_prs3_busy = _RANDOM[10'h105][17];	// lsu.scala:210:16
        ldq_15_bits_uop_ppred_busy = _RANDOM[10'h105][18];	// lsu.scala:210:16
        ldq_15_bits_uop_stale_pdst = _RANDOM[10'h105][25:19];	// lsu.scala:210:16
        ldq_15_bits_uop_exception = _RANDOM[10'h105][26];	// lsu.scala:210:16
        ldq_15_bits_uop_exc_cause =
          {_RANDOM[10'h105][31:27], _RANDOM[10'h106], _RANDOM[10'h107][26:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_bypassable = _RANDOM[10'h107][27];	// lsu.scala:210:16
        ldq_15_bits_uop_mem_cmd = {_RANDOM[10'h107][31:28], _RANDOM[10'h108][0]};	// lsu.scala:210:16
        ldq_15_bits_uop_mem_size = _RANDOM[10'h108][2:1];	// lsu.scala:210:16
        ldq_15_bits_uop_mem_signed = _RANDOM[10'h108][3];	// lsu.scala:210:16
        ldq_15_bits_uop_is_fence = _RANDOM[10'h108][4];	// lsu.scala:210:16
        ldq_15_bits_uop_is_fencei = _RANDOM[10'h108][5];	// lsu.scala:210:16
        ldq_15_bits_uop_is_amo = _RANDOM[10'h108][6];	// lsu.scala:210:16
        ldq_15_bits_uop_uses_ldq = _RANDOM[10'h108][7];	// lsu.scala:210:16
        ldq_15_bits_uop_uses_stq = _RANDOM[10'h108][8];	// lsu.scala:210:16
        ldq_15_bits_uop_is_sys_pc2epc = _RANDOM[10'h108][9];	// lsu.scala:210:16
        ldq_15_bits_uop_is_unique = _RANDOM[10'h108][10];	// lsu.scala:210:16
        ldq_15_bits_uop_flush_on_commit = _RANDOM[10'h108][11];	// lsu.scala:210:16
        ldq_15_bits_uop_ldst_is_rs1 = _RANDOM[10'h108][12];	// lsu.scala:210:16
        ldq_15_bits_uop_ldst = _RANDOM[10'h108][18:13];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs1 = _RANDOM[10'h108][24:19];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs2 = _RANDOM[10'h108][30:25];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs3 = {_RANDOM[10'h108][31], _RANDOM[10'h109][4:0]};	// lsu.scala:210:16
        ldq_15_bits_uop_ldst_val = _RANDOM[10'h109][5];	// lsu.scala:210:16
        ldq_15_bits_uop_dst_rtype = _RANDOM[10'h109][7:6];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs1_rtype = _RANDOM[10'h109][9:8];	// lsu.scala:210:16
        ldq_15_bits_uop_lrs2_rtype = _RANDOM[10'h109][11:10];	// lsu.scala:210:16
        ldq_15_bits_uop_frs3_en = _RANDOM[10'h109][12];	// lsu.scala:210:16
        ldq_15_bits_uop_fp_val = _RANDOM[10'h109][13];	// lsu.scala:210:16
        ldq_15_bits_uop_fp_single = _RANDOM[10'h109][14];	// lsu.scala:210:16
        ldq_15_bits_uop_xcpt_pf_if = _RANDOM[10'h109][15];	// lsu.scala:210:16
        ldq_15_bits_uop_xcpt_ae_if = _RANDOM[10'h109][16];	// lsu.scala:210:16
        ldq_15_bits_uop_xcpt_ma_if = _RANDOM[10'h109][17];	// lsu.scala:210:16
        ldq_15_bits_uop_bp_debug_if = _RANDOM[10'h109][18];	// lsu.scala:210:16
        ldq_15_bits_uop_bp_xcpt_if = _RANDOM[10'h109][19];	// lsu.scala:210:16
        ldq_15_bits_uop_debug_fsrc = _RANDOM[10'h109][21:20];	// lsu.scala:210:16
        ldq_15_bits_uop_debug_tsrc = _RANDOM[10'h109][23:22];	// lsu.scala:210:16
        ldq_15_bits_addr_valid = _RANDOM[10'h109][24];	// lsu.scala:210:16
        ldq_15_bits_addr_bits =
          {_RANDOM[10'h109][31:25], _RANDOM[10'h10A], _RANDOM[10'h10B][0]};	// lsu.scala:210:16
        ldq_15_bits_addr_is_virtual = _RANDOM[10'h10B][1];	// lsu.scala:210:16
        ldq_15_bits_addr_is_uncacheable = _RANDOM[10'h10B][2];	// lsu.scala:210:16
        ldq_15_bits_executed = _RANDOM[10'h10B][3];	// lsu.scala:210:16
        ldq_15_bits_succeeded = _RANDOM[10'h10B][4];	// lsu.scala:210:16
        ldq_15_bits_order_fail = _RANDOM[10'h10B][5];	// lsu.scala:210:16
        ldq_15_bits_observed = _RANDOM[10'h10B][6];	// lsu.scala:210:16
        ldq_15_bits_st_dep_mask = _RANDOM[10'h10B][22:7];	// lsu.scala:210:16
        ldq_15_bits_youngest_stq_idx = _RANDOM[10'h10B][26:23];	// lsu.scala:210:16
        ldq_15_bits_forward_std_val = _RANDOM[10'h10B][27];	// lsu.scala:210:16
        ldq_15_bits_forward_stq_idx = _RANDOM[10'h10B][31:28];	// lsu.scala:210:16
        stq_0_valid = _RANDOM[10'h10E][0];	// lsu.scala:211:16
        stq_0_bits_uop_uopc = _RANDOM[10'h10E][7:1];	// lsu.scala:211:16
        stq_0_bits_uop_inst = {_RANDOM[10'h10E][31:8], _RANDOM[10'h10F][7:0]};	// lsu.scala:211:16
        stq_0_bits_uop_debug_inst = {_RANDOM[10'h10F][31:8], _RANDOM[10'h110][7:0]};	// lsu.scala:211:16
        stq_0_bits_uop_is_rvc = _RANDOM[10'h110][8];	// lsu.scala:211:16
        stq_0_bits_uop_debug_pc = {_RANDOM[10'h110][31:9], _RANDOM[10'h111][16:0]};	// lsu.scala:211:16
        stq_0_bits_uop_iq_type = _RANDOM[10'h111][19:17];	// lsu.scala:211:16
        stq_0_bits_uop_fu_code = _RANDOM[10'h111][29:20];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_br_type = {_RANDOM[10'h111][31:30], _RANDOM[10'h112][1:0]};	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op1_sel = _RANDOM[10'h112][3:2];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op2_sel = _RANDOM[10'h112][6:4];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_imm_sel = _RANDOM[10'h112][9:7];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_op_fcn = _RANDOM[10'h112][13:10];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_fcn_dw = _RANDOM[10'h112][14];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_csr_cmd = _RANDOM[10'h112][17:15];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_is_load = _RANDOM[10'h112][18];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_is_sta = _RANDOM[10'h112][19];	// lsu.scala:211:16
        stq_0_bits_uop_ctrl_is_std = _RANDOM[10'h112][20];	// lsu.scala:211:16
        stq_0_bits_uop_iw_state = _RANDOM[10'h112][22:21];	// lsu.scala:211:16
        stq_0_bits_uop_iw_p1_poisoned = _RANDOM[10'h112][23];	// lsu.scala:211:16
        stq_0_bits_uop_iw_p2_poisoned = _RANDOM[10'h112][24];	// lsu.scala:211:16
        stq_0_bits_uop_is_br = _RANDOM[10'h112][25];	// lsu.scala:211:16
        stq_0_bits_uop_is_jalr = _RANDOM[10'h112][26];	// lsu.scala:211:16
        stq_0_bits_uop_is_jal = _RANDOM[10'h112][27];	// lsu.scala:211:16
        stq_0_bits_uop_is_sfb = _RANDOM[10'h112][28];	// lsu.scala:211:16
        stq_0_bits_uop_br_mask = {_RANDOM[10'h112][31:29], _RANDOM[10'h113][8:0]};	// lsu.scala:211:16
        stq_0_bits_uop_br_tag = _RANDOM[10'h113][12:9];	// lsu.scala:211:16
        stq_0_bits_uop_ftq_idx = _RANDOM[10'h113][17:13];	// lsu.scala:211:16
        stq_0_bits_uop_edge_inst = _RANDOM[10'h113][18];	// lsu.scala:211:16
        stq_0_bits_uop_pc_lob = _RANDOM[10'h113][24:19];	// lsu.scala:211:16
        stq_0_bits_uop_taken = _RANDOM[10'h113][25];	// lsu.scala:211:16
        stq_0_bits_uop_imm_packed = {_RANDOM[10'h113][31:26], _RANDOM[10'h114][13:0]};	// lsu.scala:211:16
        stq_0_bits_uop_csr_addr = _RANDOM[10'h114][25:14];	// lsu.scala:211:16
        stq_0_bits_uop_rob_idx = _RANDOM[10'h114][31:26];	// lsu.scala:211:16
        stq_0_bits_uop_ldq_idx = _RANDOM[10'h115][3:0];	// lsu.scala:211:16
        stq_0_bits_uop_stq_idx = _RANDOM[10'h115][7:4];	// lsu.scala:211:16
        stq_0_bits_uop_rxq_idx = _RANDOM[10'h115][9:8];	// lsu.scala:211:16
        stq_0_bits_uop_pdst = _RANDOM[10'h115][16:10];	// lsu.scala:211:16
        stq_0_bits_uop_prs1 = _RANDOM[10'h115][23:17];	// lsu.scala:211:16
        stq_0_bits_uop_prs2 = _RANDOM[10'h115][30:24];	// lsu.scala:211:16
        stq_0_bits_uop_prs3 = {_RANDOM[10'h115][31], _RANDOM[10'h116][5:0]};	// lsu.scala:211:16
        stq_0_bits_uop_ppred = _RANDOM[10'h116][10:6];	// lsu.scala:211:16
        stq_0_bits_uop_prs1_busy = _RANDOM[10'h116][11];	// lsu.scala:211:16
        stq_0_bits_uop_prs2_busy = _RANDOM[10'h116][12];	// lsu.scala:211:16
        stq_0_bits_uop_prs3_busy = _RANDOM[10'h116][13];	// lsu.scala:211:16
        stq_0_bits_uop_ppred_busy = _RANDOM[10'h116][14];	// lsu.scala:211:16
        stq_0_bits_uop_stale_pdst = _RANDOM[10'h116][21:15];	// lsu.scala:211:16
        stq_0_bits_uop_exception = _RANDOM[10'h116][22];	// lsu.scala:211:16
        stq_0_bits_uop_exc_cause =
          {_RANDOM[10'h116][31:23], _RANDOM[10'h117], _RANDOM[10'h118][22:0]};	// lsu.scala:211:16
        stq_0_bits_uop_bypassable = _RANDOM[10'h118][23];	// lsu.scala:211:16
        stq_0_bits_uop_mem_cmd = _RANDOM[10'h118][28:24];	// lsu.scala:211:16
        stq_0_bits_uop_mem_size = _RANDOM[10'h118][30:29];	// lsu.scala:211:16
        stq_0_bits_uop_mem_signed = _RANDOM[10'h118][31];	// lsu.scala:211:16
        stq_0_bits_uop_is_fence = _RANDOM[10'h119][0];	// lsu.scala:211:16
        stq_0_bits_uop_is_fencei = _RANDOM[10'h119][1];	// lsu.scala:211:16
        stq_0_bits_uop_is_amo = _RANDOM[10'h119][2];	// lsu.scala:211:16
        stq_0_bits_uop_uses_ldq = _RANDOM[10'h119][3];	// lsu.scala:211:16
        stq_0_bits_uop_uses_stq = _RANDOM[10'h119][4];	// lsu.scala:211:16
        stq_0_bits_uop_is_sys_pc2epc = _RANDOM[10'h119][5];	// lsu.scala:211:16
        stq_0_bits_uop_is_unique = _RANDOM[10'h119][6];	// lsu.scala:211:16
        stq_0_bits_uop_flush_on_commit = _RANDOM[10'h119][7];	// lsu.scala:211:16
        stq_0_bits_uop_ldst_is_rs1 = _RANDOM[10'h119][8];	// lsu.scala:211:16
        stq_0_bits_uop_ldst = _RANDOM[10'h119][14:9];	// lsu.scala:211:16
        stq_0_bits_uop_lrs1 = _RANDOM[10'h119][20:15];	// lsu.scala:211:16
        stq_0_bits_uop_lrs2 = _RANDOM[10'h119][26:21];	// lsu.scala:211:16
        stq_0_bits_uop_lrs3 = {_RANDOM[10'h119][31:27], _RANDOM[10'h11A][0]};	// lsu.scala:211:16
        stq_0_bits_uop_ldst_val = _RANDOM[10'h11A][1];	// lsu.scala:211:16
        stq_0_bits_uop_dst_rtype = _RANDOM[10'h11A][3:2];	// lsu.scala:211:16
        stq_0_bits_uop_lrs1_rtype = _RANDOM[10'h11A][5:4];	// lsu.scala:211:16
        stq_0_bits_uop_lrs2_rtype = _RANDOM[10'h11A][7:6];	// lsu.scala:211:16
        stq_0_bits_uop_frs3_en = _RANDOM[10'h11A][8];	// lsu.scala:211:16
        stq_0_bits_uop_fp_val = _RANDOM[10'h11A][9];	// lsu.scala:211:16
        stq_0_bits_uop_fp_single = _RANDOM[10'h11A][10];	// lsu.scala:211:16
        stq_0_bits_uop_xcpt_pf_if = _RANDOM[10'h11A][11];	// lsu.scala:211:16
        stq_0_bits_uop_xcpt_ae_if = _RANDOM[10'h11A][12];	// lsu.scala:211:16
        stq_0_bits_uop_xcpt_ma_if = _RANDOM[10'h11A][13];	// lsu.scala:211:16
        stq_0_bits_uop_bp_debug_if = _RANDOM[10'h11A][14];	// lsu.scala:211:16
        stq_0_bits_uop_bp_xcpt_if = _RANDOM[10'h11A][15];	// lsu.scala:211:16
        stq_0_bits_uop_debug_fsrc = _RANDOM[10'h11A][17:16];	// lsu.scala:211:16
        stq_0_bits_uop_debug_tsrc = _RANDOM[10'h11A][19:18];	// lsu.scala:211:16
        stq_0_bits_addr_valid = _RANDOM[10'h11A][20];	// lsu.scala:211:16
        stq_0_bits_addr_bits = {_RANDOM[10'h11A][31:21], _RANDOM[10'h11B][28:0]};	// lsu.scala:211:16
        stq_0_bits_addr_is_virtual = _RANDOM[10'h11B][29];	// lsu.scala:211:16
        stq_0_bits_data_valid = _RANDOM[10'h11B][30];	// lsu.scala:211:16
        stq_0_bits_data_bits =
          {_RANDOM[10'h11B][31], _RANDOM[10'h11C], _RANDOM[10'h11D][30:0]};	// lsu.scala:211:16
        stq_0_bits_committed = _RANDOM[10'h11D][31];	// lsu.scala:211:16
        stq_0_bits_succeeded = _RANDOM[10'h11E][0];	// lsu.scala:211:16
        stq_1_valid = _RANDOM[10'h120][1];	// lsu.scala:211:16
        stq_1_bits_uop_uopc = _RANDOM[10'h120][8:2];	// lsu.scala:211:16
        stq_1_bits_uop_inst = {_RANDOM[10'h120][31:9], _RANDOM[10'h121][8:0]};	// lsu.scala:211:16
        stq_1_bits_uop_debug_inst = {_RANDOM[10'h121][31:9], _RANDOM[10'h122][8:0]};	// lsu.scala:211:16
        stq_1_bits_uop_is_rvc = _RANDOM[10'h122][9];	// lsu.scala:211:16
        stq_1_bits_uop_debug_pc = {_RANDOM[10'h122][31:10], _RANDOM[10'h123][17:0]};	// lsu.scala:211:16
        stq_1_bits_uop_iq_type = _RANDOM[10'h123][20:18];	// lsu.scala:211:16
        stq_1_bits_uop_fu_code = _RANDOM[10'h123][30:21];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_br_type = {_RANDOM[10'h123][31], _RANDOM[10'h124][2:0]};	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op1_sel = _RANDOM[10'h124][4:3];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op2_sel = _RANDOM[10'h124][7:5];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_imm_sel = _RANDOM[10'h124][10:8];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_op_fcn = _RANDOM[10'h124][14:11];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_fcn_dw = _RANDOM[10'h124][15];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_csr_cmd = _RANDOM[10'h124][18:16];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_is_load = _RANDOM[10'h124][19];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_is_sta = _RANDOM[10'h124][20];	// lsu.scala:211:16
        stq_1_bits_uop_ctrl_is_std = _RANDOM[10'h124][21];	// lsu.scala:211:16
        stq_1_bits_uop_iw_state = _RANDOM[10'h124][23:22];	// lsu.scala:211:16
        stq_1_bits_uop_iw_p1_poisoned = _RANDOM[10'h124][24];	// lsu.scala:211:16
        stq_1_bits_uop_iw_p2_poisoned = _RANDOM[10'h124][25];	// lsu.scala:211:16
        stq_1_bits_uop_is_br = _RANDOM[10'h124][26];	// lsu.scala:211:16
        stq_1_bits_uop_is_jalr = _RANDOM[10'h124][27];	// lsu.scala:211:16
        stq_1_bits_uop_is_jal = _RANDOM[10'h124][28];	// lsu.scala:211:16
        stq_1_bits_uop_is_sfb = _RANDOM[10'h124][29];	// lsu.scala:211:16
        stq_1_bits_uop_br_mask = {_RANDOM[10'h124][31:30], _RANDOM[10'h125][9:0]};	// lsu.scala:211:16
        stq_1_bits_uop_br_tag = _RANDOM[10'h125][13:10];	// lsu.scala:211:16
        stq_1_bits_uop_ftq_idx = _RANDOM[10'h125][18:14];	// lsu.scala:211:16
        stq_1_bits_uop_edge_inst = _RANDOM[10'h125][19];	// lsu.scala:211:16
        stq_1_bits_uop_pc_lob = _RANDOM[10'h125][25:20];	// lsu.scala:211:16
        stq_1_bits_uop_taken = _RANDOM[10'h125][26];	// lsu.scala:211:16
        stq_1_bits_uop_imm_packed = {_RANDOM[10'h125][31:27], _RANDOM[10'h126][14:0]};	// lsu.scala:211:16
        stq_1_bits_uop_csr_addr = _RANDOM[10'h126][26:15];	// lsu.scala:211:16
        stq_1_bits_uop_rob_idx = {_RANDOM[10'h126][31:27], _RANDOM[10'h127][0]};	// lsu.scala:211:16
        stq_1_bits_uop_ldq_idx = _RANDOM[10'h127][4:1];	// lsu.scala:211:16
        stq_1_bits_uop_stq_idx = _RANDOM[10'h127][8:5];	// lsu.scala:211:16
        stq_1_bits_uop_rxq_idx = _RANDOM[10'h127][10:9];	// lsu.scala:211:16
        stq_1_bits_uop_pdst = _RANDOM[10'h127][17:11];	// lsu.scala:211:16
        stq_1_bits_uop_prs1 = _RANDOM[10'h127][24:18];	// lsu.scala:211:16
        stq_1_bits_uop_prs2 = _RANDOM[10'h127][31:25];	// lsu.scala:211:16
        stq_1_bits_uop_prs3 = _RANDOM[10'h128][6:0];	// lsu.scala:211:16
        stq_1_bits_uop_ppred = _RANDOM[10'h128][11:7];	// lsu.scala:211:16
        stq_1_bits_uop_prs1_busy = _RANDOM[10'h128][12];	// lsu.scala:211:16
        stq_1_bits_uop_prs2_busy = _RANDOM[10'h128][13];	// lsu.scala:211:16
        stq_1_bits_uop_prs3_busy = _RANDOM[10'h128][14];	// lsu.scala:211:16
        stq_1_bits_uop_ppred_busy = _RANDOM[10'h128][15];	// lsu.scala:211:16
        stq_1_bits_uop_stale_pdst = _RANDOM[10'h128][22:16];	// lsu.scala:211:16
        stq_1_bits_uop_exception = _RANDOM[10'h128][23];	// lsu.scala:211:16
        stq_1_bits_uop_exc_cause =
          {_RANDOM[10'h128][31:24], _RANDOM[10'h129], _RANDOM[10'h12A][23:0]};	// lsu.scala:211:16
        stq_1_bits_uop_bypassable = _RANDOM[10'h12A][24];	// lsu.scala:211:16
        stq_1_bits_uop_mem_cmd = _RANDOM[10'h12A][29:25];	// lsu.scala:211:16
        stq_1_bits_uop_mem_size = _RANDOM[10'h12A][31:30];	// lsu.scala:211:16
        stq_1_bits_uop_mem_signed = _RANDOM[10'h12B][0];	// lsu.scala:211:16
        stq_1_bits_uop_is_fence = _RANDOM[10'h12B][1];	// lsu.scala:211:16
        stq_1_bits_uop_is_fencei = _RANDOM[10'h12B][2];	// lsu.scala:211:16
        stq_1_bits_uop_is_amo = _RANDOM[10'h12B][3];	// lsu.scala:211:16
        stq_1_bits_uop_uses_ldq = _RANDOM[10'h12B][4];	// lsu.scala:211:16
        stq_1_bits_uop_uses_stq = _RANDOM[10'h12B][5];	// lsu.scala:211:16
        stq_1_bits_uop_is_sys_pc2epc = _RANDOM[10'h12B][6];	// lsu.scala:211:16
        stq_1_bits_uop_is_unique = _RANDOM[10'h12B][7];	// lsu.scala:211:16
        stq_1_bits_uop_flush_on_commit = _RANDOM[10'h12B][8];	// lsu.scala:211:16
        stq_1_bits_uop_ldst_is_rs1 = _RANDOM[10'h12B][9];	// lsu.scala:211:16
        stq_1_bits_uop_ldst = _RANDOM[10'h12B][15:10];	// lsu.scala:211:16
        stq_1_bits_uop_lrs1 = _RANDOM[10'h12B][21:16];	// lsu.scala:211:16
        stq_1_bits_uop_lrs2 = _RANDOM[10'h12B][27:22];	// lsu.scala:211:16
        stq_1_bits_uop_lrs3 = {_RANDOM[10'h12B][31:28], _RANDOM[10'h12C][1:0]};	// lsu.scala:211:16
        stq_1_bits_uop_ldst_val = _RANDOM[10'h12C][2];	// lsu.scala:211:16
        stq_1_bits_uop_dst_rtype = _RANDOM[10'h12C][4:3];	// lsu.scala:211:16
        stq_1_bits_uop_lrs1_rtype = _RANDOM[10'h12C][6:5];	// lsu.scala:211:16
        stq_1_bits_uop_lrs2_rtype = _RANDOM[10'h12C][8:7];	// lsu.scala:211:16
        stq_1_bits_uop_frs3_en = _RANDOM[10'h12C][9];	// lsu.scala:211:16
        stq_1_bits_uop_fp_val = _RANDOM[10'h12C][10];	// lsu.scala:211:16
        stq_1_bits_uop_fp_single = _RANDOM[10'h12C][11];	// lsu.scala:211:16
        stq_1_bits_uop_xcpt_pf_if = _RANDOM[10'h12C][12];	// lsu.scala:211:16
        stq_1_bits_uop_xcpt_ae_if = _RANDOM[10'h12C][13];	// lsu.scala:211:16
        stq_1_bits_uop_xcpt_ma_if = _RANDOM[10'h12C][14];	// lsu.scala:211:16
        stq_1_bits_uop_bp_debug_if = _RANDOM[10'h12C][15];	// lsu.scala:211:16
        stq_1_bits_uop_bp_xcpt_if = _RANDOM[10'h12C][16];	// lsu.scala:211:16
        stq_1_bits_uop_debug_fsrc = _RANDOM[10'h12C][18:17];	// lsu.scala:211:16
        stq_1_bits_uop_debug_tsrc = _RANDOM[10'h12C][20:19];	// lsu.scala:211:16
        stq_1_bits_addr_valid = _RANDOM[10'h12C][21];	// lsu.scala:211:16
        stq_1_bits_addr_bits = {_RANDOM[10'h12C][31:22], _RANDOM[10'h12D][29:0]};	// lsu.scala:211:16
        stq_1_bits_addr_is_virtual = _RANDOM[10'h12D][30];	// lsu.scala:211:16
        stq_1_bits_data_valid = _RANDOM[10'h12D][31];	// lsu.scala:211:16
        stq_1_bits_data_bits = {_RANDOM[10'h12E], _RANDOM[10'h12F]};	// lsu.scala:211:16
        stq_1_bits_committed = _RANDOM[10'h130][0];	// lsu.scala:211:16
        stq_1_bits_succeeded = _RANDOM[10'h130][1];	// lsu.scala:211:16
        stq_2_valid = _RANDOM[10'h132][2];	// lsu.scala:211:16
        stq_2_bits_uop_uopc = _RANDOM[10'h132][9:3];	// lsu.scala:211:16
        stq_2_bits_uop_inst = {_RANDOM[10'h132][31:10], _RANDOM[10'h133][9:0]};	// lsu.scala:211:16
        stq_2_bits_uop_debug_inst = {_RANDOM[10'h133][31:10], _RANDOM[10'h134][9:0]};	// lsu.scala:211:16
        stq_2_bits_uop_is_rvc = _RANDOM[10'h134][10];	// lsu.scala:211:16
        stq_2_bits_uop_debug_pc = {_RANDOM[10'h134][31:11], _RANDOM[10'h135][18:0]};	// lsu.scala:211:16
        stq_2_bits_uop_iq_type = _RANDOM[10'h135][21:19];	// lsu.scala:211:16
        stq_2_bits_uop_fu_code = _RANDOM[10'h135][31:22];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_br_type = _RANDOM[10'h136][3:0];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op1_sel = _RANDOM[10'h136][5:4];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op2_sel = _RANDOM[10'h136][8:6];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_imm_sel = _RANDOM[10'h136][11:9];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_op_fcn = _RANDOM[10'h136][15:12];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_fcn_dw = _RANDOM[10'h136][16];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_csr_cmd = _RANDOM[10'h136][19:17];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_is_load = _RANDOM[10'h136][20];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_is_sta = _RANDOM[10'h136][21];	// lsu.scala:211:16
        stq_2_bits_uop_ctrl_is_std = _RANDOM[10'h136][22];	// lsu.scala:211:16
        stq_2_bits_uop_iw_state = _RANDOM[10'h136][24:23];	// lsu.scala:211:16
        stq_2_bits_uop_iw_p1_poisoned = _RANDOM[10'h136][25];	// lsu.scala:211:16
        stq_2_bits_uop_iw_p2_poisoned = _RANDOM[10'h136][26];	// lsu.scala:211:16
        stq_2_bits_uop_is_br = _RANDOM[10'h136][27];	// lsu.scala:211:16
        stq_2_bits_uop_is_jalr = _RANDOM[10'h136][28];	// lsu.scala:211:16
        stq_2_bits_uop_is_jal = _RANDOM[10'h136][29];	// lsu.scala:211:16
        stq_2_bits_uop_is_sfb = _RANDOM[10'h136][30];	// lsu.scala:211:16
        stq_2_bits_uop_br_mask = {_RANDOM[10'h136][31], _RANDOM[10'h137][10:0]};	// lsu.scala:211:16
        stq_2_bits_uop_br_tag = _RANDOM[10'h137][14:11];	// lsu.scala:211:16
        stq_2_bits_uop_ftq_idx = _RANDOM[10'h137][19:15];	// lsu.scala:211:16
        stq_2_bits_uop_edge_inst = _RANDOM[10'h137][20];	// lsu.scala:211:16
        stq_2_bits_uop_pc_lob = _RANDOM[10'h137][26:21];	// lsu.scala:211:16
        stq_2_bits_uop_taken = _RANDOM[10'h137][27];	// lsu.scala:211:16
        stq_2_bits_uop_imm_packed = {_RANDOM[10'h137][31:28], _RANDOM[10'h138][15:0]};	// lsu.scala:211:16
        stq_2_bits_uop_csr_addr = _RANDOM[10'h138][27:16];	// lsu.scala:211:16
        stq_2_bits_uop_rob_idx = {_RANDOM[10'h138][31:28], _RANDOM[10'h139][1:0]};	// lsu.scala:211:16
        stq_2_bits_uop_ldq_idx = _RANDOM[10'h139][5:2];	// lsu.scala:211:16
        stq_2_bits_uop_stq_idx = _RANDOM[10'h139][9:6];	// lsu.scala:211:16
        stq_2_bits_uop_rxq_idx = _RANDOM[10'h139][11:10];	// lsu.scala:211:16
        stq_2_bits_uop_pdst = _RANDOM[10'h139][18:12];	// lsu.scala:211:16
        stq_2_bits_uop_prs1 = _RANDOM[10'h139][25:19];	// lsu.scala:211:16
        stq_2_bits_uop_prs2 = {_RANDOM[10'h139][31:26], _RANDOM[10'h13A][0]};	// lsu.scala:211:16
        stq_2_bits_uop_prs3 = _RANDOM[10'h13A][7:1];	// lsu.scala:211:16
        stq_2_bits_uop_ppred = _RANDOM[10'h13A][12:8];	// lsu.scala:211:16
        stq_2_bits_uop_prs1_busy = _RANDOM[10'h13A][13];	// lsu.scala:211:16
        stq_2_bits_uop_prs2_busy = _RANDOM[10'h13A][14];	// lsu.scala:211:16
        stq_2_bits_uop_prs3_busy = _RANDOM[10'h13A][15];	// lsu.scala:211:16
        stq_2_bits_uop_ppred_busy = _RANDOM[10'h13A][16];	// lsu.scala:211:16
        stq_2_bits_uop_stale_pdst = _RANDOM[10'h13A][23:17];	// lsu.scala:211:16
        stq_2_bits_uop_exception = _RANDOM[10'h13A][24];	// lsu.scala:211:16
        stq_2_bits_uop_exc_cause =
          {_RANDOM[10'h13A][31:25], _RANDOM[10'h13B], _RANDOM[10'h13C][24:0]};	// lsu.scala:211:16
        stq_2_bits_uop_bypassable = _RANDOM[10'h13C][25];	// lsu.scala:211:16
        stq_2_bits_uop_mem_cmd = _RANDOM[10'h13C][30:26];	// lsu.scala:211:16
        stq_2_bits_uop_mem_size = {_RANDOM[10'h13C][31], _RANDOM[10'h13D][0]};	// lsu.scala:211:16
        stq_2_bits_uop_mem_signed = _RANDOM[10'h13D][1];	// lsu.scala:211:16
        stq_2_bits_uop_is_fence = _RANDOM[10'h13D][2];	// lsu.scala:211:16
        stq_2_bits_uop_is_fencei = _RANDOM[10'h13D][3];	// lsu.scala:211:16
        stq_2_bits_uop_is_amo = _RANDOM[10'h13D][4];	// lsu.scala:211:16
        stq_2_bits_uop_uses_ldq = _RANDOM[10'h13D][5];	// lsu.scala:211:16
        stq_2_bits_uop_uses_stq = _RANDOM[10'h13D][6];	// lsu.scala:211:16
        stq_2_bits_uop_is_sys_pc2epc = _RANDOM[10'h13D][7];	// lsu.scala:211:16
        stq_2_bits_uop_is_unique = _RANDOM[10'h13D][8];	// lsu.scala:211:16
        stq_2_bits_uop_flush_on_commit = _RANDOM[10'h13D][9];	// lsu.scala:211:16
        stq_2_bits_uop_ldst_is_rs1 = _RANDOM[10'h13D][10];	// lsu.scala:211:16
        stq_2_bits_uop_ldst = _RANDOM[10'h13D][16:11];	// lsu.scala:211:16
        stq_2_bits_uop_lrs1 = _RANDOM[10'h13D][22:17];	// lsu.scala:211:16
        stq_2_bits_uop_lrs2 = _RANDOM[10'h13D][28:23];	// lsu.scala:211:16
        stq_2_bits_uop_lrs3 = {_RANDOM[10'h13D][31:29], _RANDOM[10'h13E][2:0]};	// lsu.scala:211:16
        stq_2_bits_uop_ldst_val = _RANDOM[10'h13E][3];	// lsu.scala:211:16
        stq_2_bits_uop_dst_rtype = _RANDOM[10'h13E][5:4];	// lsu.scala:211:16
        stq_2_bits_uop_lrs1_rtype = _RANDOM[10'h13E][7:6];	// lsu.scala:211:16
        stq_2_bits_uop_lrs2_rtype = _RANDOM[10'h13E][9:8];	// lsu.scala:211:16
        stq_2_bits_uop_frs3_en = _RANDOM[10'h13E][10];	// lsu.scala:211:16
        stq_2_bits_uop_fp_val = _RANDOM[10'h13E][11];	// lsu.scala:211:16
        stq_2_bits_uop_fp_single = _RANDOM[10'h13E][12];	// lsu.scala:211:16
        stq_2_bits_uop_xcpt_pf_if = _RANDOM[10'h13E][13];	// lsu.scala:211:16
        stq_2_bits_uop_xcpt_ae_if = _RANDOM[10'h13E][14];	// lsu.scala:211:16
        stq_2_bits_uop_xcpt_ma_if = _RANDOM[10'h13E][15];	// lsu.scala:211:16
        stq_2_bits_uop_bp_debug_if = _RANDOM[10'h13E][16];	// lsu.scala:211:16
        stq_2_bits_uop_bp_xcpt_if = _RANDOM[10'h13E][17];	// lsu.scala:211:16
        stq_2_bits_uop_debug_fsrc = _RANDOM[10'h13E][19:18];	// lsu.scala:211:16
        stq_2_bits_uop_debug_tsrc = _RANDOM[10'h13E][21:20];	// lsu.scala:211:16
        stq_2_bits_addr_valid = _RANDOM[10'h13E][22];	// lsu.scala:211:16
        stq_2_bits_addr_bits = {_RANDOM[10'h13E][31:23], _RANDOM[10'h13F][30:0]};	// lsu.scala:211:16
        stq_2_bits_addr_is_virtual = _RANDOM[10'h13F][31];	// lsu.scala:211:16
        stq_2_bits_data_valid = _RANDOM[10'h140][0];	// lsu.scala:211:16
        stq_2_bits_data_bits =
          {_RANDOM[10'h140][31:1], _RANDOM[10'h141], _RANDOM[10'h142][0]};	// lsu.scala:211:16
        stq_2_bits_committed = _RANDOM[10'h142][1];	// lsu.scala:211:16
        stq_2_bits_succeeded = _RANDOM[10'h142][2];	// lsu.scala:211:16
        stq_3_valid = _RANDOM[10'h144][3];	// lsu.scala:211:16
        stq_3_bits_uop_uopc = _RANDOM[10'h144][10:4];	// lsu.scala:211:16
        stq_3_bits_uop_inst = {_RANDOM[10'h144][31:11], _RANDOM[10'h145][10:0]};	// lsu.scala:211:16
        stq_3_bits_uop_debug_inst = {_RANDOM[10'h145][31:11], _RANDOM[10'h146][10:0]};	// lsu.scala:211:16
        stq_3_bits_uop_is_rvc = _RANDOM[10'h146][11];	// lsu.scala:211:16
        stq_3_bits_uop_debug_pc = {_RANDOM[10'h146][31:12], _RANDOM[10'h147][19:0]};	// lsu.scala:211:16
        stq_3_bits_uop_iq_type = _RANDOM[10'h147][22:20];	// lsu.scala:211:16
        stq_3_bits_uop_fu_code = {_RANDOM[10'h147][31:23], _RANDOM[10'h148][0]};	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_br_type = _RANDOM[10'h148][4:1];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op1_sel = _RANDOM[10'h148][6:5];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op2_sel = _RANDOM[10'h148][9:7];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_imm_sel = _RANDOM[10'h148][12:10];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_op_fcn = _RANDOM[10'h148][16:13];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_fcn_dw = _RANDOM[10'h148][17];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_csr_cmd = _RANDOM[10'h148][20:18];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_is_load = _RANDOM[10'h148][21];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_is_sta = _RANDOM[10'h148][22];	// lsu.scala:211:16
        stq_3_bits_uop_ctrl_is_std = _RANDOM[10'h148][23];	// lsu.scala:211:16
        stq_3_bits_uop_iw_state = _RANDOM[10'h148][25:24];	// lsu.scala:211:16
        stq_3_bits_uop_iw_p1_poisoned = _RANDOM[10'h148][26];	// lsu.scala:211:16
        stq_3_bits_uop_iw_p2_poisoned = _RANDOM[10'h148][27];	// lsu.scala:211:16
        stq_3_bits_uop_is_br = _RANDOM[10'h148][28];	// lsu.scala:211:16
        stq_3_bits_uop_is_jalr = _RANDOM[10'h148][29];	// lsu.scala:211:16
        stq_3_bits_uop_is_jal = _RANDOM[10'h148][30];	// lsu.scala:211:16
        stq_3_bits_uop_is_sfb = _RANDOM[10'h148][31];	// lsu.scala:211:16
        stq_3_bits_uop_br_mask = _RANDOM[10'h149][11:0];	// lsu.scala:211:16
        stq_3_bits_uop_br_tag = _RANDOM[10'h149][15:12];	// lsu.scala:211:16
        stq_3_bits_uop_ftq_idx = _RANDOM[10'h149][20:16];	// lsu.scala:211:16
        stq_3_bits_uop_edge_inst = _RANDOM[10'h149][21];	// lsu.scala:211:16
        stq_3_bits_uop_pc_lob = _RANDOM[10'h149][27:22];	// lsu.scala:211:16
        stq_3_bits_uop_taken = _RANDOM[10'h149][28];	// lsu.scala:211:16
        stq_3_bits_uop_imm_packed = {_RANDOM[10'h149][31:29], _RANDOM[10'h14A][16:0]};	// lsu.scala:211:16
        stq_3_bits_uop_csr_addr = _RANDOM[10'h14A][28:17];	// lsu.scala:211:16
        stq_3_bits_uop_rob_idx = {_RANDOM[10'h14A][31:29], _RANDOM[10'h14B][2:0]};	// lsu.scala:211:16
        stq_3_bits_uop_ldq_idx = _RANDOM[10'h14B][6:3];	// lsu.scala:211:16
        stq_3_bits_uop_stq_idx = _RANDOM[10'h14B][10:7];	// lsu.scala:211:16
        stq_3_bits_uop_rxq_idx = _RANDOM[10'h14B][12:11];	// lsu.scala:211:16
        stq_3_bits_uop_pdst = _RANDOM[10'h14B][19:13];	// lsu.scala:211:16
        stq_3_bits_uop_prs1 = _RANDOM[10'h14B][26:20];	// lsu.scala:211:16
        stq_3_bits_uop_prs2 = {_RANDOM[10'h14B][31:27], _RANDOM[10'h14C][1:0]};	// lsu.scala:211:16
        stq_3_bits_uop_prs3 = _RANDOM[10'h14C][8:2];	// lsu.scala:211:16
        stq_3_bits_uop_ppred = _RANDOM[10'h14C][13:9];	// lsu.scala:211:16
        stq_3_bits_uop_prs1_busy = _RANDOM[10'h14C][14];	// lsu.scala:211:16
        stq_3_bits_uop_prs2_busy = _RANDOM[10'h14C][15];	// lsu.scala:211:16
        stq_3_bits_uop_prs3_busy = _RANDOM[10'h14C][16];	// lsu.scala:211:16
        stq_3_bits_uop_ppred_busy = _RANDOM[10'h14C][17];	// lsu.scala:211:16
        stq_3_bits_uop_stale_pdst = _RANDOM[10'h14C][24:18];	// lsu.scala:211:16
        stq_3_bits_uop_exception = _RANDOM[10'h14C][25];	// lsu.scala:211:16
        stq_3_bits_uop_exc_cause =
          {_RANDOM[10'h14C][31:26], _RANDOM[10'h14D], _RANDOM[10'h14E][25:0]};	// lsu.scala:211:16
        stq_3_bits_uop_bypassable = _RANDOM[10'h14E][26];	// lsu.scala:211:16
        stq_3_bits_uop_mem_cmd = _RANDOM[10'h14E][31:27];	// lsu.scala:211:16
        stq_3_bits_uop_mem_size = _RANDOM[10'h14F][1:0];	// lsu.scala:211:16
        stq_3_bits_uop_mem_signed = _RANDOM[10'h14F][2];	// lsu.scala:211:16
        stq_3_bits_uop_is_fence = _RANDOM[10'h14F][3];	// lsu.scala:211:16
        stq_3_bits_uop_is_fencei = _RANDOM[10'h14F][4];	// lsu.scala:211:16
        stq_3_bits_uop_is_amo = _RANDOM[10'h14F][5];	// lsu.scala:211:16
        stq_3_bits_uop_uses_ldq = _RANDOM[10'h14F][6];	// lsu.scala:211:16
        stq_3_bits_uop_uses_stq = _RANDOM[10'h14F][7];	// lsu.scala:211:16
        stq_3_bits_uop_is_sys_pc2epc = _RANDOM[10'h14F][8];	// lsu.scala:211:16
        stq_3_bits_uop_is_unique = _RANDOM[10'h14F][9];	// lsu.scala:211:16
        stq_3_bits_uop_flush_on_commit = _RANDOM[10'h14F][10];	// lsu.scala:211:16
        stq_3_bits_uop_ldst_is_rs1 = _RANDOM[10'h14F][11];	// lsu.scala:211:16
        stq_3_bits_uop_ldst = _RANDOM[10'h14F][17:12];	// lsu.scala:211:16
        stq_3_bits_uop_lrs1 = _RANDOM[10'h14F][23:18];	// lsu.scala:211:16
        stq_3_bits_uop_lrs2 = _RANDOM[10'h14F][29:24];	// lsu.scala:211:16
        stq_3_bits_uop_lrs3 = {_RANDOM[10'h14F][31:30], _RANDOM[10'h150][3:0]};	// lsu.scala:211:16
        stq_3_bits_uop_ldst_val = _RANDOM[10'h150][4];	// lsu.scala:211:16
        stq_3_bits_uop_dst_rtype = _RANDOM[10'h150][6:5];	// lsu.scala:211:16
        stq_3_bits_uop_lrs1_rtype = _RANDOM[10'h150][8:7];	// lsu.scala:211:16
        stq_3_bits_uop_lrs2_rtype = _RANDOM[10'h150][10:9];	// lsu.scala:211:16
        stq_3_bits_uop_frs3_en = _RANDOM[10'h150][11];	// lsu.scala:211:16
        stq_3_bits_uop_fp_val = _RANDOM[10'h150][12];	// lsu.scala:211:16
        stq_3_bits_uop_fp_single = _RANDOM[10'h150][13];	// lsu.scala:211:16
        stq_3_bits_uop_xcpt_pf_if = _RANDOM[10'h150][14];	// lsu.scala:211:16
        stq_3_bits_uop_xcpt_ae_if = _RANDOM[10'h150][15];	// lsu.scala:211:16
        stq_3_bits_uop_xcpt_ma_if = _RANDOM[10'h150][16];	// lsu.scala:211:16
        stq_3_bits_uop_bp_debug_if = _RANDOM[10'h150][17];	// lsu.scala:211:16
        stq_3_bits_uop_bp_xcpt_if = _RANDOM[10'h150][18];	// lsu.scala:211:16
        stq_3_bits_uop_debug_fsrc = _RANDOM[10'h150][20:19];	// lsu.scala:211:16
        stq_3_bits_uop_debug_tsrc = _RANDOM[10'h150][22:21];	// lsu.scala:211:16
        stq_3_bits_addr_valid = _RANDOM[10'h150][23];	// lsu.scala:211:16
        stq_3_bits_addr_bits = {_RANDOM[10'h150][31:24], _RANDOM[10'h151]};	// lsu.scala:211:16
        stq_3_bits_addr_is_virtual = _RANDOM[10'h152][0];	// lsu.scala:211:16
        stq_3_bits_data_valid = _RANDOM[10'h152][1];	// lsu.scala:211:16
        stq_3_bits_data_bits =
          {_RANDOM[10'h152][31:2], _RANDOM[10'h153], _RANDOM[10'h154][1:0]};	// lsu.scala:211:16
        stq_3_bits_committed = _RANDOM[10'h154][2];	// lsu.scala:211:16
        stq_3_bits_succeeded = _RANDOM[10'h154][3];	// lsu.scala:211:16
        stq_4_valid = _RANDOM[10'h156][4];	// lsu.scala:211:16
        stq_4_bits_uop_uopc = _RANDOM[10'h156][11:5];	// lsu.scala:211:16
        stq_4_bits_uop_inst = {_RANDOM[10'h156][31:12], _RANDOM[10'h157][11:0]};	// lsu.scala:211:16
        stq_4_bits_uop_debug_inst = {_RANDOM[10'h157][31:12], _RANDOM[10'h158][11:0]};	// lsu.scala:211:16
        stq_4_bits_uop_is_rvc = _RANDOM[10'h158][12];	// lsu.scala:211:16
        stq_4_bits_uop_debug_pc = {_RANDOM[10'h158][31:13], _RANDOM[10'h159][20:0]};	// lsu.scala:211:16
        stq_4_bits_uop_iq_type = _RANDOM[10'h159][23:21];	// lsu.scala:211:16
        stq_4_bits_uop_fu_code = {_RANDOM[10'h159][31:24], _RANDOM[10'h15A][1:0]};	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_br_type = _RANDOM[10'h15A][5:2];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op1_sel = _RANDOM[10'h15A][7:6];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op2_sel = _RANDOM[10'h15A][10:8];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_imm_sel = _RANDOM[10'h15A][13:11];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_op_fcn = _RANDOM[10'h15A][17:14];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_fcn_dw = _RANDOM[10'h15A][18];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_csr_cmd = _RANDOM[10'h15A][21:19];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_is_load = _RANDOM[10'h15A][22];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_is_sta = _RANDOM[10'h15A][23];	// lsu.scala:211:16
        stq_4_bits_uop_ctrl_is_std = _RANDOM[10'h15A][24];	// lsu.scala:211:16
        stq_4_bits_uop_iw_state = _RANDOM[10'h15A][26:25];	// lsu.scala:211:16
        stq_4_bits_uop_iw_p1_poisoned = _RANDOM[10'h15A][27];	// lsu.scala:211:16
        stq_4_bits_uop_iw_p2_poisoned = _RANDOM[10'h15A][28];	// lsu.scala:211:16
        stq_4_bits_uop_is_br = _RANDOM[10'h15A][29];	// lsu.scala:211:16
        stq_4_bits_uop_is_jalr = _RANDOM[10'h15A][30];	// lsu.scala:211:16
        stq_4_bits_uop_is_jal = _RANDOM[10'h15A][31];	// lsu.scala:211:16
        stq_4_bits_uop_is_sfb = _RANDOM[10'h15B][0];	// lsu.scala:211:16
        stq_4_bits_uop_br_mask = _RANDOM[10'h15B][12:1];	// lsu.scala:211:16
        stq_4_bits_uop_br_tag = _RANDOM[10'h15B][16:13];	// lsu.scala:211:16
        stq_4_bits_uop_ftq_idx = _RANDOM[10'h15B][21:17];	// lsu.scala:211:16
        stq_4_bits_uop_edge_inst = _RANDOM[10'h15B][22];	// lsu.scala:211:16
        stq_4_bits_uop_pc_lob = _RANDOM[10'h15B][28:23];	// lsu.scala:211:16
        stq_4_bits_uop_taken = _RANDOM[10'h15B][29];	// lsu.scala:211:16
        stq_4_bits_uop_imm_packed = {_RANDOM[10'h15B][31:30], _RANDOM[10'h15C][17:0]};	// lsu.scala:211:16
        stq_4_bits_uop_csr_addr = _RANDOM[10'h15C][29:18];	// lsu.scala:211:16
        stq_4_bits_uop_rob_idx = {_RANDOM[10'h15C][31:30], _RANDOM[10'h15D][3:0]};	// lsu.scala:211:16
        stq_4_bits_uop_ldq_idx = _RANDOM[10'h15D][7:4];	// lsu.scala:211:16
        stq_4_bits_uop_stq_idx = _RANDOM[10'h15D][11:8];	// lsu.scala:211:16
        stq_4_bits_uop_rxq_idx = _RANDOM[10'h15D][13:12];	// lsu.scala:211:16
        stq_4_bits_uop_pdst = _RANDOM[10'h15D][20:14];	// lsu.scala:211:16
        stq_4_bits_uop_prs1 = _RANDOM[10'h15D][27:21];	// lsu.scala:211:16
        stq_4_bits_uop_prs2 = {_RANDOM[10'h15D][31:28], _RANDOM[10'h15E][2:0]};	// lsu.scala:211:16
        stq_4_bits_uop_prs3 = _RANDOM[10'h15E][9:3];	// lsu.scala:211:16
        stq_4_bits_uop_ppred = _RANDOM[10'h15E][14:10];	// lsu.scala:211:16
        stq_4_bits_uop_prs1_busy = _RANDOM[10'h15E][15];	// lsu.scala:211:16
        stq_4_bits_uop_prs2_busy = _RANDOM[10'h15E][16];	// lsu.scala:211:16
        stq_4_bits_uop_prs3_busy = _RANDOM[10'h15E][17];	// lsu.scala:211:16
        stq_4_bits_uop_ppred_busy = _RANDOM[10'h15E][18];	// lsu.scala:211:16
        stq_4_bits_uop_stale_pdst = _RANDOM[10'h15E][25:19];	// lsu.scala:211:16
        stq_4_bits_uop_exception = _RANDOM[10'h15E][26];	// lsu.scala:211:16
        stq_4_bits_uop_exc_cause =
          {_RANDOM[10'h15E][31:27], _RANDOM[10'h15F], _RANDOM[10'h160][26:0]};	// lsu.scala:211:16
        stq_4_bits_uop_bypassable = _RANDOM[10'h160][27];	// lsu.scala:211:16
        stq_4_bits_uop_mem_cmd = {_RANDOM[10'h160][31:28], _RANDOM[10'h161][0]};	// lsu.scala:211:16
        stq_4_bits_uop_mem_size = _RANDOM[10'h161][2:1];	// lsu.scala:211:16
        stq_4_bits_uop_mem_signed = _RANDOM[10'h161][3];	// lsu.scala:211:16
        stq_4_bits_uop_is_fence = _RANDOM[10'h161][4];	// lsu.scala:211:16
        stq_4_bits_uop_is_fencei = _RANDOM[10'h161][5];	// lsu.scala:211:16
        stq_4_bits_uop_is_amo = _RANDOM[10'h161][6];	// lsu.scala:211:16
        stq_4_bits_uop_uses_ldq = _RANDOM[10'h161][7];	// lsu.scala:211:16
        stq_4_bits_uop_uses_stq = _RANDOM[10'h161][8];	// lsu.scala:211:16
        stq_4_bits_uop_is_sys_pc2epc = _RANDOM[10'h161][9];	// lsu.scala:211:16
        stq_4_bits_uop_is_unique = _RANDOM[10'h161][10];	// lsu.scala:211:16
        stq_4_bits_uop_flush_on_commit = _RANDOM[10'h161][11];	// lsu.scala:211:16
        stq_4_bits_uop_ldst_is_rs1 = _RANDOM[10'h161][12];	// lsu.scala:211:16
        stq_4_bits_uop_ldst = _RANDOM[10'h161][18:13];	// lsu.scala:211:16
        stq_4_bits_uop_lrs1 = _RANDOM[10'h161][24:19];	// lsu.scala:211:16
        stq_4_bits_uop_lrs2 = _RANDOM[10'h161][30:25];	// lsu.scala:211:16
        stq_4_bits_uop_lrs3 = {_RANDOM[10'h161][31], _RANDOM[10'h162][4:0]};	// lsu.scala:211:16
        stq_4_bits_uop_ldst_val = _RANDOM[10'h162][5];	// lsu.scala:211:16
        stq_4_bits_uop_dst_rtype = _RANDOM[10'h162][7:6];	// lsu.scala:211:16
        stq_4_bits_uop_lrs1_rtype = _RANDOM[10'h162][9:8];	// lsu.scala:211:16
        stq_4_bits_uop_lrs2_rtype = _RANDOM[10'h162][11:10];	// lsu.scala:211:16
        stq_4_bits_uop_frs3_en = _RANDOM[10'h162][12];	// lsu.scala:211:16
        stq_4_bits_uop_fp_val = _RANDOM[10'h162][13];	// lsu.scala:211:16
        stq_4_bits_uop_fp_single = _RANDOM[10'h162][14];	// lsu.scala:211:16
        stq_4_bits_uop_xcpt_pf_if = _RANDOM[10'h162][15];	// lsu.scala:211:16
        stq_4_bits_uop_xcpt_ae_if = _RANDOM[10'h162][16];	// lsu.scala:211:16
        stq_4_bits_uop_xcpt_ma_if = _RANDOM[10'h162][17];	// lsu.scala:211:16
        stq_4_bits_uop_bp_debug_if = _RANDOM[10'h162][18];	// lsu.scala:211:16
        stq_4_bits_uop_bp_xcpt_if = _RANDOM[10'h162][19];	// lsu.scala:211:16
        stq_4_bits_uop_debug_fsrc = _RANDOM[10'h162][21:20];	// lsu.scala:211:16
        stq_4_bits_uop_debug_tsrc = _RANDOM[10'h162][23:22];	// lsu.scala:211:16
        stq_4_bits_addr_valid = _RANDOM[10'h162][24];	// lsu.scala:211:16
        stq_4_bits_addr_bits =
          {_RANDOM[10'h162][31:25], _RANDOM[10'h163], _RANDOM[10'h164][0]};	// lsu.scala:211:16
        stq_4_bits_addr_is_virtual = _RANDOM[10'h164][1];	// lsu.scala:211:16
        stq_4_bits_data_valid = _RANDOM[10'h164][2];	// lsu.scala:211:16
        stq_4_bits_data_bits =
          {_RANDOM[10'h164][31:3], _RANDOM[10'h165], _RANDOM[10'h166][2:0]};	// lsu.scala:211:16
        stq_4_bits_committed = _RANDOM[10'h166][3];	// lsu.scala:211:16
        stq_4_bits_succeeded = _RANDOM[10'h166][4];	// lsu.scala:211:16
        stq_5_valid = _RANDOM[10'h168][5];	// lsu.scala:211:16
        stq_5_bits_uop_uopc = _RANDOM[10'h168][12:6];	// lsu.scala:211:16
        stq_5_bits_uop_inst = {_RANDOM[10'h168][31:13], _RANDOM[10'h169][12:0]};	// lsu.scala:211:16
        stq_5_bits_uop_debug_inst = {_RANDOM[10'h169][31:13], _RANDOM[10'h16A][12:0]};	// lsu.scala:211:16
        stq_5_bits_uop_is_rvc = _RANDOM[10'h16A][13];	// lsu.scala:211:16
        stq_5_bits_uop_debug_pc = {_RANDOM[10'h16A][31:14], _RANDOM[10'h16B][21:0]};	// lsu.scala:211:16
        stq_5_bits_uop_iq_type = _RANDOM[10'h16B][24:22];	// lsu.scala:211:16
        stq_5_bits_uop_fu_code = {_RANDOM[10'h16B][31:25], _RANDOM[10'h16C][2:0]};	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_br_type = _RANDOM[10'h16C][6:3];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op1_sel = _RANDOM[10'h16C][8:7];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op2_sel = _RANDOM[10'h16C][11:9];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_imm_sel = _RANDOM[10'h16C][14:12];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_op_fcn = _RANDOM[10'h16C][18:15];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_fcn_dw = _RANDOM[10'h16C][19];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_csr_cmd = _RANDOM[10'h16C][22:20];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_is_load = _RANDOM[10'h16C][23];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_is_sta = _RANDOM[10'h16C][24];	// lsu.scala:211:16
        stq_5_bits_uop_ctrl_is_std = _RANDOM[10'h16C][25];	// lsu.scala:211:16
        stq_5_bits_uop_iw_state = _RANDOM[10'h16C][27:26];	// lsu.scala:211:16
        stq_5_bits_uop_iw_p1_poisoned = _RANDOM[10'h16C][28];	// lsu.scala:211:16
        stq_5_bits_uop_iw_p2_poisoned = _RANDOM[10'h16C][29];	// lsu.scala:211:16
        stq_5_bits_uop_is_br = _RANDOM[10'h16C][30];	// lsu.scala:211:16
        stq_5_bits_uop_is_jalr = _RANDOM[10'h16C][31];	// lsu.scala:211:16
        stq_5_bits_uop_is_jal = _RANDOM[10'h16D][0];	// lsu.scala:211:16
        stq_5_bits_uop_is_sfb = _RANDOM[10'h16D][1];	// lsu.scala:211:16
        stq_5_bits_uop_br_mask = _RANDOM[10'h16D][13:2];	// lsu.scala:211:16
        stq_5_bits_uop_br_tag = _RANDOM[10'h16D][17:14];	// lsu.scala:211:16
        stq_5_bits_uop_ftq_idx = _RANDOM[10'h16D][22:18];	// lsu.scala:211:16
        stq_5_bits_uop_edge_inst = _RANDOM[10'h16D][23];	// lsu.scala:211:16
        stq_5_bits_uop_pc_lob = _RANDOM[10'h16D][29:24];	// lsu.scala:211:16
        stq_5_bits_uop_taken = _RANDOM[10'h16D][30];	// lsu.scala:211:16
        stq_5_bits_uop_imm_packed = {_RANDOM[10'h16D][31], _RANDOM[10'h16E][18:0]};	// lsu.scala:211:16
        stq_5_bits_uop_csr_addr = _RANDOM[10'h16E][30:19];	// lsu.scala:211:16
        stq_5_bits_uop_rob_idx = {_RANDOM[10'h16E][31], _RANDOM[10'h16F][4:0]};	// lsu.scala:211:16
        stq_5_bits_uop_ldq_idx = _RANDOM[10'h16F][8:5];	// lsu.scala:211:16
        stq_5_bits_uop_stq_idx = _RANDOM[10'h16F][12:9];	// lsu.scala:211:16
        stq_5_bits_uop_rxq_idx = _RANDOM[10'h16F][14:13];	// lsu.scala:211:16
        stq_5_bits_uop_pdst = _RANDOM[10'h16F][21:15];	// lsu.scala:211:16
        stq_5_bits_uop_prs1 = _RANDOM[10'h16F][28:22];	// lsu.scala:211:16
        stq_5_bits_uop_prs2 = {_RANDOM[10'h16F][31:29], _RANDOM[10'h170][3:0]};	// lsu.scala:211:16
        stq_5_bits_uop_prs3 = _RANDOM[10'h170][10:4];	// lsu.scala:211:16
        stq_5_bits_uop_ppred = _RANDOM[10'h170][15:11];	// lsu.scala:211:16
        stq_5_bits_uop_prs1_busy = _RANDOM[10'h170][16];	// lsu.scala:211:16
        stq_5_bits_uop_prs2_busy = _RANDOM[10'h170][17];	// lsu.scala:211:16
        stq_5_bits_uop_prs3_busy = _RANDOM[10'h170][18];	// lsu.scala:211:16
        stq_5_bits_uop_ppred_busy = _RANDOM[10'h170][19];	// lsu.scala:211:16
        stq_5_bits_uop_stale_pdst = _RANDOM[10'h170][26:20];	// lsu.scala:211:16
        stq_5_bits_uop_exception = _RANDOM[10'h170][27];	// lsu.scala:211:16
        stq_5_bits_uop_exc_cause =
          {_RANDOM[10'h170][31:28], _RANDOM[10'h171], _RANDOM[10'h172][27:0]};	// lsu.scala:211:16
        stq_5_bits_uop_bypassable = _RANDOM[10'h172][28];	// lsu.scala:211:16
        stq_5_bits_uop_mem_cmd = {_RANDOM[10'h172][31:29], _RANDOM[10'h173][1:0]};	// lsu.scala:211:16
        stq_5_bits_uop_mem_size = _RANDOM[10'h173][3:2];	// lsu.scala:211:16
        stq_5_bits_uop_mem_signed = _RANDOM[10'h173][4];	// lsu.scala:211:16
        stq_5_bits_uop_is_fence = _RANDOM[10'h173][5];	// lsu.scala:211:16
        stq_5_bits_uop_is_fencei = _RANDOM[10'h173][6];	// lsu.scala:211:16
        stq_5_bits_uop_is_amo = _RANDOM[10'h173][7];	// lsu.scala:211:16
        stq_5_bits_uop_uses_ldq = _RANDOM[10'h173][8];	// lsu.scala:211:16
        stq_5_bits_uop_uses_stq = _RANDOM[10'h173][9];	// lsu.scala:211:16
        stq_5_bits_uop_is_sys_pc2epc = _RANDOM[10'h173][10];	// lsu.scala:211:16
        stq_5_bits_uop_is_unique = _RANDOM[10'h173][11];	// lsu.scala:211:16
        stq_5_bits_uop_flush_on_commit = _RANDOM[10'h173][12];	// lsu.scala:211:16
        stq_5_bits_uop_ldst_is_rs1 = _RANDOM[10'h173][13];	// lsu.scala:211:16
        stq_5_bits_uop_ldst = _RANDOM[10'h173][19:14];	// lsu.scala:211:16
        stq_5_bits_uop_lrs1 = _RANDOM[10'h173][25:20];	// lsu.scala:211:16
        stq_5_bits_uop_lrs2 = _RANDOM[10'h173][31:26];	// lsu.scala:211:16
        stq_5_bits_uop_lrs3 = _RANDOM[10'h174][5:0];	// lsu.scala:211:16
        stq_5_bits_uop_ldst_val = _RANDOM[10'h174][6];	// lsu.scala:211:16
        stq_5_bits_uop_dst_rtype = _RANDOM[10'h174][8:7];	// lsu.scala:211:16
        stq_5_bits_uop_lrs1_rtype = _RANDOM[10'h174][10:9];	// lsu.scala:211:16
        stq_5_bits_uop_lrs2_rtype = _RANDOM[10'h174][12:11];	// lsu.scala:211:16
        stq_5_bits_uop_frs3_en = _RANDOM[10'h174][13];	// lsu.scala:211:16
        stq_5_bits_uop_fp_val = _RANDOM[10'h174][14];	// lsu.scala:211:16
        stq_5_bits_uop_fp_single = _RANDOM[10'h174][15];	// lsu.scala:211:16
        stq_5_bits_uop_xcpt_pf_if = _RANDOM[10'h174][16];	// lsu.scala:211:16
        stq_5_bits_uop_xcpt_ae_if = _RANDOM[10'h174][17];	// lsu.scala:211:16
        stq_5_bits_uop_xcpt_ma_if = _RANDOM[10'h174][18];	// lsu.scala:211:16
        stq_5_bits_uop_bp_debug_if = _RANDOM[10'h174][19];	// lsu.scala:211:16
        stq_5_bits_uop_bp_xcpt_if = _RANDOM[10'h174][20];	// lsu.scala:211:16
        stq_5_bits_uop_debug_fsrc = _RANDOM[10'h174][22:21];	// lsu.scala:211:16
        stq_5_bits_uop_debug_tsrc = _RANDOM[10'h174][24:23];	// lsu.scala:211:16
        stq_5_bits_addr_valid = _RANDOM[10'h174][25];	// lsu.scala:211:16
        stq_5_bits_addr_bits =
          {_RANDOM[10'h174][31:26], _RANDOM[10'h175], _RANDOM[10'h176][1:0]};	// lsu.scala:211:16
        stq_5_bits_addr_is_virtual = _RANDOM[10'h176][2];	// lsu.scala:211:16
        stq_5_bits_data_valid = _RANDOM[10'h176][3];	// lsu.scala:211:16
        stq_5_bits_data_bits =
          {_RANDOM[10'h176][31:4], _RANDOM[10'h177], _RANDOM[10'h178][3:0]};	// lsu.scala:211:16
        stq_5_bits_committed = _RANDOM[10'h178][4];	// lsu.scala:211:16
        stq_5_bits_succeeded = _RANDOM[10'h178][5];	// lsu.scala:211:16
        stq_6_valid = _RANDOM[10'h17A][6];	// lsu.scala:211:16
        stq_6_bits_uop_uopc = _RANDOM[10'h17A][13:7];	// lsu.scala:211:16
        stq_6_bits_uop_inst = {_RANDOM[10'h17A][31:14], _RANDOM[10'h17B][13:0]};	// lsu.scala:211:16
        stq_6_bits_uop_debug_inst = {_RANDOM[10'h17B][31:14], _RANDOM[10'h17C][13:0]};	// lsu.scala:211:16
        stq_6_bits_uop_is_rvc = _RANDOM[10'h17C][14];	// lsu.scala:211:16
        stq_6_bits_uop_debug_pc = {_RANDOM[10'h17C][31:15], _RANDOM[10'h17D][22:0]};	// lsu.scala:211:16
        stq_6_bits_uop_iq_type = _RANDOM[10'h17D][25:23];	// lsu.scala:211:16
        stq_6_bits_uop_fu_code = {_RANDOM[10'h17D][31:26], _RANDOM[10'h17E][3:0]};	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_br_type = _RANDOM[10'h17E][7:4];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op1_sel = _RANDOM[10'h17E][9:8];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op2_sel = _RANDOM[10'h17E][12:10];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_imm_sel = _RANDOM[10'h17E][15:13];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_op_fcn = _RANDOM[10'h17E][19:16];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_fcn_dw = _RANDOM[10'h17E][20];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_csr_cmd = _RANDOM[10'h17E][23:21];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_is_load = _RANDOM[10'h17E][24];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_is_sta = _RANDOM[10'h17E][25];	// lsu.scala:211:16
        stq_6_bits_uop_ctrl_is_std = _RANDOM[10'h17E][26];	// lsu.scala:211:16
        stq_6_bits_uop_iw_state = _RANDOM[10'h17E][28:27];	// lsu.scala:211:16
        stq_6_bits_uop_iw_p1_poisoned = _RANDOM[10'h17E][29];	// lsu.scala:211:16
        stq_6_bits_uop_iw_p2_poisoned = _RANDOM[10'h17E][30];	// lsu.scala:211:16
        stq_6_bits_uop_is_br = _RANDOM[10'h17E][31];	// lsu.scala:211:16
        stq_6_bits_uop_is_jalr = _RANDOM[10'h17F][0];	// lsu.scala:211:16
        stq_6_bits_uop_is_jal = _RANDOM[10'h17F][1];	// lsu.scala:211:16
        stq_6_bits_uop_is_sfb = _RANDOM[10'h17F][2];	// lsu.scala:211:16
        stq_6_bits_uop_br_mask = _RANDOM[10'h17F][14:3];	// lsu.scala:211:16
        stq_6_bits_uop_br_tag = _RANDOM[10'h17F][18:15];	// lsu.scala:211:16
        stq_6_bits_uop_ftq_idx = _RANDOM[10'h17F][23:19];	// lsu.scala:211:16
        stq_6_bits_uop_edge_inst = _RANDOM[10'h17F][24];	// lsu.scala:211:16
        stq_6_bits_uop_pc_lob = _RANDOM[10'h17F][30:25];	// lsu.scala:211:16
        stq_6_bits_uop_taken = _RANDOM[10'h17F][31];	// lsu.scala:211:16
        stq_6_bits_uop_imm_packed = _RANDOM[10'h180][19:0];	// lsu.scala:211:16
        stq_6_bits_uop_csr_addr = _RANDOM[10'h180][31:20];	// lsu.scala:211:16
        stq_6_bits_uop_rob_idx = _RANDOM[10'h181][5:0];	// lsu.scala:211:16
        stq_6_bits_uop_ldq_idx = _RANDOM[10'h181][9:6];	// lsu.scala:211:16
        stq_6_bits_uop_stq_idx = _RANDOM[10'h181][13:10];	// lsu.scala:211:16
        stq_6_bits_uop_rxq_idx = _RANDOM[10'h181][15:14];	// lsu.scala:211:16
        stq_6_bits_uop_pdst = _RANDOM[10'h181][22:16];	// lsu.scala:211:16
        stq_6_bits_uop_prs1 = _RANDOM[10'h181][29:23];	// lsu.scala:211:16
        stq_6_bits_uop_prs2 = {_RANDOM[10'h181][31:30], _RANDOM[10'h182][4:0]};	// lsu.scala:211:16
        stq_6_bits_uop_prs3 = _RANDOM[10'h182][11:5];	// lsu.scala:211:16
        stq_6_bits_uop_ppred = _RANDOM[10'h182][16:12];	// lsu.scala:211:16
        stq_6_bits_uop_prs1_busy = _RANDOM[10'h182][17];	// lsu.scala:211:16
        stq_6_bits_uop_prs2_busy = _RANDOM[10'h182][18];	// lsu.scala:211:16
        stq_6_bits_uop_prs3_busy = _RANDOM[10'h182][19];	// lsu.scala:211:16
        stq_6_bits_uop_ppred_busy = _RANDOM[10'h182][20];	// lsu.scala:211:16
        stq_6_bits_uop_stale_pdst = _RANDOM[10'h182][27:21];	// lsu.scala:211:16
        stq_6_bits_uop_exception = _RANDOM[10'h182][28];	// lsu.scala:211:16
        stq_6_bits_uop_exc_cause =
          {_RANDOM[10'h182][31:29], _RANDOM[10'h183], _RANDOM[10'h184][28:0]};	// lsu.scala:211:16
        stq_6_bits_uop_bypassable = _RANDOM[10'h184][29];	// lsu.scala:211:16
        stq_6_bits_uop_mem_cmd = {_RANDOM[10'h184][31:30], _RANDOM[10'h185][2:0]};	// lsu.scala:211:16
        stq_6_bits_uop_mem_size = _RANDOM[10'h185][4:3];	// lsu.scala:211:16
        stq_6_bits_uop_mem_signed = _RANDOM[10'h185][5];	// lsu.scala:211:16
        stq_6_bits_uop_is_fence = _RANDOM[10'h185][6];	// lsu.scala:211:16
        stq_6_bits_uop_is_fencei = _RANDOM[10'h185][7];	// lsu.scala:211:16
        stq_6_bits_uop_is_amo = _RANDOM[10'h185][8];	// lsu.scala:211:16
        stq_6_bits_uop_uses_ldq = _RANDOM[10'h185][9];	// lsu.scala:211:16
        stq_6_bits_uop_uses_stq = _RANDOM[10'h185][10];	// lsu.scala:211:16
        stq_6_bits_uop_is_sys_pc2epc = _RANDOM[10'h185][11];	// lsu.scala:211:16
        stq_6_bits_uop_is_unique = _RANDOM[10'h185][12];	// lsu.scala:211:16
        stq_6_bits_uop_flush_on_commit = _RANDOM[10'h185][13];	// lsu.scala:211:16
        stq_6_bits_uop_ldst_is_rs1 = _RANDOM[10'h185][14];	// lsu.scala:211:16
        stq_6_bits_uop_ldst = _RANDOM[10'h185][20:15];	// lsu.scala:211:16
        stq_6_bits_uop_lrs1 = _RANDOM[10'h185][26:21];	// lsu.scala:211:16
        stq_6_bits_uop_lrs2 = {_RANDOM[10'h185][31:27], _RANDOM[10'h186][0]};	// lsu.scala:211:16
        stq_6_bits_uop_lrs3 = _RANDOM[10'h186][6:1];	// lsu.scala:211:16
        stq_6_bits_uop_ldst_val = _RANDOM[10'h186][7];	// lsu.scala:211:16
        stq_6_bits_uop_dst_rtype = _RANDOM[10'h186][9:8];	// lsu.scala:211:16
        stq_6_bits_uop_lrs1_rtype = _RANDOM[10'h186][11:10];	// lsu.scala:211:16
        stq_6_bits_uop_lrs2_rtype = _RANDOM[10'h186][13:12];	// lsu.scala:211:16
        stq_6_bits_uop_frs3_en = _RANDOM[10'h186][14];	// lsu.scala:211:16
        stq_6_bits_uop_fp_val = _RANDOM[10'h186][15];	// lsu.scala:211:16
        stq_6_bits_uop_fp_single = _RANDOM[10'h186][16];	// lsu.scala:211:16
        stq_6_bits_uop_xcpt_pf_if = _RANDOM[10'h186][17];	// lsu.scala:211:16
        stq_6_bits_uop_xcpt_ae_if = _RANDOM[10'h186][18];	// lsu.scala:211:16
        stq_6_bits_uop_xcpt_ma_if = _RANDOM[10'h186][19];	// lsu.scala:211:16
        stq_6_bits_uop_bp_debug_if = _RANDOM[10'h186][20];	// lsu.scala:211:16
        stq_6_bits_uop_bp_xcpt_if = _RANDOM[10'h186][21];	// lsu.scala:211:16
        stq_6_bits_uop_debug_fsrc = _RANDOM[10'h186][23:22];	// lsu.scala:211:16
        stq_6_bits_uop_debug_tsrc = _RANDOM[10'h186][25:24];	// lsu.scala:211:16
        stq_6_bits_addr_valid = _RANDOM[10'h186][26];	// lsu.scala:211:16
        stq_6_bits_addr_bits =
          {_RANDOM[10'h186][31:27], _RANDOM[10'h187], _RANDOM[10'h188][2:0]};	// lsu.scala:211:16
        stq_6_bits_addr_is_virtual = _RANDOM[10'h188][3];	// lsu.scala:211:16
        stq_6_bits_data_valid = _RANDOM[10'h188][4];	// lsu.scala:211:16
        stq_6_bits_data_bits =
          {_RANDOM[10'h188][31:5], _RANDOM[10'h189], _RANDOM[10'h18A][4:0]};	// lsu.scala:211:16
        stq_6_bits_committed = _RANDOM[10'h18A][5];	// lsu.scala:211:16
        stq_6_bits_succeeded = _RANDOM[10'h18A][6];	// lsu.scala:211:16
        stq_7_valid = _RANDOM[10'h18C][7];	// lsu.scala:211:16
        stq_7_bits_uop_uopc = _RANDOM[10'h18C][14:8];	// lsu.scala:211:16
        stq_7_bits_uop_inst = {_RANDOM[10'h18C][31:15], _RANDOM[10'h18D][14:0]};	// lsu.scala:211:16
        stq_7_bits_uop_debug_inst = {_RANDOM[10'h18D][31:15], _RANDOM[10'h18E][14:0]};	// lsu.scala:211:16
        stq_7_bits_uop_is_rvc = _RANDOM[10'h18E][15];	// lsu.scala:211:16
        stq_7_bits_uop_debug_pc = {_RANDOM[10'h18E][31:16], _RANDOM[10'h18F][23:0]};	// lsu.scala:211:16
        stq_7_bits_uop_iq_type = _RANDOM[10'h18F][26:24];	// lsu.scala:211:16
        stq_7_bits_uop_fu_code = {_RANDOM[10'h18F][31:27], _RANDOM[10'h190][4:0]};	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_br_type = _RANDOM[10'h190][8:5];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op1_sel = _RANDOM[10'h190][10:9];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op2_sel = _RANDOM[10'h190][13:11];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_imm_sel = _RANDOM[10'h190][16:14];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_op_fcn = _RANDOM[10'h190][20:17];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_fcn_dw = _RANDOM[10'h190][21];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_csr_cmd = _RANDOM[10'h190][24:22];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_is_load = _RANDOM[10'h190][25];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_is_sta = _RANDOM[10'h190][26];	// lsu.scala:211:16
        stq_7_bits_uop_ctrl_is_std = _RANDOM[10'h190][27];	// lsu.scala:211:16
        stq_7_bits_uop_iw_state = _RANDOM[10'h190][29:28];	// lsu.scala:211:16
        stq_7_bits_uop_iw_p1_poisoned = _RANDOM[10'h190][30];	// lsu.scala:211:16
        stq_7_bits_uop_iw_p2_poisoned = _RANDOM[10'h190][31];	// lsu.scala:211:16
        stq_7_bits_uop_is_br = _RANDOM[10'h191][0];	// lsu.scala:211:16
        stq_7_bits_uop_is_jalr = _RANDOM[10'h191][1];	// lsu.scala:211:16
        stq_7_bits_uop_is_jal = _RANDOM[10'h191][2];	// lsu.scala:211:16
        stq_7_bits_uop_is_sfb = _RANDOM[10'h191][3];	// lsu.scala:211:16
        stq_7_bits_uop_br_mask = _RANDOM[10'h191][15:4];	// lsu.scala:211:16
        stq_7_bits_uop_br_tag = _RANDOM[10'h191][19:16];	// lsu.scala:211:16
        stq_7_bits_uop_ftq_idx = _RANDOM[10'h191][24:20];	// lsu.scala:211:16
        stq_7_bits_uop_edge_inst = _RANDOM[10'h191][25];	// lsu.scala:211:16
        stq_7_bits_uop_pc_lob = _RANDOM[10'h191][31:26];	// lsu.scala:211:16
        stq_7_bits_uop_taken = _RANDOM[10'h192][0];	// lsu.scala:211:16
        stq_7_bits_uop_imm_packed = _RANDOM[10'h192][20:1];	// lsu.scala:211:16
        stq_7_bits_uop_csr_addr = {_RANDOM[10'h192][31:21], _RANDOM[10'h193][0]};	// lsu.scala:211:16
        stq_7_bits_uop_rob_idx = _RANDOM[10'h193][6:1];	// lsu.scala:211:16
        stq_7_bits_uop_ldq_idx = _RANDOM[10'h193][10:7];	// lsu.scala:211:16
        stq_7_bits_uop_stq_idx = _RANDOM[10'h193][14:11];	// lsu.scala:211:16
        stq_7_bits_uop_rxq_idx = _RANDOM[10'h193][16:15];	// lsu.scala:211:16
        stq_7_bits_uop_pdst = _RANDOM[10'h193][23:17];	// lsu.scala:211:16
        stq_7_bits_uop_prs1 = _RANDOM[10'h193][30:24];	// lsu.scala:211:16
        stq_7_bits_uop_prs2 = {_RANDOM[10'h193][31], _RANDOM[10'h194][5:0]};	// lsu.scala:211:16
        stq_7_bits_uop_prs3 = _RANDOM[10'h194][12:6];	// lsu.scala:211:16
        stq_7_bits_uop_ppred = _RANDOM[10'h194][17:13];	// lsu.scala:211:16
        stq_7_bits_uop_prs1_busy = _RANDOM[10'h194][18];	// lsu.scala:211:16
        stq_7_bits_uop_prs2_busy = _RANDOM[10'h194][19];	// lsu.scala:211:16
        stq_7_bits_uop_prs3_busy = _RANDOM[10'h194][20];	// lsu.scala:211:16
        stq_7_bits_uop_ppred_busy = _RANDOM[10'h194][21];	// lsu.scala:211:16
        stq_7_bits_uop_stale_pdst = _RANDOM[10'h194][28:22];	// lsu.scala:211:16
        stq_7_bits_uop_exception = _RANDOM[10'h194][29];	// lsu.scala:211:16
        stq_7_bits_uop_exc_cause =
          {_RANDOM[10'h194][31:30], _RANDOM[10'h195], _RANDOM[10'h196][29:0]};	// lsu.scala:211:16
        stq_7_bits_uop_bypassable = _RANDOM[10'h196][30];	// lsu.scala:211:16
        stq_7_bits_uop_mem_cmd = {_RANDOM[10'h196][31], _RANDOM[10'h197][3:0]};	// lsu.scala:211:16
        stq_7_bits_uop_mem_size = _RANDOM[10'h197][5:4];	// lsu.scala:211:16
        stq_7_bits_uop_mem_signed = _RANDOM[10'h197][6];	// lsu.scala:211:16
        stq_7_bits_uop_is_fence = _RANDOM[10'h197][7];	// lsu.scala:211:16
        stq_7_bits_uop_is_fencei = _RANDOM[10'h197][8];	// lsu.scala:211:16
        stq_7_bits_uop_is_amo = _RANDOM[10'h197][9];	// lsu.scala:211:16
        stq_7_bits_uop_uses_ldq = _RANDOM[10'h197][10];	// lsu.scala:211:16
        stq_7_bits_uop_uses_stq = _RANDOM[10'h197][11];	// lsu.scala:211:16
        stq_7_bits_uop_is_sys_pc2epc = _RANDOM[10'h197][12];	// lsu.scala:211:16
        stq_7_bits_uop_is_unique = _RANDOM[10'h197][13];	// lsu.scala:211:16
        stq_7_bits_uop_flush_on_commit = _RANDOM[10'h197][14];	// lsu.scala:211:16
        stq_7_bits_uop_ldst_is_rs1 = _RANDOM[10'h197][15];	// lsu.scala:211:16
        stq_7_bits_uop_ldst = _RANDOM[10'h197][21:16];	// lsu.scala:211:16
        stq_7_bits_uop_lrs1 = _RANDOM[10'h197][27:22];	// lsu.scala:211:16
        stq_7_bits_uop_lrs2 = {_RANDOM[10'h197][31:28], _RANDOM[10'h198][1:0]};	// lsu.scala:211:16
        stq_7_bits_uop_lrs3 = _RANDOM[10'h198][7:2];	// lsu.scala:211:16
        stq_7_bits_uop_ldst_val = _RANDOM[10'h198][8];	// lsu.scala:211:16
        stq_7_bits_uop_dst_rtype = _RANDOM[10'h198][10:9];	// lsu.scala:211:16
        stq_7_bits_uop_lrs1_rtype = _RANDOM[10'h198][12:11];	// lsu.scala:211:16
        stq_7_bits_uop_lrs2_rtype = _RANDOM[10'h198][14:13];	// lsu.scala:211:16
        stq_7_bits_uop_frs3_en = _RANDOM[10'h198][15];	// lsu.scala:211:16
        stq_7_bits_uop_fp_val = _RANDOM[10'h198][16];	// lsu.scala:211:16
        stq_7_bits_uop_fp_single = _RANDOM[10'h198][17];	// lsu.scala:211:16
        stq_7_bits_uop_xcpt_pf_if = _RANDOM[10'h198][18];	// lsu.scala:211:16
        stq_7_bits_uop_xcpt_ae_if = _RANDOM[10'h198][19];	// lsu.scala:211:16
        stq_7_bits_uop_xcpt_ma_if = _RANDOM[10'h198][20];	// lsu.scala:211:16
        stq_7_bits_uop_bp_debug_if = _RANDOM[10'h198][21];	// lsu.scala:211:16
        stq_7_bits_uop_bp_xcpt_if = _RANDOM[10'h198][22];	// lsu.scala:211:16
        stq_7_bits_uop_debug_fsrc = _RANDOM[10'h198][24:23];	// lsu.scala:211:16
        stq_7_bits_uop_debug_tsrc = _RANDOM[10'h198][26:25];	// lsu.scala:211:16
        stq_7_bits_addr_valid = _RANDOM[10'h198][27];	// lsu.scala:211:16
        stq_7_bits_addr_bits =
          {_RANDOM[10'h198][31:28], _RANDOM[10'h199], _RANDOM[10'h19A][3:0]};	// lsu.scala:211:16
        stq_7_bits_addr_is_virtual = _RANDOM[10'h19A][4];	// lsu.scala:211:16
        stq_7_bits_data_valid = _RANDOM[10'h19A][5];	// lsu.scala:211:16
        stq_7_bits_data_bits =
          {_RANDOM[10'h19A][31:6], _RANDOM[10'h19B], _RANDOM[10'h19C][5:0]};	// lsu.scala:211:16
        stq_7_bits_committed = _RANDOM[10'h19C][6];	// lsu.scala:211:16
        stq_7_bits_succeeded = _RANDOM[10'h19C][7];	// lsu.scala:211:16
        stq_8_valid = _RANDOM[10'h19E][8];	// lsu.scala:211:16
        stq_8_bits_uop_uopc = _RANDOM[10'h19E][15:9];	// lsu.scala:211:16
        stq_8_bits_uop_inst = {_RANDOM[10'h19E][31:16], _RANDOM[10'h19F][15:0]};	// lsu.scala:211:16
        stq_8_bits_uop_debug_inst = {_RANDOM[10'h19F][31:16], _RANDOM[10'h1A0][15:0]};	// lsu.scala:211:16
        stq_8_bits_uop_is_rvc = _RANDOM[10'h1A0][16];	// lsu.scala:211:16
        stq_8_bits_uop_debug_pc = {_RANDOM[10'h1A0][31:17], _RANDOM[10'h1A1][24:0]};	// lsu.scala:211:16
        stq_8_bits_uop_iq_type = _RANDOM[10'h1A1][27:25];	// lsu.scala:211:16
        stq_8_bits_uop_fu_code = {_RANDOM[10'h1A1][31:28], _RANDOM[10'h1A2][5:0]};	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_br_type = _RANDOM[10'h1A2][9:6];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op1_sel = _RANDOM[10'h1A2][11:10];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op2_sel = _RANDOM[10'h1A2][14:12];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_imm_sel = _RANDOM[10'h1A2][17:15];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_op_fcn = _RANDOM[10'h1A2][21:18];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1A2][22];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1A2][25:23];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_is_load = _RANDOM[10'h1A2][26];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_is_sta = _RANDOM[10'h1A2][27];	// lsu.scala:211:16
        stq_8_bits_uop_ctrl_is_std = _RANDOM[10'h1A2][28];	// lsu.scala:211:16
        stq_8_bits_uop_iw_state = _RANDOM[10'h1A2][30:29];	// lsu.scala:211:16
        stq_8_bits_uop_iw_p1_poisoned = _RANDOM[10'h1A2][31];	// lsu.scala:211:16
        stq_8_bits_uop_iw_p2_poisoned = _RANDOM[10'h1A3][0];	// lsu.scala:211:16
        stq_8_bits_uop_is_br = _RANDOM[10'h1A3][1];	// lsu.scala:211:16
        stq_8_bits_uop_is_jalr = _RANDOM[10'h1A3][2];	// lsu.scala:211:16
        stq_8_bits_uop_is_jal = _RANDOM[10'h1A3][3];	// lsu.scala:211:16
        stq_8_bits_uop_is_sfb = _RANDOM[10'h1A3][4];	// lsu.scala:211:16
        stq_8_bits_uop_br_mask = _RANDOM[10'h1A3][16:5];	// lsu.scala:211:16
        stq_8_bits_uop_br_tag = _RANDOM[10'h1A3][20:17];	// lsu.scala:211:16
        stq_8_bits_uop_ftq_idx = _RANDOM[10'h1A3][25:21];	// lsu.scala:211:16
        stq_8_bits_uop_edge_inst = _RANDOM[10'h1A3][26];	// lsu.scala:211:16
        stq_8_bits_uop_pc_lob = {_RANDOM[10'h1A3][31:27], _RANDOM[10'h1A4][0]};	// lsu.scala:211:16
        stq_8_bits_uop_taken = _RANDOM[10'h1A4][1];	// lsu.scala:211:16
        stq_8_bits_uop_imm_packed = _RANDOM[10'h1A4][21:2];	// lsu.scala:211:16
        stq_8_bits_uop_csr_addr = {_RANDOM[10'h1A4][31:22], _RANDOM[10'h1A5][1:0]};	// lsu.scala:211:16
        stq_8_bits_uop_rob_idx = _RANDOM[10'h1A5][7:2];	// lsu.scala:211:16
        stq_8_bits_uop_ldq_idx = _RANDOM[10'h1A5][11:8];	// lsu.scala:211:16
        stq_8_bits_uop_stq_idx = _RANDOM[10'h1A5][15:12];	// lsu.scala:211:16
        stq_8_bits_uop_rxq_idx = _RANDOM[10'h1A5][17:16];	// lsu.scala:211:16
        stq_8_bits_uop_pdst = _RANDOM[10'h1A5][24:18];	// lsu.scala:211:16
        stq_8_bits_uop_prs1 = _RANDOM[10'h1A5][31:25];	// lsu.scala:211:16
        stq_8_bits_uop_prs2 = _RANDOM[10'h1A6][6:0];	// lsu.scala:211:16
        stq_8_bits_uop_prs3 = _RANDOM[10'h1A6][13:7];	// lsu.scala:211:16
        stq_8_bits_uop_ppred = _RANDOM[10'h1A6][18:14];	// lsu.scala:211:16
        stq_8_bits_uop_prs1_busy = _RANDOM[10'h1A6][19];	// lsu.scala:211:16
        stq_8_bits_uop_prs2_busy = _RANDOM[10'h1A6][20];	// lsu.scala:211:16
        stq_8_bits_uop_prs3_busy = _RANDOM[10'h1A6][21];	// lsu.scala:211:16
        stq_8_bits_uop_ppred_busy = _RANDOM[10'h1A6][22];	// lsu.scala:211:16
        stq_8_bits_uop_stale_pdst = _RANDOM[10'h1A6][29:23];	// lsu.scala:211:16
        stq_8_bits_uop_exception = _RANDOM[10'h1A6][30];	// lsu.scala:211:16
        stq_8_bits_uop_exc_cause =
          {_RANDOM[10'h1A6][31], _RANDOM[10'h1A7], _RANDOM[10'h1A8][30:0]};	// lsu.scala:211:16
        stq_8_bits_uop_bypassable = _RANDOM[10'h1A8][31];	// lsu.scala:211:16
        stq_8_bits_uop_mem_cmd = _RANDOM[10'h1A9][4:0];	// lsu.scala:211:16
        stq_8_bits_uop_mem_size = _RANDOM[10'h1A9][6:5];	// lsu.scala:211:16
        stq_8_bits_uop_mem_signed = _RANDOM[10'h1A9][7];	// lsu.scala:211:16
        stq_8_bits_uop_is_fence = _RANDOM[10'h1A9][8];	// lsu.scala:211:16
        stq_8_bits_uop_is_fencei = _RANDOM[10'h1A9][9];	// lsu.scala:211:16
        stq_8_bits_uop_is_amo = _RANDOM[10'h1A9][10];	// lsu.scala:211:16
        stq_8_bits_uop_uses_ldq = _RANDOM[10'h1A9][11];	// lsu.scala:211:16
        stq_8_bits_uop_uses_stq = _RANDOM[10'h1A9][12];	// lsu.scala:211:16
        stq_8_bits_uop_is_sys_pc2epc = _RANDOM[10'h1A9][13];	// lsu.scala:211:16
        stq_8_bits_uop_is_unique = _RANDOM[10'h1A9][14];	// lsu.scala:211:16
        stq_8_bits_uop_flush_on_commit = _RANDOM[10'h1A9][15];	// lsu.scala:211:16
        stq_8_bits_uop_ldst_is_rs1 = _RANDOM[10'h1A9][16];	// lsu.scala:211:16
        stq_8_bits_uop_ldst = _RANDOM[10'h1A9][22:17];	// lsu.scala:211:16
        stq_8_bits_uop_lrs1 = _RANDOM[10'h1A9][28:23];	// lsu.scala:211:16
        stq_8_bits_uop_lrs2 = {_RANDOM[10'h1A9][31:29], _RANDOM[10'h1AA][2:0]};	// lsu.scala:211:16
        stq_8_bits_uop_lrs3 = _RANDOM[10'h1AA][8:3];	// lsu.scala:211:16
        stq_8_bits_uop_ldst_val = _RANDOM[10'h1AA][9];	// lsu.scala:211:16
        stq_8_bits_uop_dst_rtype = _RANDOM[10'h1AA][11:10];	// lsu.scala:211:16
        stq_8_bits_uop_lrs1_rtype = _RANDOM[10'h1AA][13:12];	// lsu.scala:211:16
        stq_8_bits_uop_lrs2_rtype = _RANDOM[10'h1AA][15:14];	// lsu.scala:211:16
        stq_8_bits_uop_frs3_en = _RANDOM[10'h1AA][16];	// lsu.scala:211:16
        stq_8_bits_uop_fp_val = _RANDOM[10'h1AA][17];	// lsu.scala:211:16
        stq_8_bits_uop_fp_single = _RANDOM[10'h1AA][18];	// lsu.scala:211:16
        stq_8_bits_uop_xcpt_pf_if = _RANDOM[10'h1AA][19];	// lsu.scala:211:16
        stq_8_bits_uop_xcpt_ae_if = _RANDOM[10'h1AA][20];	// lsu.scala:211:16
        stq_8_bits_uop_xcpt_ma_if = _RANDOM[10'h1AA][21];	// lsu.scala:211:16
        stq_8_bits_uop_bp_debug_if = _RANDOM[10'h1AA][22];	// lsu.scala:211:16
        stq_8_bits_uop_bp_xcpt_if = _RANDOM[10'h1AA][23];	// lsu.scala:211:16
        stq_8_bits_uop_debug_fsrc = _RANDOM[10'h1AA][25:24];	// lsu.scala:211:16
        stq_8_bits_uop_debug_tsrc = _RANDOM[10'h1AA][27:26];	// lsu.scala:211:16
        stq_8_bits_addr_valid = _RANDOM[10'h1AA][28];	// lsu.scala:211:16
        stq_8_bits_addr_bits =
          {_RANDOM[10'h1AA][31:29], _RANDOM[10'h1AB], _RANDOM[10'h1AC][4:0]};	// lsu.scala:211:16
        stq_8_bits_addr_is_virtual = _RANDOM[10'h1AC][5];	// lsu.scala:211:16
        stq_8_bits_data_valid = _RANDOM[10'h1AC][6];	// lsu.scala:211:16
        stq_8_bits_data_bits =
          {_RANDOM[10'h1AC][31:7], _RANDOM[10'h1AD], _RANDOM[10'h1AE][6:0]};	// lsu.scala:211:16
        stq_8_bits_committed = _RANDOM[10'h1AE][7];	// lsu.scala:211:16
        stq_8_bits_succeeded = _RANDOM[10'h1AE][8];	// lsu.scala:211:16
        stq_9_valid = _RANDOM[10'h1B0][9];	// lsu.scala:211:16
        stq_9_bits_uop_uopc = _RANDOM[10'h1B0][16:10];	// lsu.scala:211:16
        stq_9_bits_uop_inst = {_RANDOM[10'h1B0][31:17], _RANDOM[10'h1B1][16:0]};	// lsu.scala:211:16
        stq_9_bits_uop_debug_inst = {_RANDOM[10'h1B1][31:17], _RANDOM[10'h1B2][16:0]};	// lsu.scala:211:16
        stq_9_bits_uop_is_rvc = _RANDOM[10'h1B2][17];	// lsu.scala:211:16
        stq_9_bits_uop_debug_pc = {_RANDOM[10'h1B2][31:18], _RANDOM[10'h1B3][25:0]};	// lsu.scala:211:16
        stq_9_bits_uop_iq_type = _RANDOM[10'h1B3][28:26];	// lsu.scala:211:16
        stq_9_bits_uop_fu_code = {_RANDOM[10'h1B3][31:29], _RANDOM[10'h1B4][6:0]};	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_br_type = _RANDOM[10'h1B4][10:7];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op1_sel = _RANDOM[10'h1B4][12:11];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op2_sel = _RANDOM[10'h1B4][15:13];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_imm_sel = _RANDOM[10'h1B4][18:16];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_op_fcn = _RANDOM[10'h1B4][22:19];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1B4][23];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1B4][26:24];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_is_load = _RANDOM[10'h1B4][27];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_is_sta = _RANDOM[10'h1B4][28];	// lsu.scala:211:16
        stq_9_bits_uop_ctrl_is_std = _RANDOM[10'h1B4][29];	// lsu.scala:211:16
        stq_9_bits_uop_iw_state = _RANDOM[10'h1B4][31:30];	// lsu.scala:211:16
        stq_9_bits_uop_iw_p1_poisoned = _RANDOM[10'h1B5][0];	// lsu.scala:211:16
        stq_9_bits_uop_iw_p2_poisoned = _RANDOM[10'h1B5][1];	// lsu.scala:211:16
        stq_9_bits_uop_is_br = _RANDOM[10'h1B5][2];	// lsu.scala:211:16
        stq_9_bits_uop_is_jalr = _RANDOM[10'h1B5][3];	// lsu.scala:211:16
        stq_9_bits_uop_is_jal = _RANDOM[10'h1B5][4];	// lsu.scala:211:16
        stq_9_bits_uop_is_sfb = _RANDOM[10'h1B5][5];	// lsu.scala:211:16
        stq_9_bits_uop_br_mask = _RANDOM[10'h1B5][17:6];	// lsu.scala:211:16
        stq_9_bits_uop_br_tag = _RANDOM[10'h1B5][21:18];	// lsu.scala:211:16
        stq_9_bits_uop_ftq_idx = _RANDOM[10'h1B5][26:22];	// lsu.scala:211:16
        stq_9_bits_uop_edge_inst = _RANDOM[10'h1B5][27];	// lsu.scala:211:16
        stq_9_bits_uop_pc_lob = {_RANDOM[10'h1B5][31:28], _RANDOM[10'h1B6][1:0]};	// lsu.scala:211:16
        stq_9_bits_uop_taken = _RANDOM[10'h1B6][2];	// lsu.scala:211:16
        stq_9_bits_uop_imm_packed = _RANDOM[10'h1B6][22:3];	// lsu.scala:211:16
        stq_9_bits_uop_csr_addr = {_RANDOM[10'h1B6][31:23], _RANDOM[10'h1B7][2:0]};	// lsu.scala:211:16
        stq_9_bits_uop_rob_idx = _RANDOM[10'h1B7][8:3];	// lsu.scala:211:16
        stq_9_bits_uop_ldq_idx = _RANDOM[10'h1B7][12:9];	// lsu.scala:211:16
        stq_9_bits_uop_stq_idx = _RANDOM[10'h1B7][16:13];	// lsu.scala:211:16
        stq_9_bits_uop_rxq_idx = _RANDOM[10'h1B7][18:17];	// lsu.scala:211:16
        stq_9_bits_uop_pdst = _RANDOM[10'h1B7][25:19];	// lsu.scala:211:16
        stq_9_bits_uop_prs1 = {_RANDOM[10'h1B7][31:26], _RANDOM[10'h1B8][0]};	// lsu.scala:211:16
        stq_9_bits_uop_prs2 = _RANDOM[10'h1B8][7:1];	// lsu.scala:211:16
        stq_9_bits_uop_prs3 = _RANDOM[10'h1B8][14:8];	// lsu.scala:211:16
        stq_9_bits_uop_ppred = _RANDOM[10'h1B8][19:15];	// lsu.scala:211:16
        stq_9_bits_uop_prs1_busy = _RANDOM[10'h1B8][20];	// lsu.scala:211:16
        stq_9_bits_uop_prs2_busy = _RANDOM[10'h1B8][21];	// lsu.scala:211:16
        stq_9_bits_uop_prs3_busy = _RANDOM[10'h1B8][22];	// lsu.scala:211:16
        stq_9_bits_uop_ppred_busy = _RANDOM[10'h1B8][23];	// lsu.scala:211:16
        stq_9_bits_uop_stale_pdst = _RANDOM[10'h1B8][30:24];	// lsu.scala:211:16
        stq_9_bits_uop_exception = _RANDOM[10'h1B8][31];	// lsu.scala:211:16
        stq_9_bits_uop_exc_cause = {_RANDOM[10'h1B9], _RANDOM[10'h1BA]};	// lsu.scala:211:16
        stq_9_bits_uop_bypassable = _RANDOM[10'h1BB][0];	// lsu.scala:211:16
        stq_9_bits_uop_mem_cmd = _RANDOM[10'h1BB][5:1];	// lsu.scala:211:16
        stq_9_bits_uop_mem_size = _RANDOM[10'h1BB][7:6];	// lsu.scala:211:16
        stq_9_bits_uop_mem_signed = _RANDOM[10'h1BB][8];	// lsu.scala:211:16
        stq_9_bits_uop_is_fence = _RANDOM[10'h1BB][9];	// lsu.scala:211:16
        stq_9_bits_uop_is_fencei = _RANDOM[10'h1BB][10];	// lsu.scala:211:16
        stq_9_bits_uop_is_amo = _RANDOM[10'h1BB][11];	// lsu.scala:211:16
        stq_9_bits_uop_uses_ldq = _RANDOM[10'h1BB][12];	// lsu.scala:211:16
        stq_9_bits_uop_uses_stq = _RANDOM[10'h1BB][13];	// lsu.scala:211:16
        stq_9_bits_uop_is_sys_pc2epc = _RANDOM[10'h1BB][14];	// lsu.scala:211:16
        stq_9_bits_uop_is_unique = _RANDOM[10'h1BB][15];	// lsu.scala:211:16
        stq_9_bits_uop_flush_on_commit = _RANDOM[10'h1BB][16];	// lsu.scala:211:16
        stq_9_bits_uop_ldst_is_rs1 = _RANDOM[10'h1BB][17];	// lsu.scala:211:16
        stq_9_bits_uop_ldst = _RANDOM[10'h1BB][23:18];	// lsu.scala:211:16
        stq_9_bits_uop_lrs1 = _RANDOM[10'h1BB][29:24];	// lsu.scala:211:16
        stq_9_bits_uop_lrs2 = {_RANDOM[10'h1BB][31:30], _RANDOM[10'h1BC][3:0]};	// lsu.scala:211:16
        stq_9_bits_uop_lrs3 = _RANDOM[10'h1BC][9:4];	// lsu.scala:211:16
        stq_9_bits_uop_ldst_val = _RANDOM[10'h1BC][10];	// lsu.scala:211:16
        stq_9_bits_uop_dst_rtype = _RANDOM[10'h1BC][12:11];	// lsu.scala:211:16
        stq_9_bits_uop_lrs1_rtype = _RANDOM[10'h1BC][14:13];	// lsu.scala:211:16
        stq_9_bits_uop_lrs2_rtype = _RANDOM[10'h1BC][16:15];	// lsu.scala:211:16
        stq_9_bits_uop_frs3_en = _RANDOM[10'h1BC][17];	// lsu.scala:211:16
        stq_9_bits_uop_fp_val = _RANDOM[10'h1BC][18];	// lsu.scala:211:16
        stq_9_bits_uop_fp_single = _RANDOM[10'h1BC][19];	// lsu.scala:211:16
        stq_9_bits_uop_xcpt_pf_if = _RANDOM[10'h1BC][20];	// lsu.scala:211:16
        stq_9_bits_uop_xcpt_ae_if = _RANDOM[10'h1BC][21];	// lsu.scala:211:16
        stq_9_bits_uop_xcpt_ma_if = _RANDOM[10'h1BC][22];	// lsu.scala:211:16
        stq_9_bits_uop_bp_debug_if = _RANDOM[10'h1BC][23];	// lsu.scala:211:16
        stq_9_bits_uop_bp_xcpt_if = _RANDOM[10'h1BC][24];	// lsu.scala:211:16
        stq_9_bits_uop_debug_fsrc = _RANDOM[10'h1BC][26:25];	// lsu.scala:211:16
        stq_9_bits_uop_debug_tsrc = _RANDOM[10'h1BC][28:27];	// lsu.scala:211:16
        stq_9_bits_addr_valid = _RANDOM[10'h1BC][29];	// lsu.scala:211:16
        stq_9_bits_addr_bits =
          {_RANDOM[10'h1BC][31:30], _RANDOM[10'h1BD], _RANDOM[10'h1BE][5:0]};	// lsu.scala:211:16
        stq_9_bits_addr_is_virtual = _RANDOM[10'h1BE][6];	// lsu.scala:211:16
        stq_9_bits_data_valid = _RANDOM[10'h1BE][7];	// lsu.scala:211:16
        stq_9_bits_data_bits =
          {_RANDOM[10'h1BE][31:8], _RANDOM[10'h1BF], _RANDOM[10'h1C0][7:0]};	// lsu.scala:211:16
        stq_9_bits_committed = _RANDOM[10'h1C0][8];	// lsu.scala:211:16
        stq_9_bits_succeeded = _RANDOM[10'h1C0][9];	// lsu.scala:211:16
        stq_10_valid = _RANDOM[10'h1C2][10];	// lsu.scala:211:16
        stq_10_bits_uop_uopc = _RANDOM[10'h1C2][17:11];	// lsu.scala:211:16
        stq_10_bits_uop_inst = {_RANDOM[10'h1C2][31:18], _RANDOM[10'h1C3][17:0]};	// lsu.scala:211:16
        stq_10_bits_uop_debug_inst = {_RANDOM[10'h1C3][31:18], _RANDOM[10'h1C4][17:0]};	// lsu.scala:211:16
        stq_10_bits_uop_is_rvc = _RANDOM[10'h1C4][18];	// lsu.scala:211:16
        stq_10_bits_uop_debug_pc = {_RANDOM[10'h1C4][31:19], _RANDOM[10'h1C5][26:0]};	// lsu.scala:211:16
        stq_10_bits_uop_iq_type = _RANDOM[10'h1C5][29:27];	// lsu.scala:211:16
        stq_10_bits_uop_fu_code = {_RANDOM[10'h1C5][31:30], _RANDOM[10'h1C6][7:0]};	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_br_type = _RANDOM[10'h1C6][11:8];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op1_sel = _RANDOM[10'h1C6][13:12];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op2_sel = _RANDOM[10'h1C6][16:14];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_imm_sel = _RANDOM[10'h1C6][19:17];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_op_fcn = _RANDOM[10'h1C6][23:20];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1C6][24];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1C6][27:25];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_is_load = _RANDOM[10'h1C6][28];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_is_sta = _RANDOM[10'h1C6][29];	// lsu.scala:211:16
        stq_10_bits_uop_ctrl_is_std = _RANDOM[10'h1C6][30];	// lsu.scala:211:16
        stq_10_bits_uop_iw_state = {_RANDOM[10'h1C6][31], _RANDOM[10'h1C7][0]};	// lsu.scala:211:16
        stq_10_bits_uop_iw_p1_poisoned = _RANDOM[10'h1C7][1];	// lsu.scala:211:16
        stq_10_bits_uop_iw_p2_poisoned = _RANDOM[10'h1C7][2];	// lsu.scala:211:16
        stq_10_bits_uop_is_br = _RANDOM[10'h1C7][3];	// lsu.scala:211:16
        stq_10_bits_uop_is_jalr = _RANDOM[10'h1C7][4];	// lsu.scala:211:16
        stq_10_bits_uop_is_jal = _RANDOM[10'h1C7][5];	// lsu.scala:211:16
        stq_10_bits_uop_is_sfb = _RANDOM[10'h1C7][6];	// lsu.scala:211:16
        stq_10_bits_uop_br_mask = _RANDOM[10'h1C7][18:7];	// lsu.scala:211:16
        stq_10_bits_uop_br_tag = _RANDOM[10'h1C7][22:19];	// lsu.scala:211:16
        stq_10_bits_uop_ftq_idx = _RANDOM[10'h1C7][27:23];	// lsu.scala:211:16
        stq_10_bits_uop_edge_inst = _RANDOM[10'h1C7][28];	// lsu.scala:211:16
        stq_10_bits_uop_pc_lob = {_RANDOM[10'h1C7][31:29], _RANDOM[10'h1C8][2:0]};	// lsu.scala:211:16
        stq_10_bits_uop_taken = _RANDOM[10'h1C8][3];	// lsu.scala:211:16
        stq_10_bits_uop_imm_packed = _RANDOM[10'h1C8][23:4];	// lsu.scala:211:16
        stq_10_bits_uop_csr_addr = {_RANDOM[10'h1C8][31:24], _RANDOM[10'h1C9][3:0]};	// lsu.scala:211:16
        stq_10_bits_uop_rob_idx = _RANDOM[10'h1C9][9:4];	// lsu.scala:211:16
        stq_10_bits_uop_ldq_idx = _RANDOM[10'h1C9][13:10];	// lsu.scala:211:16
        stq_10_bits_uop_stq_idx = _RANDOM[10'h1C9][17:14];	// lsu.scala:211:16
        stq_10_bits_uop_rxq_idx = _RANDOM[10'h1C9][19:18];	// lsu.scala:211:16
        stq_10_bits_uop_pdst = _RANDOM[10'h1C9][26:20];	// lsu.scala:211:16
        stq_10_bits_uop_prs1 = {_RANDOM[10'h1C9][31:27], _RANDOM[10'h1CA][1:0]};	// lsu.scala:211:16
        stq_10_bits_uop_prs2 = _RANDOM[10'h1CA][8:2];	// lsu.scala:211:16
        stq_10_bits_uop_prs3 = _RANDOM[10'h1CA][15:9];	// lsu.scala:211:16
        stq_10_bits_uop_ppred = _RANDOM[10'h1CA][20:16];	// lsu.scala:211:16
        stq_10_bits_uop_prs1_busy = _RANDOM[10'h1CA][21];	// lsu.scala:211:16
        stq_10_bits_uop_prs2_busy = _RANDOM[10'h1CA][22];	// lsu.scala:211:16
        stq_10_bits_uop_prs3_busy = _RANDOM[10'h1CA][23];	// lsu.scala:211:16
        stq_10_bits_uop_ppred_busy = _RANDOM[10'h1CA][24];	// lsu.scala:211:16
        stq_10_bits_uop_stale_pdst = _RANDOM[10'h1CA][31:25];	// lsu.scala:211:16
        stq_10_bits_uop_exception = _RANDOM[10'h1CB][0];	// lsu.scala:211:16
        stq_10_bits_uop_exc_cause =
          {_RANDOM[10'h1CB][31:1], _RANDOM[10'h1CC], _RANDOM[10'h1CD][0]};	// lsu.scala:211:16
        stq_10_bits_uop_bypassable = _RANDOM[10'h1CD][1];	// lsu.scala:211:16
        stq_10_bits_uop_mem_cmd = _RANDOM[10'h1CD][6:2];	// lsu.scala:211:16
        stq_10_bits_uop_mem_size = _RANDOM[10'h1CD][8:7];	// lsu.scala:211:16
        stq_10_bits_uop_mem_signed = _RANDOM[10'h1CD][9];	// lsu.scala:211:16
        stq_10_bits_uop_is_fence = _RANDOM[10'h1CD][10];	// lsu.scala:211:16
        stq_10_bits_uop_is_fencei = _RANDOM[10'h1CD][11];	// lsu.scala:211:16
        stq_10_bits_uop_is_amo = _RANDOM[10'h1CD][12];	// lsu.scala:211:16
        stq_10_bits_uop_uses_ldq = _RANDOM[10'h1CD][13];	// lsu.scala:211:16
        stq_10_bits_uop_uses_stq = _RANDOM[10'h1CD][14];	// lsu.scala:211:16
        stq_10_bits_uop_is_sys_pc2epc = _RANDOM[10'h1CD][15];	// lsu.scala:211:16
        stq_10_bits_uop_is_unique = _RANDOM[10'h1CD][16];	// lsu.scala:211:16
        stq_10_bits_uop_flush_on_commit = _RANDOM[10'h1CD][17];	// lsu.scala:211:16
        stq_10_bits_uop_ldst_is_rs1 = _RANDOM[10'h1CD][18];	// lsu.scala:211:16
        stq_10_bits_uop_ldst = _RANDOM[10'h1CD][24:19];	// lsu.scala:211:16
        stq_10_bits_uop_lrs1 = _RANDOM[10'h1CD][30:25];	// lsu.scala:211:16
        stq_10_bits_uop_lrs2 = {_RANDOM[10'h1CD][31], _RANDOM[10'h1CE][4:0]};	// lsu.scala:211:16
        stq_10_bits_uop_lrs3 = _RANDOM[10'h1CE][10:5];	// lsu.scala:211:16
        stq_10_bits_uop_ldst_val = _RANDOM[10'h1CE][11];	// lsu.scala:211:16
        stq_10_bits_uop_dst_rtype = _RANDOM[10'h1CE][13:12];	// lsu.scala:211:16
        stq_10_bits_uop_lrs1_rtype = _RANDOM[10'h1CE][15:14];	// lsu.scala:211:16
        stq_10_bits_uop_lrs2_rtype = _RANDOM[10'h1CE][17:16];	// lsu.scala:211:16
        stq_10_bits_uop_frs3_en = _RANDOM[10'h1CE][18];	// lsu.scala:211:16
        stq_10_bits_uop_fp_val = _RANDOM[10'h1CE][19];	// lsu.scala:211:16
        stq_10_bits_uop_fp_single = _RANDOM[10'h1CE][20];	// lsu.scala:211:16
        stq_10_bits_uop_xcpt_pf_if = _RANDOM[10'h1CE][21];	// lsu.scala:211:16
        stq_10_bits_uop_xcpt_ae_if = _RANDOM[10'h1CE][22];	// lsu.scala:211:16
        stq_10_bits_uop_xcpt_ma_if = _RANDOM[10'h1CE][23];	// lsu.scala:211:16
        stq_10_bits_uop_bp_debug_if = _RANDOM[10'h1CE][24];	// lsu.scala:211:16
        stq_10_bits_uop_bp_xcpt_if = _RANDOM[10'h1CE][25];	// lsu.scala:211:16
        stq_10_bits_uop_debug_fsrc = _RANDOM[10'h1CE][27:26];	// lsu.scala:211:16
        stq_10_bits_uop_debug_tsrc = _RANDOM[10'h1CE][29:28];	// lsu.scala:211:16
        stq_10_bits_addr_valid = _RANDOM[10'h1CE][30];	// lsu.scala:211:16
        stq_10_bits_addr_bits =
          {_RANDOM[10'h1CE][31], _RANDOM[10'h1CF], _RANDOM[10'h1D0][6:0]};	// lsu.scala:211:16
        stq_10_bits_addr_is_virtual = _RANDOM[10'h1D0][7];	// lsu.scala:211:16
        stq_10_bits_data_valid = _RANDOM[10'h1D0][8];	// lsu.scala:211:16
        stq_10_bits_data_bits =
          {_RANDOM[10'h1D0][31:9], _RANDOM[10'h1D1], _RANDOM[10'h1D2][8:0]};	// lsu.scala:211:16
        stq_10_bits_committed = _RANDOM[10'h1D2][9];	// lsu.scala:211:16
        stq_10_bits_succeeded = _RANDOM[10'h1D2][10];	// lsu.scala:211:16
        stq_11_valid = _RANDOM[10'h1D4][11];	// lsu.scala:211:16
        stq_11_bits_uop_uopc = _RANDOM[10'h1D4][18:12];	// lsu.scala:211:16
        stq_11_bits_uop_inst = {_RANDOM[10'h1D4][31:19], _RANDOM[10'h1D5][18:0]};	// lsu.scala:211:16
        stq_11_bits_uop_debug_inst = {_RANDOM[10'h1D5][31:19], _RANDOM[10'h1D6][18:0]};	// lsu.scala:211:16
        stq_11_bits_uop_is_rvc = _RANDOM[10'h1D6][19];	// lsu.scala:211:16
        stq_11_bits_uop_debug_pc = {_RANDOM[10'h1D6][31:20], _RANDOM[10'h1D7][27:0]};	// lsu.scala:211:16
        stq_11_bits_uop_iq_type = _RANDOM[10'h1D7][30:28];	// lsu.scala:211:16
        stq_11_bits_uop_fu_code = {_RANDOM[10'h1D7][31], _RANDOM[10'h1D8][8:0]};	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_br_type = _RANDOM[10'h1D8][12:9];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op1_sel = _RANDOM[10'h1D8][14:13];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op2_sel = _RANDOM[10'h1D8][17:15];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_imm_sel = _RANDOM[10'h1D8][20:18];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_op_fcn = _RANDOM[10'h1D8][24:21];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1D8][25];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1D8][28:26];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_is_load = _RANDOM[10'h1D8][29];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_is_sta = _RANDOM[10'h1D8][30];	// lsu.scala:211:16
        stq_11_bits_uop_ctrl_is_std = _RANDOM[10'h1D8][31];	// lsu.scala:211:16
        stq_11_bits_uop_iw_state = _RANDOM[10'h1D9][1:0];	// lsu.scala:211:16
        stq_11_bits_uop_iw_p1_poisoned = _RANDOM[10'h1D9][2];	// lsu.scala:211:16
        stq_11_bits_uop_iw_p2_poisoned = _RANDOM[10'h1D9][3];	// lsu.scala:211:16
        stq_11_bits_uop_is_br = _RANDOM[10'h1D9][4];	// lsu.scala:211:16
        stq_11_bits_uop_is_jalr = _RANDOM[10'h1D9][5];	// lsu.scala:211:16
        stq_11_bits_uop_is_jal = _RANDOM[10'h1D9][6];	// lsu.scala:211:16
        stq_11_bits_uop_is_sfb = _RANDOM[10'h1D9][7];	// lsu.scala:211:16
        stq_11_bits_uop_br_mask = _RANDOM[10'h1D9][19:8];	// lsu.scala:211:16
        stq_11_bits_uop_br_tag = _RANDOM[10'h1D9][23:20];	// lsu.scala:211:16
        stq_11_bits_uop_ftq_idx = _RANDOM[10'h1D9][28:24];	// lsu.scala:211:16
        stq_11_bits_uop_edge_inst = _RANDOM[10'h1D9][29];	// lsu.scala:211:16
        stq_11_bits_uop_pc_lob = {_RANDOM[10'h1D9][31:30], _RANDOM[10'h1DA][3:0]};	// lsu.scala:211:16
        stq_11_bits_uop_taken = _RANDOM[10'h1DA][4];	// lsu.scala:211:16
        stq_11_bits_uop_imm_packed = _RANDOM[10'h1DA][24:5];	// lsu.scala:211:16
        stq_11_bits_uop_csr_addr = {_RANDOM[10'h1DA][31:25], _RANDOM[10'h1DB][4:0]};	// lsu.scala:211:16
        stq_11_bits_uop_rob_idx = _RANDOM[10'h1DB][10:5];	// lsu.scala:211:16
        stq_11_bits_uop_ldq_idx = _RANDOM[10'h1DB][14:11];	// lsu.scala:211:16
        stq_11_bits_uop_stq_idx = _RANDOM[10'h1DB][18:15];	// lsu.scala:211:16
        stq_11_bits_uop_rxq_idx = _RANDOM[10'h1DB][20:19];	// lsu.scala:211:16
        stq_11_bits_uop_pdst = _RANDOM[10'h1DB][27:21];	// lsu.scala:211:16
        stq_11_bits_uop_prs1 = {_RANDOM[10'h1DB][31:28], _RANDOM[10'h1DC][2:0]};	// lsu.scala:211:16
        stq_11_bits_uop_prs2 = _RANDOM[10'h1DC][9:3];	// lsu.scala:211:16
        stq_11_bits_uop_prs3 = _RANDOM[10'h1DC][16:10];	// lsu.scala:211:16
        stq_11_bits_uop_ppred = _RANDOM[10'h1DC][21:17];	// lsu.scala:211:16
        stq_11_bits_uop_prs1_busy = _RANDOM[10'h1DC][22];	// lsu.scala:211:16
        stq_11_bits_uop_prs2_busy = _RANDOM[10'h1DC][23];	// lsu.scala:211:16
        stq_11_bits_uop_prs3_busy = _RANDOM[10'h1DC][24];	// lsu.scala:211:16
        stq_11_bits_uop_ppred_busy = _RANDOM[10'h1DC][25];	// lsu.scala:211:16
        stq_11_bits_uop_stale_pdst = {_RANDOM[10'h1DC][31:26], _RANDOM[10'h1DD][0]};	// lsu.scala:211:16
        stq_11_bits_uop_exception = _RANDOM[10'h1DD][1];	// lsu.scala:211:16
        stq_11_bits_uop_exc_cause =
          {_RANDOM[10'h1DD][31:2], _RANDOM[10'h1DE], _RANDOM[10'h1DF][1:0]};	// lsu.scala:211:16
        stq_11_bits_uop_bypassable = _RANDOM[10'h1DF][2];	// lsu.scala:211:16
        stq_11_bits_uop_mem_cmd = _RANDOM[10'h1DF][7:3];	// lsu.scala:211:16
        stq_11_bits_uop_mem_size = _RANDOM[10'h1DF][9:8];	// lsu.scala:211:16
        stq_11_bits_uop_mem_signed = _RANDOM[10'h1DF][10];	// lsu.scala:211:16
        stq_11_bits_uop_is_fence = _RANDOM[10'h1DF][11];	// lsu.scala:211:16
        stq_11_bits_uop_is_fencei = _RANDOM[10'h1DF][12];	// lsu.scala:211:16
        stq_11_bits_uop_is_amo = _RANDOM[10'h1DF][13];	// lsu.scala:211:16
        stq_11_bits_uop_uses_ldq = _RANDOM[10'h1DF][14];	// lsu.scala:211:16
        stq_11_bits_uop_uses_stq = _RANDOM[10'h1DF][15];	// lsu.scala:211:16
        stq_11_bits_uop_is_sys_pc2epc = _RANDOM[10'h1DF][16];	// lsu.scala:211:16
        stq_11_bits_uop_is_unique = _RANDOM[10'h1DF][17];	// lsu.scala:211:16
        stq_11_bits_uop_flush_on_commit = _RANDOM[10'h1DF][18];	// lsu.scala:211:16
        stq_11_bits_uop_ldst_is_rs1 = _RANDOM[10'h1DF][19];	// lsu.scala:211:16
        stq_11_bits_uop_ldst = _RANDOM[10'h1DF][25:20];	// lsu.scala:211:16
        stq_11_bits_uop_lrs1 = _RANDOM[10'h1DF][31:26];	// lsu.scala:211:16
        stq_11_bits_uop_lrs2 = _RANDOM[10'h1E0][5:0];	// lsu.scala:211:16
        stq_11_bits_uop_lrs3 = _RANDOM[10'h1E0][11:6];	// lsu.scala:211:16
        stq_11_bits_uop_ldst_val = _RANDOM[10'h1E0][12];	// lsu.scala:211:16
        stq_11_bits_uop_dst_rtype = _RANDOM[10'h1E0][14:13];	// lsu.scala:211:16
        stq_11_bits_uop_lrs1_rtype = _RANDOM[10'h1E0][16:15];	// lsu.scala:211:16
        stq_11_bits_uop_lrs2_rtype = _RANDOM[10'h1E0][18:17];	// lsu.scala:211:16
        stq_11_bits_uop_frs3_en = _RANDOM[10'h1E0][19];	// lsu.scala:211:16
        stq_11_bits_uop_fp_val = _RANDOM[10'h1E0][20];	// lsu.scala:211:16
        stq_11_bits_uop_fp_single = _RANDOM[10'h1E0][21];	// lsu.scala:211:16
        stq_11_bits_uop_xcpt_pf_if = _RANDOM[10'h1E0][22];	// lsu.scala:211:16
        stq_11_bits_uop_xcpt_ae_if = _RANDOM[10'h1E0][23];	// lsu.scala:211:16
        stq_11_bits_uop_xcpt_ma_if = _RANDOM[10'h1E0][24];	// lsu.scala:211:16
        stq_11_bits_uop_bp_debug_if = _RANDOM[10'h1E0][25];	// lsu.scala:211:16
        stq_11_bits_uop_bp_xcpt_if = _RANDOM[10'h1E0][26];	// lsu.scala:211:16
        stq_11_bits_uop_debug_fsrc = _RANDOM[10'h1E0][28:27];	// lsu.scala:211:16
        stq_11_bits_uop_debug_tsrc = _RANDOM[10'h1E0][30:29];	// lsu.scala:211:16
        stq_11_bits_addr_valid = _RANDOM[10'h1E0][31];	// lsu.scala:211:16
        stq_11_bits_addr_bits = {_RANDOM[10'h1E1], _RANDOM[10'h1E2][7:0]};	// lsu.scala:211:16
        stq_11_bits_addr_is_virtual = _RANDOM[10'h1E2][8];	// lsu.scala:211:16
        stq_11_bits_data_valid = _RANDOM[10'h1E2][9];	// lsu.scala:211:16
        stq_11_bits_data_bits =
          {_RANDOM[10'h1E2][31:10], _RANDOM[10'h1E3], _RANDOM[10'h1E4][9:0]};	// lsu.scala:211:16
        stq_11_bits_committed = _RANDOM[10'h1E4][10];	// lsu.scala:211:16
        stq_11_bits_succeeded = _RANDOM[10'h1E4][11];	// lsu.scala:211:16
        stq_12_valid = _RANDOM[10'h1E6][12];	// lsu.scala:211:16
        stq_12_bits_uop_uopc = _RANDOM[10'h1E6][19:13];	// lsu.scala:211:16
        stq_12_bits_uop_inst = {_RANDOM[10'h1E6][31:20], _RANDOM[10'h1E7][19:0]};	// lsu.scala:211:16
        stq_12_bits_uop_debug_inst = {_RANDOM[10'h1E7][31:20], _RANDOM[10'h1E8][19:0]};	// lsu.scala:211:16
        stq_12_bits_uop_is_rvc = _RANDOM[10'h1E8][20];	// lsu.scala:211:16
        stq_12_bits_uop_debug_pc = {_RANDOM[10'h1E8][31:21], _RANDOM[10'h1E9][28:0]};	// lsu.scala:211:16
        stq_12_bits_uop_iq_type = _RANDOM[10'h1E9][31:29];	// lsu.scala:211:16
        stq_12_bits_uop_fu_code = _RANDOM[10'h1EA][9:0];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_br_type = _RANDOM[10'h1EA][13:10];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op1_sel = _RANDOM[10'h1EA][15:14];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op2_sel = _RANDOM[10'h1EA][18:16];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_imm_sel = _RANDOM[10'h1EA][21:19];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_op_fcn = _RANDOM[10'h1EA][25:22];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1EA][26];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1EA][29:27];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_is_load = _RANDOM[10'h1EA][30];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_is_sta = _RANDOM[10'h1EA][31];	// lsu.scala:211:16
        stq_12_bits_uop_ctrl_is_std = _RANDOM[10'h1EB][0];	// lsu.scala:211:16
        stq_12_bits_uop_iw_state = _RANDOM[10'h1EB][2:1];	// lsu.scala:211:16
        stq_12_bits_uop_iw_p1_poisoned = _RANDOM[10'h1EB][3];	// lsu.scala:211:16
        stq_12_bits_uop_iw_p2_poisoned = _RANDOM[10'h1EB][4];	// lsu.scala:211:16
        stq_12_bits_uop_is_br = _RANDOM[10'h1EB][5];	// lsu.scala:211:16
        stq_12_bits_uop_is_jalr = _RANDOM[10'h1EB][6];	// lsu.scala:211:16
        stq_12_bits_uop_is_jal = _RANDOM[10'h1EB][7];	// lsu.scala:211:16
        stq_12_bits_uop_is_sfb = _RANDOM[10'h1EB][8];	// lsu.scala:211:16
        stq_12_bits_uop_br_mask = _RANDOM[10'h1EB][20:9];	// lsu.scala:211:16
        stq_12_bits_uop_br_tag = _RANDOM[10'h1EB][24:21];	// lsu.scala:211:16
        stq_12_bits_uop_ftq_idx = _RANDOM[10'h1EB][29:25];	// lsu.scala:211:16
        stq_12_bits_uop_edge_inst = _RANDOM[10'h1EB][30];	// lsu.scala:211:16
        stq_12_bits_uop_pc_lob = {_RANDOM[10'h1EB][31], _RANDOM[10'h1EC][4:0]};	// lsu.scala:211:16
        stq_12_bits_uop_taken = _RANDOM[10'h1EC][5];	// lsu.scala:211:16
        stq_12_bits_uop_imm_packed = _RANDOM[10'h1EC][25:6];	// lsu.scala:211:16
        stq_12_bits_uop_csr_addr = {_RANDOM[10'h1EC][31:26], _RANDOM[10'h1ED][5:0]};	// lsu.scala:211:16
        stq_12_bits_uop_rob_idx = _RANDOM[10'h1ED][11:6];	// lsu.scala:211:16
        stq_12_bits_uop_ldq_idx = _RANDOM[10'h1ED][15:12];	// lsu.scala:211:16
        stq_12_bits_uop_stq_idx = _RANDOM[10'h1ED][19:16];	// lsu.scala:211:16
        stq_12_bits_uop_rxq_idx = _RANDOM[10'h1ED][21:20];	// lsu.scala:211:16
        stq_12_bits_uop_pdst = _RANDOM[10'h1ED][28:22];	// lsu.scala:211:16
        stq_12_bits_uop_prs1 = {_RANDOM[10'h1ED][31:29], _RANDOM[10'h1EE][3:0]};	// lsu.scala:211:16
        stq_12_bits_uop_prs2 = _RANDOM[10'h1EE][10:4];	// lsu.scala:211:16
        stq_12_bits_uop_prs3 = _RANDOM[10'h1EE][17:11];	// lsu.scala:211:16
        stq_12_bits_uop_ppred = _RANDOM[10'h1EE][22:18];	// lsu.scala:211:16
        stq_12_bits_uop_prs1_busy = _RANDOM[10'h1EE][23];	// lsu.scala:211:16
        stq_12_bits_uop_prs2_busy = _RANDOM[10'h1EE][24];	// lsu.scala:211:16
        stq_12_bits_uop_prs3_busy = _RANDOM[10'h1EE][25];	// lsu.scala:211:16
        stq_12_bits_uop_ppred_busy = _RANDOM[10'h1EE][26];	// lsu.scala:211:16
        stq_12_bits_uop_stale_pdst = {_RANDOM[10'h1EE][31:27], _RANDOM[10'h1EF][1:0]};	// lsu.scala:211:16
        stq_12_bits_uop_exception = _RANDOM[10'h1EF][2];	// lsu.scala:211:16
        stq_12_bits_uop_exc_cause =
          {_RANDOM[10'h1EF][31:3], _RANDOM[10'h1F0], _RANDOM[10'h1F1][2:0]};	// lsu.scala:211:16
        stq_12_bits_uop_bypassable = _RANDOM[10'h1F1][3];	// lsu.scala:211:16
        stq_12_bits_uop_mem_cmd = _RANDOM[10'h1F1][8:4];	// lsu.scala:211:16
        stq_12_bits_uop_mem_size = _RANDOM[10'h1F1][10:9];	// lsu.scala:211:16
        stq_12_bits_uop_mem_signed = _RANDOM[10'h1F1][11];	// lsu.scala:211:16
        stq_12_bits_uop_is_fence = _RANDOM[10'h1F1][12];	// lsu.scala:211:16
        stq_12_bits_uop_is_fencei = _RANDOM[10'h1F1][13];	// lsu.scala:211:16
        stq_12_bits_uop_is_amo = _RANDOM[10'h1F1][14];	// lsu.scala:211:16
        stq_12_bits_uop_uses_ldq = _RANDOM[10'h1F1][15];	// lsu.scala:211:16
        stq_12_bits_uop_uses_stq = _RANDOM[10'h1F1][16];	// lsu.scala:211:16
        stq_12_bits_uop_is_sys_pc2epc = _RANDOM[10'h1F1][17];	// lsu.scala:211:16
        stq_12_bits_uop_is_unique = _RANDOM[10'h1F1][18];	// lsu.scala:211:16
        stq_12_bits_uop_flush_on_commit = _RANDOM[10'h1F1][19];	// lsu.scala:211:16
        stq_12_bits_uop_ldst_is_rs1 = _RANDOM[10'h1F1][20];	// lsu.scala:211:16
        stq_12_bits_uop_ldst = _RANDOM[10'h1F1][26:21];	// lsu.scala:211:16
        stq_12_bits_uop_lrs1 = {_RANDOM[10'h1F1][31:27], _RANDOM[10'h1F2][0]};	// lsu.scala:211:16
        stq_12_bits_uop_lrs2 = _RANDOM[10'h1F2][6:1];	// lsu.scala:211:16
        stq_12_bits_uop_lrs3 = _RANDOM[10'h1F2][12:7];	// lsu.scala:211:16
        stq_12_bits_uop_ldst_val = _RANDOM[10'h1F2][13];	// lsu.scala:211:16
        stq_12_bits_uop_dst_rtype = _RANDOM[10'h1F2][15:14];	// lsu.scala:211:16
        stq_12_bits_uop_lrs1_rtype = _RANDOM[10'h1F2][17:16];	// lsu.scala:211:16
        stq_12_bits_uop_lrs2_rtype = _RANDOM[10'h1F2][19:18];	// lsu.scala:211:16
        stq_12_bits_uop_frs3_en = _RANDOM[10'h1F2][20];	// lsu.scala:211:16
        stq_12_bits_uop_fp_val = _RANDOM[10'h1F2][21];	// lsu.scala:211:16
        stq_12_bits_uop_fp_single = _RANDOM[10'h1F2][22];	// lsu.scala:211:16
        stq_12_bits_uop_xcpt_pf_if = _RANDOM[10'h1F2][23];	// lsu.scala:211:16
        stq_12_bits_uop_xcpt_ae_if = _RANDOM[10'h1F2][24];	// lsu.scala:211:16
        stq_12_bits_uop_xcpt_ma_if = _RANDOM[10'h1F2][25];	// lsu.scala:211:16
        stq_12_bits_uop_bp_debug_if = _RANDOM[10'h1F2][26];	// lsu.scala:211:16
        stq_12_bits_uop_bp_xcpt_if = _RANDOM[10'h1F2][27];	// lsu.scala:211:16
        stq_12_bits_uop_debug_fsrc = _RANDOM[10'h1F2][29:28];	// lsu.scala:211:16
        stq_12_bits_uop_debug_tsrc = _RANDOM[10'h1F2][31:30];	// lsu.scala:211:16
        stq_12_bits_addr_valid = _RANDOM[10'h1F3][0];	// lsu.scala:211:16
        stq_12_bits_addr_bits = {_RANDOM[10'h1F3][31:1], _RANDOM[10'h1F4][8:0]};	// lsu.scala:211:16
        stq_12_bits_addr_is_virtual = _RANDOM[10'h1F4][9];	// lsu.scala:211:16
        stq_12_bits_data_valid = _RANDOM[10'h1F4][10];	// lsu.scala:211:16
        stq_12_bits_data_bits =
          {_RANDOM[10'h1F4][31:11], _RANDOM[10'h1F5], _RANDOM[10'h1F6][10:0]};	// lsu.scala:211:16
        stq_12_bits_committed = _RANDOM[10'h1F6][11];	// lsu.scala:211:16
        stq_12_bits_succeeded = _RANDOM[10'h1F6][12];	// lsu.scala:211:16
        stq_13_valid = _RANDOM[10'h1F8][13];	// lsu.scala:211:16
        stq_13_bits_uop_uopc = _RANDOM[10'h1F8][20:14];	// lsu.scala:211:16
        stq_13_bits_uop_inst = {_RANDOM[10'h1F8][31:21], _RANDOM[10'h1F9][20:0]};	// lsu.scala:211:16
        stq_13_bits_uop_debug_inst = {_RANDOM[10'h1F9][31:21], _RANDOM[10'h1FA][20:0]};	// lsu.scala:211:16
        stq_13_bits_uop_is_rvc = _RANDOM[10'h1FA][21];	// lsu.scala:211:16
        stq_13_bits_uop_debug_pc = {_RANDOM[10'h1FA][31:22], _RANDOM[10'h1FB][29:0]};	// lsu.scala:211:16
        stq_13_bits_uop_iq_type = {_RANDOM[10'h1FB][31:30], _RANDOM[10'h1FC][0]};	// lsu.scala:211:16
        stq_13_bits_uop_fu_code = _RANDOM[10'h1FC][10:1];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_br_type = _RANDOM[10'h1FC][14:11];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op1_sel = _RANDOM[10'h1FC][16:15];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op2_sel = _RANDOM[10'h1FC][19:17];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_imm_sel = _RANDOM[10'h1FC][22:20];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_op_fcn = _RANDOM[10'h1FC][26:23];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_fcn_dw = _RANDOM[10'h1FC][27];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_csr_cmd = _RANDOM[10'h1FC][30:28];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_is_load = _RANDOM[10'h1FC][31];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_is_sta = _RANDOM[10'h1FD][0];	// lsu.scala:211:16
        stq_13_bits_uop_ctrl_is_std = _RANDOM[10'h1FD][1];	// lsu.scala:211:16
        stq_13_bits_uop_iw_state = _RANDOM[10'h1FD][3:2];	// lsu.scala:211:16
        stq_13_bits_uop_iw_p1_poisoned = _RANDOM[10'h1FD][4];	// lsu.scala:211:16
        stq_13_bits_uop_iw_p2_poisoned = _RANDOM[10'h1FD][5];	// lsu.scala:211:16
        stq_13_bits_uop_is_br = _RANDOM[10'h1FD][6];	// lsu.scala:211:16
        stq_13_bits_uop_is_jalr = _RANDOM[10'h1FD][7];	// lsu.scala:211:16
        stq_13_bits_uop_is_jal = _RANDOM[10'h1FD][8];	// lsu.scala:211:16
        stq_13_bits_uop_is_sfb = _RANDOM[10'h1FD][9];	// lsu.scala:211:16
        stq_13_bits_uop_br_mask = _RANDOM[10'h1FD][21:10];	// lsu.scala:211:16
        stq_13_bits_uop_br_tag = _RANDOM[10'h1FD][25:22];	// lsu.scala:211:16
        stq_13_bits_uop_ftq_idx = _RANDOM[10'h1FD][30:26];	// lsu.scala:211:16
        stq_13_bits_uop_edge_inst = _RANDOM[10'h1FD][31];	// lsu.scala:211:16
        stq_13_bits_uop_pc_lob = _RANDOM[10'h1FE][5:0];	// lsu.scala:211:16
        stq_13_bits_uop_taken = _RANDOM[10'h1FE][6];	// lsu.scala:211:16
        stq_13_bits_uop_imm_packed = _RANDOM[10'h1FE][26:7];	// lsu.scala:211:16
        stq_13_bits_uop_csr_addr = {_RANDOM[10'h1FE][31:27], _RANDOM[10'h1FF][6:0]};	// lsu.scala:211:16
        stq_13_bits_uop_rob_idx = _RANDOM[10'h1FF][12:7];	// lsu.scala:211:16
        stq_13_bits_uop_ldq_idx = _RANDOM[10'h1FF][16:13];	// lsu.scala:211:16
        stq_13_bits_uop_stq_idx = _RANDOM[10'h1FF][20:17];	// lsu.scala:211:16
        stq_13_bits_uop_rxq_idx = _RANDOM[10'h1FF][22:21];	// lsu.scala:211:16
        stq_13_bits_uop_pdst = _RANDOM[10'h1FF][29:23];	// lsu.scala:211:16
        stq_13_bits_uop_prs1 = {_RANDOM[10'h1FF][31:30], _RANDOM[10'h200][4:0]};	// lsu.scala:211:16
        stq_13_bits_uop_prs2 = _RANDOM[10'h200][11:5];	// lsu.scala:211:16
        stq_13_bits_uop_prs3 = _RANDOM[10'h200][18:12];	// lsu.scala:211:16
        stq_13_bits_uop_ppred = _RANDOM[10'h200][23:19];	// lsu.scala:211:16
        stq_13_bits_uop_prs1_busy = _RANDOM[10'h200][24];	// lsu.scala:211:16
        stq_13_bits_uop_prs2_busy = _RANDOM[10'h200][25];	// lsu.scala:211:16
        stq_13_bits_uop_prs3_busy = _RANDOM[10'h200][26];	// lsu.scala:211:16
        stq_13_bits_uop_ppred_busy = _RANDOM[10'h200][27];	// lsu.scala:211:16
        stq_13_bits_uop_stale_pdst = {_RANDOM[10'h200][31:28], _RANDOM[10'h201][2:0]};	// lsu.scala:211:16
        stq_13_bits_uop_exception = _RANDOM[10'h201][3];	// lsu.scala:211:16
        stq_13_bits_uop_exc_cause =
          {_RANDOM[10'h201][31:4], _RANDOM[10'h202], _RANDOM[10'h203][3:0]};	// lsu.scala:211:16
        stq_13_bits_uop_bypassable = _RANDOM[10'h203][4];	// lsu.scala:211:16
        stq_13_bits_uop_mem_cmd = _RANDOM[10'h203][9:5];	// lsu.scala:211:16
        stq_13_bits_uop_mem_size = _RANDOM[10'h203][11:10];	// lsu.scala:211:16
        stq_13_bits_uop_mem_signed = _RANDOM[10'h203][12];	// lsu.scala:211:16
        stq_13_bits_uop_is_fence = _RANDOM[10'h203][13];	// lsu.scala:211:16
        stq_13_bits_uop_is_fencei = _RANDOM[10'h203][14];	// lsu.scala:211:16
        stq_13_bits_uop_is_amo = _RANDOM[10'h203][15];	// lsu.scala:211:16
        stq_13_bits_uop_uses_ldq = _RANDOM[10'h203][16];	// lsu.scala:211:16
        stq_13_bits_uop_uses_stq = _RANDOM[10'h203][17];	// lsu.scala:211:16
        stq_13_bits_uop_is_sys_pc2epc = _RANDOM[10'h203][18];	// lsu.scala:211:16
        stq_13_bits_uop_is_unique = _RANDOM[10'h203][19];	// lsu.scala:211:16
        stq_13_bits_uop_flush_on_commit = _RANDOM[10'h203][20];	// lsu.scala:211:16
        stq_13_bits_uop_ldst_is_rs1 = _RANDOM[10'h203][21];	// lsu.scala:211:16
        stq_13_bits_uop_ldst = _RANDOM[10'h203][27:22];	// lsu.scala:211:16
        stq_13_bits_uop_lrs1 = {_RANDOM[10'h203][31:28], _RANDOM[10'h204][1:0]};	// lsu.scala:211:16
        stq_13_bits_uop_lrs2 = _RANDOM[10'h204][7:2];	// lsu.scala:211:16
        stq_13_bits_uop_lrs3 = _RANDOM[10'h204][13:8];	// lsu.scala:211:16
        stq_13_bits_uop_ldst_val = _RANDOM[10'h204][14];	// lsu.scala:211:16
        stq_13_bits_uop_dst_rtype = _RANDOM[10'h204][16:15];	// lsu.scala:211:16
        stq_13_bits_uop_lrs1_rtype = _RANDOM[10'h204][18:17];	// lsu.scala:211:16
        stq_13_bits_uop_lrs2_rtype = _RANDOM[10'h204][20:19];	// lsu.scala:211:16
        stq_13_bits_uop_frs3_en = _RANDOM[10'h204][21];	// lsu.scala:211:16
        stq_13_bits_uop_fp_val = _RANDOM[10'h204][22];	// lsu.scala:211:16
        stq_13_bits_uop_fp_single = _RANDOM[10'h204][23];	// lsu.scala:211:16
        stq_13_bits_uop_xcpt_pf_if = _RANDOM[10'h204][24];	// lsu.scala:211:16
        stq_13_bits_uop_xcpt_ae_if = _RANDOM[10'h204][25];	// lsu.scala:211:16
        stq_13_bits_uop_xcpt_ma_if = _RANDOM[10'h204][26];	// lsu.scala:211:16
        stq_13_bits_uop_bp_debug_if = _RANDOM[10'h204][27];	// lsu.scala:211:16
        stq_13_bits_uop_bp_xcpt_if = _RANDOM[10'h204][28];	// lsu.scala:211:16
        stq_13_bits_uop_debug_fsrc = _RANDOM[10'h204][30:29];	// lsu.scala:211:16
        stq_13_bits_uop_debug_tsrc = {_RANDOM[10'h204][31], _RANDOM[10'h205][0]};	// lsu.scala:211:16
        stq_13_bits_addr_valid = _RANDOM[10'h205][1];	// lsu.scala:211:16
        stq_13_bits_addr_bits = {_RANDOM[10'h205][31:2], _RANDOM[10'h206][9:0]};	// lsu.scala:211:16
        stq_13_bits_addr_is_virtual = _RANDOM[10'h206][10];	// lsu.scala:211:16
        stq_13_bits_data_valid = _RANDOM[10'h206][11];	// lsu.scala:211:16
        stq_13_bits_data_bits =
          {_RANDOM[10'h206][31:12], _RANDOM[10'h207], _RANDOM[10'h208][11:0]};	// lsu.scala:211:16
        stq_13_bits_committed = _RANDOM[10'h208][12];	// lsu.scala:211:16
        stq_13_bits_succeeded = _RANDOM[10'h208][13];	// lsu.scala:211:16
        stq_14_valid = _RANDOM[10'h20A][14];	// lsu.scala:211:16
        stq_14_bits_uop_uopc = _RANDOM[10'h20A][21:15];	// lsu.scala:211:16
        stq_14_bits_uop_inst = {_RANDOM[10'h20A][31:22], _RANDOM[10'h20B][21:0]};	// lsu.scala:211:16
        stq_14_bits_uop_debug_inst = {_RANDOM[10'h20B][31:22], _RANDOM[10'h20C][21:0]};	// lsu.scala:211:16
        stq_14_bits_uop_is_rvc = _RANDOM[10'h20C][22];	// lsu.scala:211:16
        stq_14_bits_uop_debug_pc = {_RANDOM[10'h20C][31:23], _RANDOM[10'h20D][30:0]};	// lsu.scala:211:16
        stq_14_bits_uop_iq_type = {_RANDOM[10'h20D][31], _RANDOM[10'h20E][1:0]};	// lsu.scala:211:16
        stq_14_bits_uop_fu_code = _RANDOM[10'h20E][11:2];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_br_type = _RANDOM[10'h20E][15:12];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op1_sel = _RANDOM[10'h20E][17:16];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op2_sel = _RANDOM[10'h20E][20:18];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_imm_sel = _RANDOM[10'h20E][23:21];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_op_fcn = _RANDOM[10'h20E][27:24];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_fcn_dw = _RANDOM[10'h20E][28];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_csr_cmd = _RANDOM[10'h20E][31:29];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_is_load = _RANDOM[10'h20F][0];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_is_sta = _RANDOM[10'h20F][1];	// lsu.scala:211:16
        stq_14_bits_uop_ctrl_is_std = _RANDOM[10'h20F][2];	// lsu.scala:211:16
        stq_14_bits_uop_iw_state = _RANDOM[10'h20F][4:3];	// lsu.scala:211:16
        stq_14_bits_uop_iw_p1_poisoned = _RANDOM[10'h20F][5];	// lsu.scala:211:16
        stq_14_bits_uop_iw_p2_poisoned = _RANDOM[10'h20F][6];	// lsu.scala:211:16
        stq_14_bits_uop_is_br = _RANDOM[10'h20F][7];	// lsu.scala:211:16
        stq_14_bits_uop_is_jalr = _RANDOM[10'h20F][8];	// lsu.scala:211:16
        stq_14_bits_uop_is_jal = _RANDOM[10'h20F][9];	// lsu.scala:211:16
        stq_14_bits_uop_is_sfb = _RANDOM[10'h20F][10];	// lsu.scala:211:16
        stq_14_bits_uop_br_mask = _RANDOM[10'h20F][22:11];	// lsu.scala:211:16
        stq_14_bits_uop_br_tag = _RANDOM[10'h20F][26:23];	// lsu.scala:211:16
        stq_14_bits_uop_ftq_idx = _RANDOM[10'h20F][31:27];	// lsu.scala:211:16
        stq_14_bits_uop_edge_inst = _RANDOM[10'h210][0];	// lsu.scala:211:16
        stq_14_bits_uop_pc_lob = _RANDOM[10'h210][6:1];	// lsu.scala:211:16
        stq_14_bits_uop_taken = _RANDOM[10'h210][7];	// lsu.scala:211:16
        stq_14_bits_uop_imm_packed = _RANDOM[10'h210][27:8];	// lsu.scala:211:16
        stq_14_bits_uop_csr_addr = {_RANDOM[10'h210][31:28], _RANDOM[10'h211][7:0]};	// lsu.scala:211:16
        stq_14_bits_uop_rob_idx = _RANDOM[10'h211][13:8];	// lsu.scala:211:16
        stq_14_bits_uop_ldq_idx = _RANDOM[10'h211][17:14];	// lsu.scala:211:16
        stq_14_bits_uop_stq_idx = _RANDOM[10'h211][21:18];	// lsu.scala:211:16
        stq_14_bits_uop_rxq_idx = _RANDOM[10'h211][23:22];	// lsu.scala:211:16
        stq_14_bits_uop_pdst = _RANDOM[10'h211][30:24];	// lsu.scala:211:16
        stq_14_bits_uop_prs1 = {_RANDOM[10'h211][31], _RANDOM[10'h212][5:0]};	// lsu.scala:211:16
        stq_14_bits_uop_prs2 = _RANDOM[10'h212][12:6];	// lsu.scala:211:16
        stq_14_bits_uop_prs3 = _RANDOM[10'h212][19:13];	// lsu.scala:211:16
        stq_14_bits_uop_ppred = _RANDOM[10'h212][24:20];	// lsu.scala:211:16
        stq_14_bits_uop_prs1_busy = _RANDOM[10'h212][25];	// lsu.scala:211:16
        stq_14_bits_uop_prs2_busy = _RANDOM[10'h212][26];	// lsu.scala:211:16
        stq_14_bits_uop_prs3_busy = _RANDOM[10'h212][27];	// lsu.scala:211:16
        stq_14_bits_uop_ppred_busy = _RANDOM[10'h212][28];	// lsu.scala:211:16
        stq_14_bits_uop_stale_pdst = {_RANDOM[10'h212][31:29], _RANDOM[10'h213][3:0]};	// lsu.scala:211:16
        stq_14_bits_uop_exception = _RANDOM[10'h213][4];	// lsu.scala:211:16
        stq_14_bits_uop_exc_cause =
          {_RANDOM[10'h213][31:5], _RANDOM[10'h214], _RANDOM[10'h215][4:0]};	// lsu.scala:211:16
        stq_14_bits_uop_bypassable = _RANDOM[10'h215][5];	// lsu.scala:211:16
        stq_14_bits_uop_mem_cmd = _RANDOM[10'h215][10:6];	// lsu.scala:211:16
        stq_14_bits_uop_mem_size = _RANDOM[10'h215][12:11];	// lsu.scala:211:16
        stq_14_bits_uop_mem_signed = _RANDOM[10'h215][13];	// lsu.scala:211:16
        stq_14_bits_uop_is_fence = _RANDOM[10'h215][14];	// lsu.scala:211:16
        stq_14_bits_uop_is_fencei = _RANDOM[10'h215][15];	// lsu.scala:211:16
        stq_14_bits_uop_is_amo = _RANDOM[10'h215][16];	// lsu.scala:211:16
        stq_14_bits_uop_uses_ldq = _RANDOM[10'h215][17];	// lsu.scala:211:16
        stq_14_bits_uop_uses_stq = _RANDOM[10'h215][18];	// lsu.scala:211:16
        stq_14_bits_uop_is_sys_pc2epc = _RANDOM[10'h215][19];	// lsu.scala:211:16
        stq_14_bits_uop_is_unique = _RANDOM[10'h215][20];	// lsu.scala:211:16
        stq_14_bits_uop_flush_on_commit = _RANDOM[10'h215][21];	// lsu.scala:211:16
        stq_14_bits_uop_ldst_is_rs1 = _RANDOM[10'h215][22];	// lsu.scala:211:16
        stq_14_bits_uop_ldst = _RANDOM[10'h215][28:23];	// lsu.scala:211:16
        stq_14_bits_uop_lrs1 = {_RANDOM[10'h215][31:29], _RANDOM[10'h216][2:0]};	// lsu.scala:211:16
        stq_14_bits_uop_lrs2 = _RANDOM[10'h216][8:3];	// lsu.scala:211:16
        stq_14_bits_uop_lrs3 = _RANDOM[10'h216][14:9];	// lsu.scala:211:16
        stq_14_bits_uop_ldst_val = _RANDOM[10'h216][15];	// lsu.scala:211:16
        stq_14_bits_uop_dst_rtype = _RANDOM[10'h216][17:16];	// lsu.scala:211:16
        stq_14_bits_uop_lrs1_rtype = _RANDOM[10'h216][19:18];	// lsu.scala:211:16
        stq_14_bits_uop_lrs2_rtype = _RANDOM[10'h216][21:20];	// lsu.scala:211:16
        stq_14_bits_uop_frs3_en = _RANDOM[10'h216][22];	// lsu.scala:211:16
        stq_14_bits_uop_fp_val = _RANDOM[10'h216][23];	// lsu.scala:211:16
        stq_14_bits_uop_fp_single = _RANDOM[10'h216][24];	// lsu.scala:211:16
        stq_14_bits_uop_xcpt_pf_if = _RANDOM[10'h216][25];	// lsu.scala:211:16
        stq_14_bits_uop_xcpt_ae_if = _RANDOM[10'h216][26];	// lsu.scala:211:16
        stq_14_bits_uop_xcpt_ma_if = _RANDOM[10'h216][27];	// lsu.scala:211:16
        stq_14_bits_uop_bp_debug_if = _RANDOM[10'h216][28];	// lsu.scala:211:16
        stq_14_bits_uop_bp_xcpt_if = _RANDOM[10'h216][29];	// lsu.scala:211:16
        stq_14_bits_uop_debug_fsrc = _RANDOM[10'h216][31:30];	// lsu.scala:211:16
        stq_14_bits_uop_debug_tsrc = _RANDOM[10'h217][1:0];	// lsu.scala:211:16
        stq_14_bits_addr_valid = _RANDOM[10'h217][2];	// lsu.scala:211:16
        stq_14_bits_addr_bits = {_RANDOM[10'h217][31:3], _RANDOM[10'h218][10:0]};	// lsu.scala:211:16
        stq_14_bits_addr_is_virtual = _RANDOM[10'h218][11];	// lsu.scala:211:16
        stq_14_bits_data_valid = _RANDOM[10'h218][12];	// lsu.scala:211:16
        stq_14_bits_data_bits =
          {_RANDOM[10'h218][31:13], _RANDOM[10'h219], _RANDOM[10'h21A][12:0]};	// lsu.scala:211:16
        stq_14_bits_committed = _RANDOM[10'h21A][13];	// lsu.scala:211:16
        stq_14_bits_succeeded = _RANDOM[10'h21A][14];	// lsu.scala:211:16
        stq_15_valid = _RANDOM[10'h21C][15];	// lsu.scala:211:16
        stq_15_bits_uop_uopc = _RANDOM[10'h21C][22:16];	// lsu.scala:211:16
        stq_15_bits_uop_inst = {_RANDOM[10'h21C][31:23], _RANDOM[10'h21D][22:0]};	// lsu.scala:211:16
        stq_15_bits_uop_debug_inst = {_RANDOM[10'h21D][31:23], _RANDOM[10'h21E][22:0]};	// lsu.scala:211:16
        stq_15_bits_uop_is_rvc = _RANDOM[10'h21E][23];	// lsu.scala:211:16
        stq_15_bits_uop_debug_pc = {_RANDOM[10'h21E][31:24], _RANDOM[10'h21F]};	// lsu.scala:211:16
        stq_15_bits_uop_iq_type = _RANDOM[10'h220][2:0];	// lsu.scala:211:16
        stq_15_bits_uop_fu_code = _RANDOM[10'h220][12:3];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_br_type = _RANDOM[10'h220][16:13];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op1_sel = _RANDOM[10'h220][18:17];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op2_sel = _RANDOM[10'h220][21:19];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_imm_sel = _RANDOM[10'h220][24:22];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_op_fcn = _RANDOM[10'h220][28:25];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_fcn_dw = _RANDOM[10'h220][29];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_csr_cmd = {_RANDOM[10'h220][31:30], _RANDOM[10'h221][0]};	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_is_load = _RANDOM[10'h221][1];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_is_sta = _RANDOM[10'h221][2];	// lsu.scala:211:16
        stq_15_bits_uop_ctrl_is_std = _RANDOM[10'h221][3];	// lsu.scala:211:16
        stq_15_bits_uop_iw_state = _RANDOM[10'h221][5:4];	// lsu.scala:211:16
        stq_15_bits_uop_iw_p1_poisoned = _RANDOM[10'h221][6];	// lsu.scala:211:16
        stq_15_bits_uop_iw_p2_poisoned = _RANDOM[10'h221][7];	// lsu.scala:211:16
        stq_15_bits_uop_is_br = _RANDOM[10'h221][8];	// lsu.scala:211:16
        stq_15_bits_uop_is_jalr = _RANDOM[10'h221][9];	// lsu.scala:211:16
        stq_15_bits_uop_is_jal = _RANDOM[10'h221][10];	// lsu.scala:211:16
        stq_15_bits_uop_is_sfb = _RANDOM[10'h221][11];	// lsu.scala:211:16
        stq_15_bits_uop_br_mask = _RANDOM[10'h221][23:12];	// lsu.scala:211:16
        stq_15_bits_uop_br_tag = _RANDOM[10'h221][27:24];	// lsu.scala:211:16
        stq_15_bits_uop_ftq_idx = {_RANDOM[10'h221][31:28], _RANDOM[10'h222][0]};	// lsu.scala:211:16
        stq_15_bits_uop_edge_inst = _RANDOM[10'h222][1];	// lsu.scala:211:16
        stq_15_bits_uop_pc_lob = _RANDOM[10'h222][7:2];	// lsu.scala:211:16
        stq_15_bits_uop_taken = _RANDOM[10'h222][8];	// lsu.scala:211:16
        stq_15_bits_uop_imm_packed = _RANDOM[10'h222][28:9];	// lsu.scala:211:16
        stq_15_bits_uop_csr_addr = {_RANDOM[10'h222][31:29], _RANDOM[10'h223][8:0]};	// lsu.scala:211:16
        stq_15_bits_uop_rob_idx = _RANDOM[10'h223][14:9];	// lsu.scala:211:16
        stq_15_bits_uop_ldq_idx = _RANDOM[10'h223][18:15];	// lsu.scala:211:16
        stq_15_bits_uop_stq_idx = _RANDOM[10'h223][22:19];	// lsu.scala:211:16
        stq_15_bits_uop_rxq_idx = _RANDOM[10'h223][24:23];	// lsu.scala:211:16
        stq_15_bits_uop_pdst = _RANDOM[10'h223][31:25];	// lsu.scala:211:16
        stq_15_bits_uop_prs1 = _RANDOM[10'h224][6:0];	// lsu.scala:211:16
        stq_15_bits_uop_prs2 = _RANDOM[10'h224][13:7];	// lsu.scala:211:16
        stq_15_bits_uop_prs3 = _RANDOM[10'h224][20:14];	// lsu.scala:211:16
        stq_15_bits_uop_ppred = _RANDOM[10'h224][25:21];	// lsu.scala:211:16
        stq_15_bits_uop_prs1_busy = _RANDOM[10'h224][26];	// lsu.scala:211:16
        stq_15_bits_uop_prs2_busy = _RANDOM[10'h224][27];	// lsu.scala:211:16
        stq_15_bits_uop_prs3_busy = _RANDOM[10'h224][28];	// lsu.scala:211:16
        stq_15_bits_uop_ppred_busy = _RANDOM[10'h224][29];	// lsu.scala:211:16
        stq_15_bits_uop_stale_pdst = {_RANDOM[10'h224][31:30], _RANDOM[10'h225][4:0]};	// lsu.scala:211:16
        stq_15_bits_uop_exception = _RANDOM[10'h225][5];	// lsu.scala:211:16
        stq_15_bits_uop_exc_cause =
          {_RANDOM[10'h225][31:6], _RANDOM[10'h226], _RANDOM[10'h227][5:0]};	// lsu.scala:211:16
        stq_15_bits_uop_bypassable = _RANDOM[10'h227][6];	// lsu.scala:211:16
        stq_15_bits_uop_mem_cmd = _RANDOM[10'h227][11:7];	// lsu.scala:211:16
        stq_15_bits_uop_mem_size = _RANDOM[10'h227][13:12];	// lsu.scala:211:16
        stq_15_bits_uop_mem_signed = _RANDOM[10'h227][14];	// lsu.scala:211:16
        stq_15_bits_uop_is_fence = _RANDOM[10'h227][15];	// lsu.scala:211:16
        stq_15_bits_uop_is_fencei = _RANDOM[10'h227][16];	// lsu.scala:211:16
        stq_15_bits_uop_is_amo = _RANDOM[10'h227][17];	// lsu.scala:211:16
        stq_15_bits_uop_uses_ldq = _RANDOM[10'h227][18];	// lsu.scala:211:16
        stq_15_bits_uop_uses_stq = _RANDOM[10'h227][19];	// lsu.scala:211:16
        stq_15_bits_uop_is_sys_pc2epc = _RANDOM[10'h227][20];	// lsu.scala:211:16
        stq_15_bits_uop_is_unique = _RANDOM[10'h227][21];	// lsu.scala:211:16
        stq_15_bits_uop_flush_on_commit = _RANDOM[10'h227][22];	// lsu.scala:211:16
        stq_15_bits_uop_ldst_is_rs1 = _RANDOM[10'h227][23];	// lsu.scala:211:16
        stq_15_bits_uop_ldst = _RANDOM[10'h227][29:24];	// lsu.scala:211:16
        stq_15_bits_uop_lrs1 = {_RANDOM[10'h227][31:30], _RANDOM[10'h228][3:0]};	// lsu.scala:211:16
        stq_15_bits_uop_lrs2 = _RANDOM[10'h228][9:4];	// lsu.scala:211:16
        stq_15_bits_uop_lrs3 = _RANDOM[10'h228][15:10];	// lsu.scala:211:16
        stq_15_bits_uop_ldst_val = _RANDOM[10'h228][16];	// lsu.scala:211:16
        stq_15_bits_uop_dst_rtype = _RANDOM[10'h228][18:17];	// lsu.scala:211:16
        stq_15_bits_uop_lrs1_rtype = _RANDOM[10'h228][20:19];	// lsu.scala:211:16
        stq_15_bits_uop_lrs2_rtype = _RANDOM[10'h228][22:21];	// lsu.scala:211:16
        stq_15_bits_uop_frs3_en = _RANDOM[10'h228][23];	// lsu.scala:211:16
        stq_15_bits_uop_fp_val = _RANDOM[10'h228][24];	// lsu.scala:211:16
        stq_15_bits_uop_fp_single = _RANDOM[10'h228][25];	// lsu.scala:211:16
        stq_15_bits_uop_xcpt_pf_if = _RANDOM[10'h228][26];	// lsu.scala:211:16
        stq_15_bits_uop_xcpt_ae_if = _RANDOM[10'h228][27];	// lsu.scala:211:16
        stq_15_bits_uop_xcpt_ma_if = _RANDOM[10'h228][28];	// lsu.scala:211:16
        stq_15_bits_uop_bp_debug_if = _RANDOM[10'h228][29];	// lsu.scala:211:16
        stq_15_bits_uop_bp_xcpt_if = _RANDOM[10'h228][30];	// lsu.scala:211:16
        stq_15_bits_uop_debug_fsrc = {_RANDOM[10'h228][31], _RANDOM[10'h229][0]};	// lsu.scala:211:16
        stq_15_bits_uop_debug_tsrc = _RANDOM[10'h229][2:1];	// lsu.scala:211:16
        stq_15_bits_addr_valid = _RANDOM[10'h229][3];	// lsu.scala:211:16
        stq_15_bits_addr_bits = {_RANDOM[10'h229][31:4], _RANDOM[10'h22A][11:0]};	// lsu.scala:211:16
        stq_15_bits_addr_is_virtual = _RANDOM[10'h22A][12];	// lsu.scala:211:16
        stq_15_bits_data_valid = _RANDOM[10'h22A][13];	// lsu.scala:211:16
        stq_15_bits_data_bits =
          {_RANDOM[10'h22A][31:14], _RANDOM[10'h22B], _RANDOM[10'h22C][13:0]};	// lsu.scala:211:16
        stq_15_bits_committed = _RANDOM[10'h22C][14];	// lsu.scala:211:16
        stq_15_bits_succeeded = _RANDOM[10'h22C][15];	// lsu.scala:211:16
        ldq_head = _RANDOM[10'h22E][19:16];	// lsu.scala:215:29
        ldq_tail = _RANDOM[10'h22E][23:20];	// lsu.scala:215:29, :216:29
        stq_head = _RANDOM[10'h22E][27:24];	// lsu.scala:215:29, :217:29
        stq_tail = _RANDOM[10'h22E][31:28];	// lsu.scala:215:29, :218:29
        stq_commit_head = _RANDOM[10'h22F][3:0];	// lsu.scala:219:29
        stq_execute_head = _RANDOM[10'h22F][7:4];	// lsu.scala:219:29, :220:29
        hella_state = _RANDOM[10'h22F][10:8];	// lsu.scala:219:29, :242:38
        hella_req_addr = {_RANDOM[10'h22F][31:11], _RANDOM[10'h230][18:0]};	// lsu.scala:219:29, :243:34
        hella_req_cmd = _RANDOM[10'h230][30:26];	// lsu.scala:243:34
        hella_req_size = {_RANDOM[10'h230][31], _RANDOM[10'h231][0]};	// lsu.scala:243:34
        hella_req_signed = _RANDOM[10'h231][1];	// lsu.scala:243:34
        hella_req_phys = _RANDOM[10'h231][4];	// lsu.scala:243:34
        hella_data_data =
          {_RANDOM[10'h233][31:15], _RANDOM[10'h234], _RANDOM[10'h235][14:0]};	// lsu.scala:244:34
        hella_paddr = {_RANDOM[10'h235][31:23], _RANDOM[10'h236][22:0]};	// lsu.scala:244:34, :245:34
        hella_xcpt_ma_ld = _RANDOM[10'h236][23];	// lsu.scala:245:34, :246:34
        hella_xcpt_ma_st = _RANDOM[10'h236][24];	// lsu.scala:245:34, :246:34
        hella_xcpt_pf_ld = _RANDOM[10'h236][25];	// lsu.scala:245:34, :246:34
        hella_xcpt_pf_st = _RANDOM[10'h236][26];	// lsu.scala:245:34, :246:34
        hella_xcpt_ae_ld = _RANDOM[10'h236][27];	// lsu.scala:245:34, :246:34
        hella_xcpt_ae_st = _RANDOM[10'h236][28];	// lsu.scala:245:34, :246:34
        live_store_mask = {_RANDOM[10'h236][31:29], _RANDOM[10'h237][12:0]};	// lsu.scala:245:34, :259:32
        p1_block_load_mask_0 = _RANDOM[10'h237][13];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_1 = _RANDOM[10'h237][14];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_2 = _RANDOM[10'h237][15];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_3 = _RANDOM[10'h237][16];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_4 = _RANDOM[10'h237][17];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_5 = _RANDOM[10'h237][18];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_6 = _RANDOM[10'h237][19];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_7 = _RANDOM[10'h237][20];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_8 = _RANDOM[10'h237][21];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_9 = _RANDOM[10'h237][22];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_10 = _RANDOM[10'h237][23];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_11 = _RANDOM[10'h237][24];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_12 = _RANDOM[10'h237][25];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_13 = _RANDOM[10'h237][26];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_14 = _RANDOM[10'h237][27];	// lsu.scala:259:32, :398:35
        p1_block_load_mask_15 = _RANDOM[10'h237][28];	// lsu.scala:259:32, :398:35
        p2_block_load_mask_0 = _RANDOM[10'h237][29];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_1 = _RANDOM[10'h237][30];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_2 = _RANDOM[10'h237][31];	// lsu.scala:259:32, :399:35
        p2_block_load_mask_3 = _RANDOM[10'h238][0];	// lsu.scala:399:35
        p2_block_load_mask_4 = _RANDOM[10'h238][1];	// lsu.scala:399:35
        p2_block_load_mask_5 = _RANDOM[10'h238][2];	// lsu.scala:399:35
        p2_block_load_mask_6 = _RANDOM[10'h238][3];	// lsu.scala:399:35
        p2_block_load_mask_7 = _RANDOM[10'h238][4];	// lsu.scala:399:35
        p2_block_load_mask_8 = _RANDOM[10'h238][5];	// lsu.scala:399:35
        p2_block_load_mask_9 = _RANDOM[10'h238][6];	// lsu.scala:399:35
        p2_block_load_mask_10 = _RANDOM[10'h238][7];	// lsu.scala:399:35
        p2_block_load_mask_11 = _RANDOM[10'h238][8];	// lsu.scala:399:35
        p2_block_load_mask_12 = _RANDOM[10'h238][9];	// lsu.scala:399:35
        p2_block_load_mask_13 = _RANDOM[10'h238][10];	// lsu.scala:399:35
        p2_block_load_mask_14 = _RANDOM[10'h238][11];	// lsu.scala:399:35
        p2_block_load_mask_15 = _RANDOM[10'h238][12];	// lsu.scala:399:35
        ldq_retry_idx = _RANDOM[10'h238][17:14];	// lsu.scala:399:35, :415:30
        stq_retry_idx = _RANDOM[10'h238][21:18];	// lsu.scala:399:35, :422:30
        ldq_wakeup_idx = _RANDOM[10'h238][25:22];	// lsu.scala:399:35, :430:31
        can_fire_load_retry_REG = _RANDOM[10'h238][26];	// lsu.scala:399:35, :470:40
        can_fire_sta_retry_REG = _RANDOM[10'h238][27];	// lsu.scala:399:35, :482:41
        mem_xcpt_valids_0 = _RANDOM[10'h238][28];	// lsu.scala:399:35, :667:32
        mem_xcpt_uops_0_br_mask = {_RANDOM[10'h23D][31:25], _RANDOM[10'h23E][4:0]};	// lsu.scala:671:32
        mem_xcpt_uops_0_rob_idx = _RANDOM[10'h23F][27:22];	// lsu.scala:671:32
        mem_xcpt_uops_0_ldq_idx = _RANDOM[10'h23F][31:28];	// lsu.scala:671:32
        mem_xcpt_uops_0_stq_idx = _RANDOM[10'h240][3:0];	// lsu.scala:671:32
        mem_xcpt_uops_0_uses_ldq = _RANDOM[10'h243][31];	// lsu.scala:671:32
        mem_xcpt_uops_0_uses_stq = _RANDOM[10'h244][0];	// lsu.scala:671:32
        mem_xcpt_causes_0 = _RANDOM[10'h245][19:16];	// lsu.scala:672:32
        mem_xcpt_vaddrs_0 = {_RANDOM[10'h245][31:20], _RANDOM[10'h246][27:0]};	// lsu.scala:672:32, :679:32
        REG = _RANDOM[10'h246][28];	// lsu.scala:679:32, :718:21
        fired_load_incoming_REG = _RANDOM[10'h246][29];	// lsu.scala:679:32, :894:51
        fired_stad_incoming_REG = _RANDOM[10'h246][30];	// lsu.scala:679:32, :895:51
        fired_sta_incoming_REG = _RANDOM[10'h246][31];	// lsu.scala:679:32, :896:51
        fired_std_incoming_REG = _RANDOM[10'h247][0];	// lsu.scala:897:51
        fired_stdf_incoming = _RANDOM[10'h247][1];	// lsu.scala:897:51, :898:37
        fired_sfence_0 = _RANDOM[10'h247][2];	// lsu.scala:897:51, :899:37
        fired_release_0 = _RANDOM[10'h247][3];	// lsu.scala:897:51, :900:37
        fired_load_retry_REG = _RANDOM[10'h247][4];	// lsu.scala:897:51, :901:51
        fired_sta_retry_REG = _RANDOM[10'h247][5];	// lsu.scala:897:51, :902:51
        fired_load_wakeup_REG = _RANDOM[10'h247][7];	// lsu.scala:897:51, :904:51
        mem_incoming_uop_0_br_mask = _RANDOM[10'h24C][17:6];	// lsu.scala:908:37
        mem_incoming_uop_0_rob_idx = _RANDOM[10'h24E][8:3];	// lsu.scala:908:37
        mem_incoming_uop_0_ldq_idx = _RANDOM[10'h24E][12:9];	// lsu.scala:908:37
        mem_incoming_uop_0_stq_idx = _RANDOM[10'h24E][16:13];	// lsu.scala:908:37
        mem_incoming_uop_0_pdst = _RANDOM[10'h24E][25:19];	// lsu.scala:908:37
        mem_incoming_uop_0_fp_val = _RANDOM[10'h253][18];	// lsu.scala:908:37
        mem_ldq_incoming_e_0_bits_uop_br_mask =
          {_RANDOM[10'h258][31:26], _RANDOM[10'h259][5:0]};	// lsu.scala:909:37
        mem_ldq_incoming_e_0_bits_uop_stq_idx = _RANDOM[10'h25B][4:1];	// lsu.scala:909:37
        mem_ldq_incoming_e_0_bits_uop_mem_size = _RANDOM[10'h25E][27:26];	// lsu.scala:909:37
        mem_ldq_incoming_e_0_bits_st_dep_mask = _RANDOM[10'h262][15:0];	// lsu.scala:909:37
        mem_stq_incoming_e_0_valid = _RANDOM[10'h264][25];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_br_mask =
          {_RANDOM[10'h269][31:22], _RANDOM[10'h26A][1:0]};	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_rob_idx = _RANDOM[10'h26B][24:19];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_stq_idx =
          {_RANDOM[10'h26B][31:29], _RANDOM[10'h26C][0]};	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_mem_size = _RANDOM[10'h26F][23:22];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_uop_is_amo = _RANDOM[10'h26F][27];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_addr_valid = _RANDOM[10'h271][13];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_addr_is_virtual = _RANDOM[10'h272][22];	// lsu.scala:910:37
        mem_stq_incoming_e_0_bits_data_valid = _RANDOM[10'h272][23];	// lsu.scala:910:37
        mem_ldq_wakeup_e_bits_uop_br_mask =
          {_RANDOM[10'h27B][31:23], _RANDOM[10'h27C][2:0]};	// lsu.scala:911:37
        mem_ldq_wakeup_e_bits_uop_stq_idx =
          {_RANDOM[10'h27D][31:30], _RANDOM[10'h27E][1:0]};	// lsu.scala:911:37
        mem_ldq_wakeup_e_bits_uop_mem_size = _RANDOM[10'h281][24:23];	// lsu.scala:911:37
        mem_ldq_wakeup_e_bits_st_dep_mask =
          {_RANDOM[10'h284][31:29], _RANDOM[10'h285][12:0]};	// lsu.scala:911:37
        mem_ldq_retry_e_bits_uop_br_mask = _RANDOM[10'h28C][30:19];	// lsu.scala:912:37
        mem_ldq_retry_e_bits_uop_stq_idx = _RANDOM[10'h28E][29:26];	// lsu.scala:912:37
        mem_ldq_retry_e_bits_uop_mem_size = _RANDOM[10'h292][20:19];	// lsu.scala:912:37
        mem_ldq_retry_e_bits_st_dep_mask =
          {_RANDOM[10'h295][31:25], _RANDOM[10'h296][8:0]};	// lsu.scala:912:37
        mem_stq_retry_e_valid = _RANDOM[10'h298][18];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_br_mask = _RANDOM[10'h29D][26:15];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_rob_idx = _RANDOM[10'h29F][17:12];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_stq_idx = _RANDOM[10'h29F][25:22];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_mem_size = _RANDOM[10'h2A3][16:15];	// lsu.scala:913:37
        mem_stq_retry_e_bits_uop_is_amo = _RANDOM[10'h2A3][20];	// lsu.scala:913:37
        mem_stq_retry_e_bits_data_valid = _RANDOM[10'h2A6][16];	// lsu.scala:913:37
        mem_stdf_uop_br_mask = _RANDOM[10'h2AF][26:15];	// lsu.scala:922:37
        mem_stdf_uop_rob_idx = _RANDOM[10'h2B1][17:12];	// lsu.scala:922:37
        mem_stdf_uop_stq_idx = _RANDOM[10'h2B1][25:22];	// lsu.scala:922:37
        mem_tlb_miss_0 = _RANDOM[10'h2B7][6];	// lsu.scala:925:41
        mem_tlb_uncacheable_0 = _RANDOM[10'h2B7][7];	// lsu.scala:925:41, :926:41
        mem_paddr_0 = {_RANDOM[10'h2B7][31:8], _RANDOM[10'h2B8][15:0]};	// lsu.scala:925:41, :927:41
        clr_bsy_valid_0 = _RANDOM[10'h2B8][16];	// lsu.scala:927:41, :930:32
        clr_bsy_rob_idx_0 = _RANDOM[10'h2B8][22:17];	// lsu.scala:927:41, :931:28
        clr_bsy_brmask_0 = {_RANDOM[10'h2B8][31:23], _RANDOM[10'h2B9][2:0]};	// lsu.scala:927:41, :932:28
        io_core_clr_bsy_0_valid_REG = _RANDOM[10'h2B9][3];	// lsu.scala:932:28, :979:62
        io_core_clr_bsy_0_valid_REG_1 = _RANDOM[10'h2B9][4];	// lsu.scala:932:28, :979:101
        io_core_clr_bsy_0_valid_REG_2 = _RANDOM[10'h2B9][5];	// lsu.scala:932:28, :979:93
        stdf_clr_bsy_valid = _RANDOM[10'h2B9][6];	// lsu.scala:932:28, :983:37
        stdf_clr_bsy_rob_idx = _RANDOM[10'h2B9][12:7];	// lsu.scala:932:28, :984:33
        stdf_clr_bsy_brmask = _RANDOM[10'h2B9][24:13];	// lsu.scala:932:28, :985:33
        io_core_clr_bsy_1_valid_REG = _RANDOM[10'h2B9][25];	// lsu.scala:932:28, :1004:67
        io_core_clr_bsy_1_valid_REG_1 = _RANDOM[10'h2B9][26];	// lsu.scala:932:28, :1004:106
        io_core_clr_bsy_1_valid_REG_2 = _RANDOM[10'h2B9][27];	// lsu.scala:932:28, :1004:98
        lcam_addr_REG = {_RANDOM[10'h2B9][31:28], _RANDOM[10'h2BA][27:0]};	// lsu.scala:932:28, :1026:45
        lcam_addr_REG_1 = {_RANDOM[10'h2BA][31:28], _RANDOM[10'h2BB][27:0]};	// lsu.scala:1026:45, :1027:67
        lcam_ldq_idx_REG = _RANDOM[10'h2BB][31:28];	// lsu.scala:1027:67, :1037:58
        lcam_ldq_idx_REG_1 = _RANDOM[10'h2BC][3:0];	// lsu.scala:1038:58
        lcam_stq_idx_REG = _RANDOM[10'h2BC][7:4];	// lsu.scala:1038:58, :1042:58
        s1_executing_loads_0 = _RANDOM[10'h2BC][8];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_1 = _RANDOM[10'h2BC][9];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_2 = _RANDOM[10'h2BC][10];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_3 = _RANDOM[10'h2BC][11];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_4 = _RANDOM[10'h2BC][12];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_5 = _RANDOM[10'h2BC][13];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_6 = _RANDOM[10'h2BC][14];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_7 = _RANDOM[10'h2BC][15];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_8 = _RANDOM[10'h2BC][16];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_9 = _RANDOM[10'h2BC][17];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_10 = _RANDOM[10'h2BC][18];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_11 = _RANDOM[10'h2BC][19];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_12 = _RANDOM[10'h2BC][20];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_13 = _RANDOM[10'h2BC][21];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_14 = _RANDOM[10'h2BC][22];	// lsu.scala:1038:58, :1056:35
        s1_executing_loads_15 = _RANDOM[10'h2BC][23];	// lsu.scala:1038:58, :1056:35
        wb_forward_valid_0 = _RANDOM[10'h2BC][24];	// lsu.scala:1038:58, :1064:36
        wb_forward_ldq_idx_0 = _RANDOM[10'h2BC][28:25];	// lsu.scala:1038:58, :1065:36
        wb_forward_ld_addr_0 =
          {_RANDOM[10'h2BC][31:29], _RANDOM[10'h2BD], _RANDOM[10'h2BE][4:0]};	// lsu.scala:1038:58, :1066:36
        wb_forward_stq_idx_0 = _RANDOM[10'h2BE][8:5];	// lsu.scala:1066:36, :1067:36
        older_nacked_REG = _RANDOM[10'h2BE][9];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG = _RANDOM[10'h2BE][10];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_1 = _RANDOM[10'h2BE][11];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_1 = _RANDOM[10'h2BE][12];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_2 = _RANDOM[10'h2BE][13];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_2 = _RANDOM[10'h2BE][14];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_3 = _RANDOM[10'h2BE][15];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_3 = _RANDOM[10'h2BE][16];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_4 = _RANDOM[10'h2BE][17];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_4 = _RANDOM[10'h2BE][18];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_5 = _RANDOM[10'h2BE][19];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_5 = _RANDOM[10'h2BE][20];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_6 = _RANDOM[10'h2BE][21];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_6 = _RANDOM[10'h2BE][22];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_7 = _RANDOM[10'h2BE][23];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_7 = _RANDOM[10'h2BE][24];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_8 = _RANDOM[10'h2BE][25];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_8 = _RANDOM[10'h2BE][26];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_9 = _RANDOM[10'h2BE][27];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_9 = _RANDOM[10'h2BE][28];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_10 = _RANDOM[10'h2BE][29];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_10 = _RANDOM[10'h2BE][30];	// lsu.scala:1066:36, :1131:58
        older_nacked_REG_11 = _RANDOM[10'h2BE][31];	// lsu.scala:1066:36, :1128:57
        io_dmem_s1_kill_0_REG_11 = _RANDOM[10'h2BF][0];	// lsu.scala:1131:58
        older_nacked_REG_12 = _RANDOM[10'h2BF][1];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_12 = _RANDOM[10'h2BF][2];	// lsu.scala:1131:58
        older_nacked_REG_13 = _RANDOM[10'h2BF][3];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_13 = _RANDOM[10'h2BF][4];	// lsu.scala:1131:58
        older_nacked_REG_14 = _RANDOM[10'h2BF][5];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_14 = _RANDOM[10'h2BF][6];	// lsu.scala:1131:58
        older_nacked_REG_15 = _RANDOM[10'h2BF][7];	// lsu.scala:1128:57, :1131:58
        io_dmem_s1_kill_0_REG_15 = _RANDOM[10'h2BF][8];	// lsu.scala:1131:58
        io_dmem_s1_kill_0_REG_16 = _RANDOM[10'h2BF][9];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_17 = _RANDOM[10'h2BF][10];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_18 = _RANDOM[10'h2BF][11];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_19 = _RANDOM[10'h2BF][12];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_20 = _RANDOM[10'h2BF][13];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_21 = _RANDOM[10'h2BF][14];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_22 = _RANDOM[10'h2BF][15];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_23 = _RANDOM[10'h2BF][16];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_24 = _RANDOM[10'h2BF][17];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_25 = _RANDOM[10'h2BF][18];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_26 = _RANDOM[10'h2BF][19];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_27 = _RANDOM[10'h2BF][20];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_28 = _RANDOM[10'h2BF][21];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_29 = _RANDOM[10'h2BF][22];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_30 = _RANDOM[10'h2BF][23];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_31 = _RANDOM[10'h2BF][24];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_32 = _RANDOM[10'h2BF][25];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_33 = _RANDOM[10'h2BF][26];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_34 = _RANDOM[10'h2BF][27];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_35 = _RANDOM[10'h2BF][28];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_36 = _RANDOM[10'h2BF][29];	// lsu.scala:1131:58, :1165:56
        io_dmem_s1_kill_0_REG_37 = _RANDOM[10'h2BF][30];	// lsu.scala:1131:58, :1153:56
        io_dmem_s1_kill_0_REG_38 = _RANDOM[10'h2BF][31];	// lsu.scala:1131:58, :1159:56
        io_dmem_s1_kill_0_REG_39 = _RANDOM[10'h2C0][0];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_40 = _RANDOM[10'h2C0][1];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_41 = _RANDOM[10'h2C0][2];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_42 = _RANDOM[10'h2C0][3];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_43 = _RANDOM[10'h2C0][4];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_44 = _RANDOM[10'h2C0][5];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_45 = _RANDOM[10'h2C0][6];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_46 = _RANDOM[10'h2C0][7];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_47 = _RANDOM[10'h2C0][8];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_48 = _RANDOM[10'h2C0][9];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_49 = _RANDOM[10'h2C0][10];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_50 = _RANDOM[10'h2C0][11];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_51 = _RANDOM[10'h2C0][12];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_52 = _RANDOM[10'h2C0][13];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_53 = _RANDOM[10'h2C0][14];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_54 = _RANDOM[10'h2C0][15];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_55 = _RANDOM[10'h2C0][16];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_56 = _RANDOM[10'h2C0][17];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_57 = _RANDOM[10'h2C0][18];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_58 = _RANDOM[10'h2C0][19];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_59 = _RANDOM[10'h2C0][20];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_60 = _RANDOM[10'h2C0][21];	// lsu.scala:1165:56
        io_dmem_s1_kill_0_REG_61 = _RANDOM[10'h2C0][22];	// lsu.scala:1153:56, :1165:56
        io_dmem_s1_kill_0_REG_62 = _RANDOM[10'h2C0][23];	// lsu.scala:1159:56, :1165:56
        io_dmem_s1_kill_0_REG_63 = _RANDOM[10'h2C0][24];	// lsu.scala:1165:56
        REG_1 = _RANDOM[10'h2C0][25];	// lsu.scala:1165:56, :1189:64
        REG_2 = _RANDOM[10'h2C0][26];	// lsu.scala:1165:56, :1199:18
        store_blocked_counter = _RANDOM[10'h2C0][30:27];	// lsu.scala:1165:56, :1204:36
        r_xcpt_valid = _RANDOM[10'h2C1][6];	// lsu.scala:1235:29
        r_xcpt_uop_br_mask = _RANDOM[10'h2C6][14:3];	// lsu.scala:1236:25
        r_xcpt_uop_rob_idx = _RANDOM[10'h2C8][5:0];	// lsu.scala:1236:25
        r_xcpt_cause = _RANDOM[10'h2CD][30:26];	// lsu.scala:1236:25
        r_xcpt_badvaddr = {_RANDOM[10'h2CD][31], _RANDOM[10'h2CE], _RANDOM[10'h2CF][6:0]};	// lsu.scala:1236:25
        io_core_ld_miss_REG = _RANDOM[10'h2CF][7];	// lsu.scala:1236:25, :1380:37
        spec_ld_succeed_REG = _RANDOM[10'h2CF][8];	// lsu.scala:1236:25, :1382:13
        spec_ld_succeed_REG_1 = _RANDOM[10'h2CF][12:9];	// lsu.scala:1236:25, :1384:56
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  NBDTLB_2 dtlb (	// lsu.scala:249:20
    .clock                        (clock),
    .reset                        (reset),
    .io_req_0_valid               (~_will_fire_store_commit_0_T_2),	// lsu.scala:538:31, :576:25
    .io_req_0_bits_vaddr          (exe_tlb_vaddr_0),	// lsu.scala:607:24
    .io_req_0_bits_passthrough    (will_fire_hella_incoming_0 & hella_req_phys),	// lsu.scala:243:34, :535:65, :643:23
    .io_req_0_bits_size
      (_exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0 | will_fire_load_retry_0
       | will_fire_sta_retry_0
         ? exe_tlb_uop_0_mem_size
         : will_fire_hella_incoming_0 ? hella_req_size : 2'h0),	// lsu.scala:243:34, :535:65, :536:61, :567:63, :597:24, :624:23, :628:52, :630:23
    .io_req_0_bits_cmd
      (_exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0 | will_fire_load_retry_0
       | will_fire_sta_retry_0
         ? exe_tlb_uop_0_mem_cmd
         : will_fire_hella_incoming_0 ? hella_req_cmd : 5'h0),	// lsu.scala:243:34, :535:65, :536:61, :567:63, :597:24, :633:23, :637:52, :639:23
    .io_sfence_valid
      (will_fire_sfence_0 & io_core_exe_0_req_bits_sfence_valid),	// lsu.scala:536:61, :618:32, :619:18
    .io_sfence_bits_rs1
      (will_fire_sfence_0 & io_core_exe_0_req_bits_sfence_bits_rs1),	// lsu.scala:536:61, :618:32, :619:18
    .io_sfence_bits_rs2
      (will_fire_sfence_0 & io_core_exe_0_req_bits_sfence_bits_rs2),	// lsu.scala:536:61, :618:32, :619:18
    .io_sfence_bits_addr
      (will_fire_sfence_0 ? io_core_exe_0_req_bits_sfence_bits_addr : 39'h0),	// lsu.scala:536:61, :616:43, :618:32, :619:18
    .io_ptw_req_ready             (io_ptw_req_ready),
    .io_ptw_resp_valid            (io_ptw_resp_valid),
    .io_ptw_resp_bits_ae          (io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn     (io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d       (io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a       (io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g       (io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u       (io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x       (io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w       (io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r       (io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v       (io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level       (io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous (io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode             (io_ptw_ptbr_mode),
    .io_ptw_status_dprv           (io_ptw_status_dprv),
    .io_ptw_status_mxr            (io_ptw_status_mxr),
    .io_ptw_status_sum            (io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l           (io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a           (io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x           (io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w           (io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r           (io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr            (io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask            (io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l           (io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a           (io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x           (io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w           (io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r           (io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr            (io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask            (io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l           (io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a           (io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x           (io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w           (io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r           (io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr            (io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask            (io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l           (io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a           (io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x           (io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w           (io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r           (io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr            (io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask            (io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l           (io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a           (io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x           (io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w           (io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r           (io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr            (io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask            (io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l           (io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a           (io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x           (io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w           (io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r           (io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr            (io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask            (io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l           (io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a           (io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x           (io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w           (io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r           (io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr            (io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask            (io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l           (io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a           (io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x           (io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w           (io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r           (io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr            (io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask            (io_ptw_pmp_7_mask),
    .io_kill                      (will_fire_hella_incoming_0 & io_hellacache_s1_kill),	// lsu.scala:535:65, :646:23
    .io_miss_rdy                  (_dtlb_io_miss_rdy),
    .io_resp_0_miss               (_dtlb_io_resp_0_miss),
    .io_resp_0_paddr              (_dtlb_io_resp_0_paddr),
    .io_resp_0_pf_ld              (_dtlb_io_resp_0_pf_ld),
    .io_resp_0_pf_st              (_dtlb_io_resp_0_pf_st),
    .io_resp_0_ae_ld              (_dtlb_io_resp_0_ae_ld),
    .io_resp_0_ae_st              (_dtlb_io_resp_0_ae_st),
    .io_resp_0_ma_ld              (_dtlb_io_resp_0_ma_ld),
    .io_resp_0_ma_st              (_dtlb_io_resp_0_ma_st),
    .io_resp_0_cacheable          (_dtlb_io_resp_0_cacheable),
    .io_ptw_req_valid             (_dtlb_io_ptw_req_valid),
    .io_ptw_req_bits_valid        (io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr    (io_ptw_req_bits_bits_addr)
  );
  ForwardingAgeLogic_3 forwarding_age_logic_0 (	// lsu.scala:1178:57
    .io_addr_matches
      ({ldst_addr_matches_0_15,
        ldst_addr_matches_0_14,
        ldst_addr_matches_0_13,
        ldst_addr_matches_0_12,
        ldst_addr_matches_0_11,
        ldst_addr_matches_0_10,
        ldst_addr_matches_0_9,
        ldst_addr_matches_0_8,
        ldst_addr_matches_0_7,
        ldst_addr_matches_0_6,
        ldst_addr_matches_0_5,
        ldst_addr_matches_0_4,
        ldst_addr_matches_0_3,
        ldst_addr_matches_0_2,
        ldst_addr_matches_0_1,
        ldst_addr_matches_0_0}),	// lsu.scala:1148:72, :1150:9, :1180:72
    .io_youngest_st_idx
      (do_st_search_0
         ? (_lcam_stq_idx_T
              ? mem_stq_incoming_e_0_bits_uop_stq_idx
              : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_stq_idx : 4'h0)
         : do_ld_search_0
             ? (fired_load_incoming_REG
                  ? mem_ldq_incoming_e_0_bits_uop_stq_idx
                  : fired_load_retry_REG
                      ? mem_ldq_retry_e_bits_uop_stq_idx
                      : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_uop_stq_idx : 4'h0)
             : 4'h0),	// lsu.scala:894:51, :901:51, :902:51, :904:51, :909:37, :910:37, :911:37, :912:37, :913:37, :915:33, :916:33, :917:33, :919:{33,57}, :921:33, :1014:108, :1016:106, :1029:37, :1030:37
    .io_forwarding_idx  (_forwarding_age_logic_0_io_forwarding_idx)
  );
  assign io_ptw_req_valid = _dtlb_io_ptw_req_valid;	// lsu.scala:249:20
  assign io_core_exe_0_iresp_valid = _io_core_exe_0_iresp_valid_output;	// lsu.scala:1306:5, :1344:5, :1348:5
  assign io_core_exe_0_iresp_bits_uop_rob_idx =
    _GEN_604
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_140[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_36[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_593;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_pdst =
    _GEN_604
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_145[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_40[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_594;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_is_amo =
    _GEN_604
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_163[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_61[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_597;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_uses_stq =
    _GEN_604
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_166[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_64[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_598;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_uop_dst_rtype =
    _GEN_604
      ? (io_dmem_resp_0_bits_uop_uses_ldq
           ? _GEN_177[io_dmem_resp_0_bits_uop_ldq_idx]
           : _GEN_74[io_dmem_resp_0_bits_uop_stq_idx])
      : _GEN_599;	// lsu.scala:224:42, :465:79, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_iresp_bits_data =
    _GEN_604
      ? io_dmem_resp_0_bits_data
      : {_ldq_bits_debug_wb_data_T_17
           ? {56{_GEN_596 & io_core_exe_0_iresp_bits_data_lo_2[7]}}
           : {_ldq_bits_debug_wb_data_T_9
                ? {48{_GEN_596 & io_core_exe_0_iresp_bits_data_lo_1[15]}}
                : {_ldq_bits_debug_wb_data_T_1
                     ? {32{_GEN_596 & io_core_exe_0_iresp_bits_data_lo[31]}}
                     : _GEN_603[63:32],
                   io_core_exe_0_iresp_bits_data_lo[31:16]},
              io_core_exe_0_iresp_bits_data_lo_1[15:8]},
         io_core_exe_0_iresp_bits_data_lo_2};	// AMOALU.scala:26:13, :39:{24,37}, :42:{20,26,76,85,98}, Bitwise.scala:72:12, Cat.scala:30:58, lsu.scala:1306:5, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_valid = _io_core_exe_0_fresp_valid_output;	// lsu.scala:1306:5, :1344:5, :1348:5
  assign io_core_exe_0_fresp_bits_uop_uopc =
    _GEN_604 ? _GEN_108[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_108[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_br_mask =
    _GEN_604 ? _GEN_102[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_592;	// lsu.scala:264:49, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_rob_idx =
    _GEN_604 ? _GEN_140[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_593;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_stq_idx =
    _GEN_604 ? _GEN_103[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_103[wb_forward_ldq_idx_0];	// lsu.scala:264:49, :1065:36, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_pdst =
    _GEN_604 ? _GEN_145[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_594;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_mem_size =
    _GEN_604 ? _GEN_104[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_595;	// lsu.scala:264:49, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_is_amo =
    _GEN_604 ? _GEN_163[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_597;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_uses_stq =
    _GEN_604 ? _GEN_166[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_598;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_dst_rtype =
    _GEN_604 ? _GEN_177[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_599;	// lsu.scala:465:79, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_uop_fp_val =
    _GEN_604 ? _GEN_181[io_dmem_resp_0_bits_uop_ldq_idx] : _GEN_181[wb_forward_ldq_idx_0];	// lsu.scala:465:79, :1065:36, :1306:5, :1311:58, :1344:5, :1348:5, util.scala:118:51
  assign io_core_exe_0_fresp_bits_data =
    {1'h0,
     _GEN_604
       ? io_dmem_resp_0_bits_data
       : {_ldq_bits_debug_wb_data_T_17
            ? {56{_GEN_596 & io_core_exe_0_fresp_bits_data_lo_2[7]}}
            : {_ldq_bits_debug_wb_data_T_9
                 ? {48{_GEN_596 & io_core_exe_0_fresp_bits_data_lo_1[15]}}
                 : {_ldq_bits_debug_wb_data_T_1
                      ? {32{_GEN_596 & io_core_exe_0_fresp_bits_data_lo[31]}}
                      : _GEN_603[63:32],
                    io_core_exe_0_fresp_bits_data_lo[31:16]},
               io_core_exe_0_fresp_bits_data_lo_1[15:8]},
          io_core_exe_0_fresp_bits_data_lo_2}};	// AMOALU.scala:26:13, :39:{24,37}, :42:{20,26,76,85,98}, Bitwise.scala:72:12, lsu.scala:249:20, :708:86, :1306:5, :1344:5, :1348:5, :1367:38, util.scala:118:51
  assign io_core_dis_ldq_idx_0 = ldq_tail;	// lsu.scala:216:29
  assign io_core_dis_ldq_idx_1 = _GEN_98;	// lsu.scala:333:21
  assign io_core_dis_stq_idx_0 = stq_tail;	// lsu.scala:218:29
  assign io_core_dis_stq_idx_1 = _GEN_99;	// lsu.scala:338:21
  assign io_core_ldq_full_0 = _GEN_95 == ldq_head;	// lsu.scala:215:29, :293:51, util.scala:203:14
  assign io_core_ldq_full_1 = _GEN_100 == ldq_head;	// lsu.scala:215:29, :293:51, util.scala:203:14
  assign io_core_stq_full_0 = _GEN_96 == stq_head;	// lsu.scala:217:29, :297:51, util.scala:203:14
  assign io_core_stq_full_1 = _GEN_101 == stq_head;	// lsu.scala:217:29, :297:51, util.scala:203:14
  assign io_core_fp_stdata_ready = _io_core_fp_stdata_ready_output;	// lsu.scala:866:61
  assign io_core_clr_bsy_0_valid =
    clr_bsy_valid_0 & (io_core_brupdate_b1_mispredict_mask & clr_bsy_brmask_0) == 12'h0
    & ~io_core_exception & ~io_core_clr_bsy_0_valid_REG & ~io_core_clr_bsy_0_valid_REG_2;	// lsu.scala:669:22, :930:32, :932:28, :979:{54,62,82,85,93}, util.scala:118:{51,59}
  assign io_core_clr_bsy_0_bits = clr_bsy_rob_idx_0;	// lsu.scala:931:28
  assign io_core_clr_bsy_1_valid =
    stdf_clr_bsy_valid
    & (io_core_brupdate_b1_mispredict_mask & stdf_clr_bsy_brmask) == 12'h0
    & ~io_core_exception & ~io_core_clr_bsy_1_valid_REG & ~io_core_clr_bsy_1_valid_REG_2;	// lsu.scala:669:22, :983:37, :985:33, :1004:{59,67,87,90,98}, util.scala:118:{51,59}
  assign io_core_clr_bsy_1_bits = stdf_clr_bsy_rob_idx;	// lsu.scala:984:33
  assign io_core_spec_ld_wakeup_0_valid = _io_core_spec_ld_wakeup_0_valid_output;	// lsu.scala:1260:69
  assign io_core_spec_ld_wakeup_0_bits = mem_incoming_uop_0_pdst;	// lsu.scala:908:37
  assign io_core_ld_miss =
    ~(~spec_ld_succeed_REG | _io_core_exe_0_iresp_valid_output
      & (_GEN_604
           ? (io_dmem_resp_0_bits_uop_uses_ldq
                ? _GEN_142[io_dmem_resp_0_bits_uop_ldq_idx]
                : _GEN_37[io_dmem_resp_0_bits_uop_stq_idx])
           : _GEN_142[wb_forward_ldq_idx_0]) == spec_ld_succeed_REG_1)
    & io_core_ld_miss_REG;	// lsu.scala:224:42, :465:79, :1065:36, :1306:5, :1308:7, :1311:58, :1314:40, :1328:7, :1330:62, :1344:5, :1348:5, :1380:{27,37}, :1382:{5,13,47}, :1383:33, :1384:{45,56}, :1387:26, :1388:21, util.scala:118:51
  assign io_core_fencei_rdy =
    ~(stq_0_valid | stq_1_valid | stq_2_valid | stq_3_valid | stq_4_valid | stq_5_valid
      | stq_6_valid | stq_7_valid | stq_8_valid | stq_9_valid | stq_10_valid
      | stq_11_valid | stq_12_valid | stq_13_valid | stq_14_valid | stq_15_valid)
    & io_dmem_ordered;	// lsu.scala:211:16, :286:79, :348:{28,42}
  assign io_core_lxcpt_valid =
    r_xcpt_valid & ~io_core_exception
    & (io_core_brupdate_b1_mispredict_mask & r_xcpt_uop_br_mask) == 12'h0;	// lsu.scala:669:22, :1235:29, :1236:25, :1253:61, util.scala:118:{51,59}
  assign io_core_lxcpt_bits_uop_br_mask = r_xcpt_uop_br_mask;	// lsu.scala:1236:25
  assign io_core_lxcpt_bits_uop_rob_idx = r_xcpt_uop_rob_idx;	// lsu.scala:1236:25
  assign io_core_lxcpt_bits_cause = r_xcpt_cause;	// lsu.scala:1236:25
  assign io_core_lxcpt_bits_badvaddr = r_xcpt_badvaddr;	// lsu.scala:1236:25
  assign io_core_perf_tlbMiss = io_ptw_req_ready & _dtlb_io_ptw_req_valid;	// Decoupled.scala:40:37, lsu.scala:249:20
  assign io_dmem_req_valid = dmem_req_0_valid;	// lsu.scala:766:39, :767:30, :773:43
  assign io_dmem_req_bits_0_valid = dmem_req_0_valid;	// lsu.scala:766:39, :767:30, :773:43
  assign io_dmem_req_bits_0_bits_uop_uopc =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_uopc
           : will_fire_load_retry_0
               ? _GEN_108[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_4[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_4[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_108[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_inst =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_inst
           : will_fire_load_retry_0
               ? _GEN_109[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_5[stq_retry_idx] : 32'h0)
      : will_fire_store_commit_0
          ? _GEN_5[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_109[ldq_wakeup_idx] : 32'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_inst =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_inst
           : will_fire_load_retry_0
               ? _GEN_110[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_6[stq_retry_idx] : 32'h0)
      : will_fire_store_commit_0
          ? _GEN_6[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_110[ldq_wakeup_idx] : 32'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_rvc =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_rvc
           : will_fire_load_retry_0
               ? _GEN_111[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_7[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_7[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_111[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_pc =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_pc
           : will_fire_load_retry_0
               ? _GEN_112[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_8[stq_retry_idx] : 40'h0)
      : will_fire_store_commit_0
          ? _GEN_8[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_112[ldq_wakeup_idx] : 40'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iq_type =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iq_type
           : will_fire_load_retry_0
               ? _GEN_113[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_9[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_9[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_113[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_fu_code =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_fu_code
           : will_fire_load_retry_0
               ? _GEN_114[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_10[stq_retry_idx] : 10'h0)
      : will_fire_store_commit_0
          ? _GEN_10[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_114[ldq_wakeup_idx] : 10'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_br_type =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_br_type
           : will_fire_load_retry_0
               ? _GEN_115[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_11[stq_retry_idx] : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_11[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_115[ldq_wakeup_idx] : 4'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_op1_sel =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_op1_sel
           : will_fire_load_retry_0
               ? _GEN_116[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_12[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_12[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_116[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_op2_sel =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_op2_sel
           : will_fire_load_retry_0
               ? _GEN_117[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_13[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_13[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_117[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_imm_sel =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_imm_sel
           : will_fire_load_retry_0
               ? _GEN_118[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_14[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_14[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_118[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_op_fcn =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_op_fcn
           : will_fire_load_retry_0
               ? _GEN_119[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_15[stq_retry_idx] : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_15[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_119[ldq_wakeup_idx] : 4'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_fcn_dw
           : will_fire_load_retry_0
               ? _GEN_120[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_16[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_16[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_120[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_csr_cmd
           : will_fire_load_retry_0
               ? _GEN_121[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_17[stq_retry_idx] : 3'h0)
      : will_fire_store_commit_0
          ? _GEN_17[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_121[ldq_wakeup_idx] : 3'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_load =
    _GEN_272
      ? exe_tlb_uop_0_ctrl_is_load
      : will_fire_store_commit_0
          ? _GEN_18[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_122[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_sta =
    _GEN_272
      ? exe_tlb_uop_0_ctrl_is_sta
      : will_fire_store_commit_0
          ? _GEN_19[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_123[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_std =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ctrl_is_std
           : will_fire_load_retry_0
               ? _GEN_124[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_20[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_20[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_124[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iw_state =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iw_state
           : will_fire_load_retry_0
               ? _GEN_125[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_21[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_21[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_125[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iw_p1_poisoned =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iw_p1_poisoned
           : will_fire_load_retry_0
               ? _GEN_126[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_22[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_22[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_126[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_iw_p2_poisoned =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_iw_p2_poisoned
           : will_fire_load_retry_0
               ? _GEN_127[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_23[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_23[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_127[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_br =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_br
           : will_fire_load_retry_0
               ? _GEN_128[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_24[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_24[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_128[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_jalr =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_jalr
           : will_fire_load_retry_0
               ? _GEN_129[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_25[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_25[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_129[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_jal =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_jal
           : will_fire_load_retry_0
               ? _GEN_130[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_26[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_26[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_130[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_sfb =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_sfb
           : will_fire_load_retry_0
               ? _GEN_131[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_27[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_27[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_131[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_br_mask =
    _GEN_272
      ? exe_tlb_uop_0_br_mask
      : will_fire_store_commit_0
          ? _GEN_28[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_201 : 12'h0;	// lsu.scala:220:29, :224:42, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_br_tag =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_br_tag
           : will_fire_load_retry_0
               ? _GEN_133[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_29[stq_retry_idx] : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_29[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_133[ldq_wakeup_idx] : 4'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ftq_idx =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ftq_idx
           : will_fire_load_retry_0
               ? _GEN_134[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_30[stq_retry_idx] : 5'h0)
      : will_fire_store_commit_0
          ? _GEN_30[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_134[ldq_wakeup_idx] : 5'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_edge_inst =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_edge_inst
           : will_fire_load_retry_0
               ? _GEN_135[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_31[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_31[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_135[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_pc_lob =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_pc_lob
           : will_fire_load_retry_0
               ? _GEN_136[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_32[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_32[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_136[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_taken =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_taken
           : will_fire_load_retry_0
               ? _GEN_137[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_33[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_33[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_137[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_imm_packed =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_imm_packed
           : will_fire_load_retry_0
               ? _GEN_138[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_34[stq_retry_idx] : 20'h0)
      : will_fire_store_commit_0
          ? _GEN_34[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_138[ldq_wakeup_idx] : 20'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_csr_addr =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_csr_addr
           : will_fire_load_retry_0
               ? _GEN_139[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_35[stq_retry_idx] : 12'h0)
      : will_fire_store_commit_0
          ? _GEN_35[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_139[ldq_wakeup_idx] : 12'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_rob_idx =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_rob_idx
           : will_fire_load_retry_0
               ? _GEN_141
               : will_fire_sta_retry_0 ? mem_stq_retry_e_out_bits_uop_rob_idx : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_36[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_140[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldq_idx =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldq_idx
           : will_fire_load_retry_0 ? _GEN_143 : will_fire_sta_retry_0 ? _GEN_198 : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_37[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_142[ldq_wakeup_idx] : 4'h0;	// lsu.scala:220:29, :224:42, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_stq_idx =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_stq_idx
           : will_fire_load_retry_0
               ? mem_ldq_retry_e_out_bits_uop_stq_idx
               : will_fire_sta_retry_0 ? mem_stq_retry_e_out_bits_uop_stq_idx : 4'h0)
      : will_fire_store_commit_0
          ? _GEN_38[stq_execute_head]
          : will_fire_load_wakeup_0 ? mem_ldq_wakeup_e_out_bits_uop_stq_idx : 4'h0;	// lsu.scala:220:29, :224:42, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_rxq_idx =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_rxq_idx
           : will_fire_load_retry_0
               ? _GEN_144[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_39[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_39[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_144[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_pdst =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_pdst
           : will_fire_load_retry_0 ? _GEN_146 : will_fire_sta_retry_0 ? _GEN_199 : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_40[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_145[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs1 =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs1
           : will_fire_load_retry_0
               ? _GEN_147[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_41[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_41[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_147[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs2 =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs2
           : will_fire_load_retry_0
               ? _GEN_148[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_42[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_42[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_148[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs3 =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs3
           : will_fire_load_retry_0
               ? _GEN_149[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_43[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_43[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_149[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ppred =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ppred
           : will_fire_load_retry_0
               ? _GEN_150[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_44[stq_retry_idx] : 5'h0)
      : will_fire_store_commit_0
          ? _GEN_44[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_150[ldq_wakeup_idx] : 5'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs1_busy =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs1_busy
           : will_fire_load_retry_0
               ? _GEN_151[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_45[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_45[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_151[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs2_busy =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs2_busy
           : will_fire_load_retry_0
               ? _GEN_152[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_46[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_46[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_152[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_prs3_busy =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_prs3_busy
           : will_fire_load_retry_0
               ? _GEN_153[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_47[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_47[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_153[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ppred_busy =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ppred_busy
           : will_fire_load_retry_0
               ? _GEN_154[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_48[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_48[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_154[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_stale_pdst =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_stale_pdst
           : will_fire_load_retry_0
               ? _GEN_155[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_49[stq_retry_idx] : 7'h0)
      : will_fire_store_commit_0
          ? _GEN_49[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_155[ldq_wakeup_idx] : 7'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_exception =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_exception
           : will_fire_load_retry_0
               ? _GEN_156[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_50[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_51
          : will_fire_load_wakeup_0 & _GEN_156[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_exc_cause =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_exc_cause
           : will_fire_load_retry_0
               ? _GEN_157[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_52[stq_retry_idx] : 64'h0)
      : will_fire_store_commit_0
          ? _GEN_52[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_157[ldq_wakeup_idx] : 64'h0;	// AMOALU.scala:26:13, lsu.scala:220:29, :224:42, :249:20, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_bypassable =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_bypassable
           : will_fire_load_retry_0
               ? _GEN_158[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_53[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_53[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_158[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_mem_cmd =
    _GEN_272
      ? exe_tlb_uop_0_mem_cmd
      : will_fire_store_commit_0
          ? _GEN_54[stq_execute_head]
          : will_fire_load_wakeup_0
              ? _GEN_159[ldq_wakeup_idx]
              : _GEN_277 ? hella_req_cmd : 5'h0;	// lsu.scala:220:29, :224:42, :243:34, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, :802:47, :811:39, :819:5, :827:39
  assign io_dmem_req_bits_0_bits_uop_mem_size =
    _GEN_272
      ? exe_tlb_uop_0_mem_size
      : will_fire_store_commit_0
          ? _GEN_56
          : will_fire_load_wakeup_0
              ? mem_ldq_wakeup_e_out_bits_uop_mem_size
              : _GEN_277 ? hella_req_size : 2'h0;	// lsu.scala:220:29, :224:42, :243:34, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, :802:47, :811:39, :812:39, :819:5, :827:39, :828:39
  assign io_dmem_req_bits_0_bits_uop_mem_signed =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_mem_signed
           : will_fire_load_retry_0
               ? _GEN_160[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_57[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_57[stq_execute_head]
          : will_fire_load_wakeup_0
              ? _GEN_160[ldq_wakeup_idx]
              : _GEN_277 & hella_req_signed;	// lsu.scala:220:29, :224:42, :243:34, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, :802:47, :811:39, :813:39, :819:5, :827:39, :829:39
  assign io_dmem_req_bits_0_bits_uop_is_fence =
    _GEN_272
      ? exe_tlb_uop_0_is_fence
      : will_fire_store_commit_0
          ? _GEN_59
          : will_fire_load_wakeup_0 & _GEN_161[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_fencei =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_fencei
           : will_fire_load_retry_0
               ? _GEN_162[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_60[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_60[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_162[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_amo =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_amo
           : will_fire_load_retry_0
               ? _GEN_163[ldq_retry_idx]
               : will_fire_sta_retry_0 & mem_stq_retry_e_out_bits_uop_is_amo)
      : will_fire_store_commit_0
          ? _GEN_62
          : will_fire_load_wakeup_0 & _GEN_163[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_uses_ldq =
    _GEN_272
      ? _mem_xcpt_uops_WIRE_0_uses_ldq
      : will_fire_store_commit_0
          ? _GEN_63[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_164[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_uses_stq =
    _GEN_272
      ? _mem_xcpt_uops_WIRE_0_uses_stq
      : will_fire_store_commit_0
          ? _GEN_64[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_166[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :430:31, :465:79, :502:88, :535:65, :597:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_sys_pc2epc =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_sys_pc2epc
           : will_fire_load_retry_0
               ? _GEN_168[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_65[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_65[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_168[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_is_unique =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_is_unique
           : will_fire_load_retry_0
               ? _GEN_169[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_66[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_66[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_169[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_flush_on_commit =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_flush_on_commit
           : will_fire_load_retry_0
               ? _GEN_170[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_67[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_67[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_170[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldst_is_rs1 =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldst_is_rs1
           : will_fire_load_retry_0
               ? _GEN_171[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_68[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_68[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_171[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldst =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldst
           : will_fire_load_retry_0
               ? _GEN_172[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_69[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_69[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_172[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs1 =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs1
           : will_fire_load_retry_0
               ? _GEN_173[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_70[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_70[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_173[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs2 =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs2
           : will_fire_load_retry_0
               ? _GEN_174[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_71[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_71[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_174[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs3 =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs3
           : will_fire_load_retry_0
               ? _GEN_175[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_72[stq_retry_idx] : 6'h0)
      : will_fire_store_commit_0
          ? _GEN_72[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_175[ldq_wakeup_idx] : 6'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_ldst_val =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_ldst_val
           : will_fire_load_retry_0
               ? _GEN_176[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_73[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_73[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_176[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_dst_rtype =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_dst_rtype
           : will_fire_load_retry_0
               ? _GEN_177[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_74[stq_retry_idx] : 2'h2)
      : will_fire_store_commit_0
          ? _GEN_74[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_177[ldq_wakeup_idx] : 2'h2;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30, util.scala:351:72
  assign io_dmem_req_bits_0_bits_uop_lrs1_rtype =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs1_rtype
           : will_fire_load_retry_0
               ? _GEN_178[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_75[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_75[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_178[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_lrs2_rtype =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_lrs2_rtype
           : will_fire_load_retry_0
               ? _GEN_179[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_76[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_76[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_179[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_frs3_en =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_frs3_en
           : will_fire_load_retry_0
               ? _GEN_180[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_77[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_77[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_180[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_fp_val =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_fp_val
           : will_fire_load_retry_0
               ? _GEN_181[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_78[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_78[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_181[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_fp_single =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_fp_single
           : will_fire_load_retry_0
               ? _GEN_182[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_79[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_79[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_182[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_xcpt_pf_if =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_xcpt_pf_if
           : will_fire_load_retry_0
               ? _GEN_183[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_80[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_80[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_183[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_xcpt_ae_if =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_xcpt_ae_if
           : will_fire_load_retry_0
               ? _GEN_184[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_81[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_81[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_184[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_xcpt_ma_if =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_xcpt_ma_if
           : will_fire_load_retry_0
               ? _GEN_185[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_82[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_82[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_185[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_bp_debug_if =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_bp_debug_if
           : will_fire_load_retry_0
               ? _GEN_186[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_83[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_83[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_186[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_bp_xcpt_if =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_bp_xcpt_if
           : will_fire_load_retry_0
               ? _GEN_187[ldq_retry_idx]
               : will_fire_sta_retry_0 & _GEN_84[stq_retry_idx])
      : will_fire_store_commit_0
          ? _GEN_84[stq_execute_head]
          : will_fire_load_wakeup_0 & _GEN_187[ldq_wakeup_idx];	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_fsrc =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_fsrc
           : will_fire_load_retry_0
               ? _GEN_188[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_85[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_85[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_188[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_uop_debug_tsrc =
    _GEN_272
      ? (_exe_tlb_uop_T_2
           ? io_core_exe_0_req_bits_uop_debug_tsrc
           : will_fire_load_retry_0
               ? _GEN_189[ldq_retry_idx]
               : will_fire_sta_retry_0 ? _GEN_86[stq_retry_idx] : 2'h0)
      : will_fire_store_commit_0
          ? _GEN_86[stq_execute_head]
          : will_fire_load_wakeup_0 ? _GEN_189[ldq_wakeup_idx] : 2'h0;	// lsu.scala:220:29, :224:42, :415:30, :422:30, :430:31, :465:79, :478:79, :502:88, :535:65, :536:61, :597:24, :599:53, :601:24, :602:24, :759:28, :766:39, :769:30, :773:43, :776:30, :780:45, :787:33, :794:44, :797:30
  assign io_dmem_req_bits_0_bits_addr =
    _GEN_275
      ? _GEN_270
      : will_fire_store_commit_0
          ? _GEN_89
          : will_fire_load_wakeup_0
              ? _GEN_202
              : will_fire_hella_incoming_0
                  ? _GEN_270
                  : will_fire_hella_wakeup_0 ? _GEN_274 : 40'h0;	// lsu.scala:224:42, :502:88, :535:65, :760:28, :766:39, :768:30, :773:43, :780:45, :782:33, :794:44, :796:30, :802:47, :806:39, :819:5, :822:39
  assign io_dmem_req_bits_0_bits_data =
    _GEN_272
      ? 64'h0
      : will_fire_store_commit_0
          ? _GEN_271[_GEN_56]
          : will_fire_load_wakeup_0 | will_fire_hella_incoming_0
            | ~will_fire_hella_wakeup_0
              ? 64'h0
              : _GEN_276[hella_req_size];	// AMOALU.scala:26:{13,19}, lsu.scala:220:29, :224:42, :243:34, :249:20, :535:65, :761:28, :766:39, :773:43, :780:45, :783:33, :794:44, :802:47, :807:39, :819:5
  assign io_dmem_req_bits_0_bits_is_hella =
    ~(_GEN_272 | will_fire_store_commit_0 | will_fire_load_wakeup_0)
    & (will_fire_hella_incoming_0 | will_fire_hella_wakeup_0);	// lsu.scala:220:29, :535:65, :762:31, :766:39, :773:43, :780:45, :794:44, :802:47, :814:39, :819:5
  assign io_dmem_s1_kill_0 =
    _GEN_565
      ? (_GEN_567
           ? io_dmem_s1_kill_0_REG_61
           : _GEN_568
               ? io_dmem_s1_kill_0_REG_62
               : _GEN_569 ? io_dmem_s1_kill_0_REG_63 : _GEN_563)
      : _GEN_563;	// lsu.scala:1148:{45,72}, :1149:106, :1150:9, :1153:{46,56}, :1156:60, :1157:9, :1159:{46,56}, :1162:37, :1163:9, :1165:{46,56}
  assign io_dmem_release_ready = will_fire_release_0;	// lsu.scala:534:63
  assign io_dmem_force_order = _GEN_636 & _GEN_637 | io_core_fence_dmem;	// lsu.scala:347:25, :1494:29, :1495:3, :1496:{43,64}, :1497:27
  assign io_hellacache_req_ready = ~(|hella_state);	// lsu.scala:242:38, :593:24, :1527:21
  assign io_hellacache_s2_nack = ~_GEN_639 & _GEN_638;	// lsu.scala:1524:27, :1527:34, :1533:38, :1550:{28,43}
  assign io_hellacache_resp_valid =
    ~(_GEN_639 | _GEN_638 | _GEN_640) & _GEN_571 & _GEN_641;	// lsu.scala:1288:28, :1524:27, :1526:28, :1527:34, :1533:38, :1550:{28,43}, :1553:{28,38}, :1560:40, :1562:35
  assign io_hellacache_s2_xcpt_ae_ld =
    ~(~(|hella_state) | _GEN_1 | _GEN_638) & _GEN_640 & hella_xcpt_ae_ld;	// lsu.scala:242:38, :246:34, :593:24, :803:26, :1525:27, :1527:{21,34}, :1533:38, :1550:{28,43}, :1553:{28,38}
endmodule

