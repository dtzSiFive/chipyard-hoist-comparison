// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module TLInterconnectCoupler_28(
  input         auto_tlserial_manager_crossing_out_a_ready,
                auto_tlserial_manager_crossing_out_d_valid,
  input  [2:0]  auto_tlserial_manager_crossing_out_d_bits_opcode,
  input  [1:0]  auto_tlserial_manager_crossing_out_d_bits_param,
  input  [2:0]  auto_tlserial_manager_crossing_out_d_bits_size,
  input  [3:0]  auto_tlserial_manager_crossing_out_d_bits_source,
  input         auto_tlserial_manager_crossing_out_d_bits_sink,
                auto_tlserial_manager_crossing_out_d_bits_denied,
  input  [63:0] auto_tlserial_manager_crossing_out_d_bits_data,
  input         auto_tlserial_manager_crossing_out_d_bits_corrupt,
                auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_opcode,
                auto_tl_in_a_bits_param,
                auto_tl_in_a_bits_size,
  input  [3:0]  auto_tl_in_a_bits_source,
  input  [28:0] auto_tl_in_a_bits_address,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input  [63:0] auto_tl_in_a_bits_data,
  input         auto_tl_in_a_bits_corrupt,
                auto_tl_in_d_ready,
  output        auto_tlserial_manager_crossing_out_a_valid,
  output [2:0]  auto_tlserial_manager_crossing_out_a_bits_opcode,
                auto_tlserial_manager_crossing_out_a_bits_param,
                auto_tlserial_manager_crossing_out_a_bits_size,
  output [3:0]  auto_tlserial_manager_crossing_out_a_bits_source,
  output [28:0] auto_tlserial_manager_crossing_out_a_bits_address,
  output [7:0]  auto_tlserial_manager_crossing_out_a_bits_mask,
  output [63:0] auto_tlserial_manager_crossing_out_a_bits_data,
  output        auto_tlserial_manager_crossing_out_a_bits_corrupt,
                auto_tlserial_manager_crossing_out_d_ready,
                auto_tl_in_a_ready,
                auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_opcode,
  output [1:0]  auto_tl_in_d_bits_param,
  output [2:0]  auto_tl_in_d_bits_size,
  output [3:0]  auto_tl_in_d_bits_source,
  output        auto_tl_in_d_bits_sink,
                auto_tl_in_d_bits_denied,
  output [63:0] auto_tl_in_d_bits_data,
  output        auto_tl_in_d_bits_corrupt
);

  wire        _widget_auto_out_a_valid;	// WidthWidget.scala:212:28
  wire [2:0]  _widget_auto_out_a_bits_opcode;	// WidthWidget.scala:212:28
  wire [2:0]  _widget_auto_out_a_bits_param;	// WidthWidget.scala:212:28
  wire [2:0]  _widget_auto_out_a_bits_size;	// WidthWidget.scala:212:28
  wire [3:0]  _widget_auto_out_a_bits_source;	// WidthWidget.scala:212:28
  wire [28:0] _widget_auto_out_a_bits_address;	// WidthWidget.scala:212:28
  wire [7:0]  _widget_auto_out_a_bits_mask;	// WidthWidget.scala:212:28
  wire [63:0] _widget_auto_out_a_bits_data;	// WidthWidget.scala:212:28
  wire        _widget_auto_out_a_bits_corrupt;	// WidthWidget.scala:212:28
  wire        _widget_auto_out_d_ready;	// WidthWidget.scala:212:28
  wire        _shrinker_auto_in_a_ready;	// SourceShrinker.scala:88:30
  wire        _shrinker_auto_in_d_valid;	// SourceShrinker.scala:88:30
  wire [2:0]  _shrinker_auto_in_d_bits_opcode;	// SourceShrinker.scala:88:30
  wire [1:0]  _shrinker_auto_in_d_bits_param;	// SourceShrinker.scala:88:30
  wire [2:0]  _shrinker_auto_in_d_bits_size;	// SourceShrinker.scala:88:30
  wire [3:0]  _shrinker_auto_in_d_bits_source;	// SourceShrinker.scala:88:30
  wire        _shrinker_auto_in_d_bits_sink;	// SourceShrinker.scala:88:30
  wire        _shrinker_auto_in_d_bits_denied;	// SourceShrinker.scala:88:30
  wire [63:0] _shrinker_auto_in_d_bits_data;	// SourceShrinker.scala:88:30
  wire        _shrinker_auto_in_d_bits_corrupt;	// SourceShrinker.scala:88:30
  TLSourceShrinker_1 shrinker (	// SourceShrinker.scala:88:30
    .auto_in_a_valid         (_widget_auto_out_a_valid),	// WidthWidget.scala:212:28
    .auto_in_a_bits_opcode   (_widget_auto_out_a_bits_opcode),	// WidthWidget.scala:212:28
    .auto_in_a_bits_param    (_widget_auto_out_a_bits_param),	// WidthWidget.scala:212:28
    .auto_in_a_bits_size     (_widget_auto_out_a_bits_size),	// WidthWidget.scala:212:28
    .auto_in_a_bits_source   (_widget_auto_out_a_bits_source),	// WidthWidget.scala:212:28
    .auto_in_a_bits_address  (_widget_auto_out_a_bits_address),	// WidthWidget.scala:212:28
    .auto_in_a_bits_mask     (_widget_auto_out_a_bits_mask),	// WidthWidget.scala:212:28
    .auto_in_a_bits_data     (_widget_auto_out_a_bits_data),	// WidthWidget.scala:212:28
    .auto_in_a_bits_corrupt  (_widget_auto_out_a_bits_corrupt),	// WidthWidget.scala:212:28
    .auto_in_d_ready         (_widget_auto_out_d_ready),	// WidthWidget.scala:212:28
    .auto_out_a_ready        (auto_tlserial_manager_crossing_out_a_ready),
    .auto_out_d_valid        (auto_tlserial_manager_crossing_out_d_valid),
    .auto_out_d_bits_opcode  (auto_tlserial_manager_crossing_out_d_bits_opcode),
    .auto_out_d_bits_param   (auto_tlserial_manager_crossing_out_d_bits_param),
    .auto_out_d_bits_size    (auto_tlserial_manager_crossing_out_d_bits_size),
    .auto_out_d_bits_source  (auto_tlserial_manager_crossing_out_d_bits_source),
    .auto_out_d_bits_sink    (auto_tlserial_manager_crossing_out_d_bits_sink),
    .auto_out_d_bits_denied  (auto_tlserial_manager_crossing_out_d_bits_denied),
    .auto_out_d_bits_data    (auto_tlserial_manager_crossing_out_d_bits_data),
    .auto_out_d_bits_corrupt (auto_tlserial_manager_crossing_out_d_bits_corrupt),
    .auto_in_a_ready         (_shrinker_auto_in_a_ready),
    .auto_in_d_valid         (_shrinker_auto_in_d_valid),
    .auto_in_d_bits_opcode   (_shrinker_auto_in_d_bits_opcode),
    .auto_in_d_bits_param    (_shrinker_auto_in_d_bits_param),
    .auto_in_d_bits_size     (_shrinker_auto_in_d_bits_size),
    .auto_in_d_bits_source   (_shrinker_auto_in_d_bits_source),
    .auto_in_d_bits_sink     (_shrinker_auto_in_d_bits_sink),
    .auto_in_d_bits_denied   (_shrinker_auto_in_d_bits_denied),
    .auto_in_d_bits_data     (_shrinker_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt  (_shrinker_auto_in_d_bits_corrupt),
    .auto_out_a_valid        (auto_tlserial_manager_crossing_out_a_valid),
    .auto_out_a_bits_opcode  (auto_tlserial_manager_crossing_out_a_bits_opcode),
    .auto_out_a_bits_param   (auto_tlserial_manager_crossing_out_a_bits_param),
    .auto_out_a_bits_size    (auto_tlserial_manager_crossing_out_a_bits_size),
    .auto_out_a_bits_source  (auto_tlserial_manager_crossing_out_a_bits_source),
    .auto_out_a_bits_address (auto_tlserial_manager_crossing_out_a_bits_address),
    .auto_out_a_bits_mask    (auto_tlserial_manager_crossing_out_a_bits_mask),
    .auto_out_a_bits_data    (auto_tlserial_manager_crossing_out_a_bits_data),
    .auto_out_a_bits_corrupt (auto_tlserial_manager_crossing_out_a_bits_corrupt),
    .auto_out_d_ready        (auto_tlserial_manager_crossing_out_d_ready)
  );
  TLWidthWidget_12 widget (	// WidthWidget.scala:212:28
    .auto_in_a_valid         (auto_tl_in_a_valid),
    .auto_in_a_bits_opcode   (auto_tl_in_a_bits_opcode),
    .auto_in_a_bits_param    (auto_tl_in_a_bits_param),
    .auto_in_a_bits_size     (auto_tl_in_a_bits_size),
    .auto_in_a_bits_source   (auto_tl_in_a_bits_source),
    .auto_in_a_bits_address  (auto_tl_in_a_bits_address),
    .auto_in_a_bits_mask     (auto_tl_in_a_bits_mask),
    .auto_in_a_bits_data     (auto_tl_in_a_bits_data),
    .auto_in_a_bits_corrupt  (auto_tl_in_a_bits_corrupt),
    .auto_in_d_ready         (auto_tl_in_d_ready),
    .auto_out_a_ready        (_shrinker_auto_in_a_ready),	// SourceShrinker.scala:88:30
    .auto_out_d_valid        (_shrinker_auto_in_d_valid),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_opcode  (_shrinker_auto_in_d_bits_opcode),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_param   (_shrinker_auto_in_d_bits_param),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_size    (_shrinker_auto_in_d_bits_size),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_source  (_shrinker_auto_in_d_bits_source),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_sink    (_shrinker_auto_in_d_bits_sink),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_denied  (_shrinker_auto_in_d_bits_denied),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_data    (_shrinker_auto_in_d_bits_data),	// SourceShrinker.scala:88:30
    .auto_out_d_bits_corrupt (_shrinker_auto_in_d_bits_corrupt),	// SourceShrinker.scala:88:30
    .auto_in_a_ready         (auto_tl_in_a_ready),
    .auto_in_d_valid         (auto_tl_in_d_valid),
    .auto_in_d_bits_opcode   (auto_tl_in_d_bits_opcode),
    .auto_in_d_bits_param    (auto_tl_in_d_bits_param),
    .auto_in_d_bits_size     (auto_tl_in_d_bits_size),
    .auto_in_d_bits_source   (auto_tl_in_d_bits_source),
    .auto_in_d_bits_sink     (auto_tl_in_d_bits_sink),
    .auto_in_d_bits_denied   (auto_tl_in_d_bits_denied),
    .auto_in_d_bits_data     (auto_tl_in_d_bits_data),
    .auto_in_d_bits_corrupt  (auto_tl_in_d_bits_corrupt),
    .auto_out_a_valid        (_widget_auto_out_a_valid),
    .auto_out_a_bits_opcode  (_widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_param   (_widget_auto_out_a_bits_param),
    .auto_out_a_bits_size    (_widget_auto_out_a_bits_size),
    .auto_out_a_bits_source  (_widget_auto_out_a_bits_source),
    .auto_out_a_bits_address (_widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask    (_widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data    (_widget_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt (_widget_auto_out_a_bits_corrupt),
    .auto_out_d_ready        (_widget_auto_out_d_ready)
  );
endmodule

