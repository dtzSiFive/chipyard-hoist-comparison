// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module TLROM(
  input         clock,
                reset,
                auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
                auto_in_a_bits_param,
  input  [1:0]  auto_in_a_bits_size,
  input  [11:0] auto_in_a_bits_source,
  input  [16:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_a_bits_corrupt,
                auto_in_d_ready,
  output        auto_in_a_ready,
                auto_in_d_valid,
  output [1:0]  auto_in_d_bits_size,
  output [11:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data
);

  wire [1023:0][63:0] _GEN =
    {64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h0,
     64'h73656D616E,
     64'h2D74757074756F2D,
     64'h6B636F6C6300736C,
     64'h6C65632D6B636F6C,
     64'h6323007374707572,
     64'h7265746E6900746E,
     64'h657261702D747075,
     64'h727265746E690073,
     64'h6B636F6C63007665,
     64'h646E2C7663736972,
     64'h797469726F6972,
     64'h702D78616D2C7663,
     64'h7369720068636174,
     64'h74612D6775626564,
     64'h6465646E657478,
     64'h652D737470757272,
     64'h65746E6900746E75,
     64'h6F632D7268736D2C,
     64'h6576696669730064,
     64'h656966696E752D65,
     64'h68636163006C6576,
     64'h656C2D6568636163,
     64'h73656D616E2D67,
     64'h6572007365676E61,
     64'h7200656C646E6168,
     64'h702C78756E696C00,
     64'h72656C6C6F72746E,
     64'h6F632D7470757272,
     64'h65746E6900736C6C,
     64'h65632D7470757272,
     64'h65746E6923007469,
     64'h6C70732D626C7400,
     64'h79636E6575716572,
     64'h662D65736162656D,
     64'h6974007375746174,
     64'h7300736E6F696765,
     64'h72706D702C766373,
     64'h6972007974697261,
     64'h6C756E617267706D,
     64'h702C766373697200,
     64'h6173692C76637369,
     64'h7200676572006568,
     64'h6361632D6C657665,
     64'h6C2D7478656E0065,
     64'h7079742D756D6D00,
     64'h657A69732D626C74,
     64'h2D6900737465732D,
     64'h626C742D6900657A,
     64'h69732D6568636163,
     64'h2D6900737465732D,
     64'h65686361632D6900,
     64'h657A69732D6B636F,
     64'h6C622D6568636163,
     64'h2D6900746E756F63,
     64'h2D746E696F706B61,
     64'h6572622D63657865,
     64'h2D65726177647261,
     64'h6800657079745F65,
     64'h636976656400657A,
     64'h69732D626C742D64,
     64'h737465732D626C,
     64'h742D6400657A6973,
     64'h2D65686361632D64,
     64'h737465732D6568,
     64'h6361632D6400657A,
     64'h69732D6B636F6C62,
     64'h2D65686361632D64,
     64'h79636E65757165,
     64'h72662D6B636F6C63,
     64'h306C6169726573,
     64'h6C65646F6D0065,
     64'h6C62697461706D6F,
     64'h6300736C6C65632D,
     64'h657A69732300736C,
     64'h6C65632D73736572,
     64'h6464612309000000,
     64'h200000002000000,
     64'h2000000006C6F72,
     64'h746E6F63A2010000,
     64'h800000003000000,
     64'h10000000001000,
     64'hF01000008000000,
     64'h300000000003030,
     64'h30303031406C7274,
     64'h632D74657365722D,
     64'h656C697401000000,
     64'h20000000B000000,
     64'h9301000004000000,
     64'h30000000B000000,
     64'h8D01000004000000,
     64'h3000000006B636F,
     64'h6C632D6465786966,
     64'h1B0000000C000000,
     64'h300000000000000,
     64'h6B636F6C635F7375,
     64'h62705F6D65747379,
     64'h7362757347020000,
     64'h1500000003000000,
     64'hE1F50534000000,
     64'h400000003000000,
     64'h3A020000,
     64'h400000003000000,
     64'h6B636F6C,
     64'h635F737562705F6D,
     64'h6574737973627573,
     64'h100000002000000,
     64'h6B636F6C632D64,
     64'h657869661B000000,
     64'hC00000003000000,
     64'h6B636F6C,
     64'h635F7375626D5F6D,
     64'h6574737973627573,
     64'h4702000015000000,
     64'h300000000E1F505,
     64'h3400000004000000,
     64'h300000000000000,
     64'h3A02000004000000,
     64'h300000000000000,
     64'h6B636F6C635F7375,
     64'h626D5F6D65747379,
     64'h7362757301000000,
     64'h2000000006C6F72,
     64'h746E6F63A2010000,
     64'h800000003000000,
     64'h10000000000054,
     64'hF01000008000000,
     64'h300000001000000,
     64'h2F02000004000000,
     64'h30000000C000000,
     64'h1E02000004000000,
     64'h300000000000000,
     64'h30747261752C6576,
     64'h696669731B000000,
     64'hD00000003000000,
     64'hB00000017020000,
     64'h400000003000000,
     64'h30303030303034,
     64'h35406C6169726573,
     64'h100000002000000,
     64'h6D656DA2010000,
     64'h400000003000000,
     64'h10000000100,
     64'hF01000008000000,
     64'h300000000306D6F,
     64'h722C657669666973,
     64'h1B0000000C000000,
     64'h300000000000030,
     64'h30303031406D6F72,
     64'h100000002000000,
     64'h400000093010000,
     64'h400000003000000,
     64'h40000008D010000,
     64'h400000003000000,
     64'h10000000200,
     64'hF01000008000000,
     64'h300000000303030,
     64'h3032406D6F722D66,
     64'h6977626C01000000,
     64'h200000003000000,
     64'h9301000004000000,
     64'h300000003000000,
     64'h8D01000004000000,
     64'h300000000100000,
     64'h100F010000,
     64'h800000003000000,
     64'h303030303030,
     64'h3031406D61722D66,
     64'h6977626C01000000,
     64'h20000000C000000,
     64'h9301000004000000,
     64'h30000000C000000,
     64'h8D01000004000000,
     64'h300000001000000,
     64'hC02000004000000,
     64'h300000001000000,
     64'hF901000004000000,
     64'h3000000006C6F72,
     64'h746E6F63A2010000,
     64'h800000003000000,
     64'h40000000C,
     64'hF01000008000000,
     64'h300000009000000,
     64'hA0000000B000000,
     64'hA00000009000000,
     64'h90000000B000000,
     64'h900000009000000,
     64'h80000000B000000,
     64'h80000000B000000,
     64'h700000009000000,
     64'h60000000B000000,
     64'h600000009000000,
     64'h50000000B000000,
     64'h5000000D8010000,
     64'h5800000003000000,
     64'h7801000000000000,
     64'h300000000306369,
     64'h6C702C7663736972,
     64'h1B0000000C000000,
     64'h300000001000000,
     64'h6701000004000000,
     64'h300000000000000,
     64'h3030303030306340,
     64'h72656C6C6F72746E,
     64'h6F632D7470757272,
     64'h65746E6901000000,
     64'h200000000100000,
     64'h3000000F010000,
     64'h800000003000000,
     64'h30726F7272,
     64'h652C657669666973,
     64'h1B0000000E000000,
     64'h300000000000030,
     64'h3030334065636976,
     64'h65642D726F727265,
     64'h100000002000000,
     64'h6C6F72746E6F63,
     64'hA201000008000000,
     64'h300000000100000,
     64'hF010000,
     64'h800000003000000,
     64'hFFFF00000A000000,
     64'hFFFF000009000000,
     64'hFFFF000008000000,
     64'hFFFF000007000000,
     64'hFFFF000006000000,
     64'hFFFF000005000000,
     64'hD801000030000000,
     64'h300000000000000,
     64'h6761746AEC010000,
     64'h500000003000000,
     64'h3331302D,
     64'h67756265642C7663,
     64'h736972003331302D,
     64'h67756265642C6576,
     64'h696669731B000000,
     64'h2100000003000000,
     64'h304072656C6C,
     64'h6F72746E6F632D67,
     64'h7562656401000000,
     64'h2000000006C6F72,
     64'h746E6F63A2010000,
     64'h800000003000000,
     64'h10000000002,
     64'hF01000008000000,
     64'h300000007000000,
     64'hA00000003000000,
     64'hA00000007000000,
     64'h900000003000000,
     64'h900000007000000,
     64'h800000003000000,
     64'h800000007000000,
     64'h700000003000000,
     64'h700000007000000,
     64'h600000003000000,
     64'h600000007000000,
     64'h500000003000000,
     64'h5000000D8010000,
     64'h6000000003000000,
     64'h30746E69,
     64'h6C632C7663736972,
     64'h1B0000000D000000,
     64'h300000000000030,
     64'h3030303030324074,
     64'h6E696C6301000000,
     64'h200000001000000,
     64'h9301000004000000,
     64'h300000001000000,
     64'h8D01000004000000,
     64'h300000007000000,
     64'hC601000004000000,
     64'h3000000006C6F72,
     64'h746E6F63A2010000,
     64'h800000003000000,
     64'h10000000000102,
     64'hF01000008000000,
     64'h300000004000000,
     64'h300000002000000,
     64'hFE0000000C000000,
     64'h300000000000000,
     64'h6568636163003065,
     64'h6863616365766973,
     64'h756C636E692C6576,
     64'h696669731B000000,
     64'h1D00000003000000,
     64'hB801000000000000,
     64'h300000000000800,
     64'h6600000004000000,
     64'h300000000040000,
     64'h5900000004000000,
     64'h300000002000000,
     64'hAC01000004000000,
     64'h300000040000000,
     64'h4600000004000000,
     64'h300000000000000,
     64'h3030303031303240,
     64'h72656C6C6F72746E,
     64'h6F632D6568636163,
     64'h100000002000000,
     64'h6C6F72746E6F63,
     64'hA201000008000000,
     64'h300000000100000,
     64'h4000000F010000,
     64'h800000003000000,
     64'h3030303440,
     64'h6765722D73736572,
     64'h6464612D746F6F62,
     64'h10000009B010000,
     64'h3000000,
     64'h7375622D656C70,
     64'h6D697300636F732D,
     64'h6E776F6E6B6E752D,
     64'h7069686374656B63,
     64'h6F722C7370696863,
     64'h656572661B000000,
     64'h2C00000003000000,
     64'h10000000F000000,
     64'h400000003000000,
     64'h100000000000000,
     64'h400000003000000,
     64'h636F7301000000,
     64'h200000002000000,
     64'h9301000004000000,
     64'h300000002000000,
     64'h8D01000004000000,
     64'h300000000000010,
     64'h800F010000,
     64'h800000003000000,
     64'h79726F6D656D,
     64'h8700000007000000,
     64'h300000000303030,
     64'h3030303038407972,
     64'h6F6D656D01000000,
     64'h200000000000030,
     64'h666974682C626375,
     64'h1B0000000A000000,
     64'h300000000000000,
     64'h6669746801000000,
     64'h200000002000000,
     64'h20000000A000000,
     64'h9301000004000000,
     64'h30000000A000000,
     64'h8D01000004000000,
     64'h300000078010000,
     64'h3000000,
     64'h63746E692D75,
     64'h70632C7663736972,
     64'h1B0000000F000000,
     64'h300000001000000,
     64'h6701000004000000,
     64'h300000000000000,
     64'h72656C6C6F72746E,
     64'h6F632D7470757272,
     64'h65746E6901000000,
     64'h5D01000000000000,
     64'h300000040420F00,
     64'h4A01000004000000,
     64'h300000000000000,
     64'h79616B6F43010000,
     64'h500000003000000,
     64'h800000032010000,
     64'h400000003000000,
     64'h40000001D010000,
     64'h400000003000000,
     64'h636466616D69,
     64'h3436767213010000,
     64'hB00000003000000,
     64'h50000000F010000,
     64'h400000003000000,
     64'h1000000FE000000,
     64'h400000003000000,
     64'h393376732C76,
     64'h63736972F5000000,
     64'hB00000003000000,
     64'h20000000EA000000,
     64'h400000003000000,
     64'h1000000DF000000,
     64'h400000003000000,
     64'h400000D2000000,
     64'h400000003000000,
     64'h40000000C5000000,
     64'h400000003000000,
     64'h40000000B2000000,
     64'h400000003000000,
     64'h93000000,
     64'h400000003000000,
     64'h75706387000000,
     64'h400000003000000,
     64'h80000007C000000,
     64'h400000003000000,
     64'h100000071000000,
     64'h400000003000000,
     64'h40000064000000,
     64'h400000003000000,
     64'h4000000057000000,
     64'h400000003000000,
     64'h4000000044000000,
     64'h400000003000000,
     64'h76637369720030,
     64'h6D6F6F622C726162,
     64'h2D6263751B000000,
     64'h1400000003000000,
     64'h34000000,
     64'h400000003000000,
     64'h3540757063,
     64'h100000002000000,
     64'h200000009000000,
     64'h9301000004000000,
     64'h300000009000000,
     64'h8D01000004000000,
     64'h300000078010000,
     64'h3000000,
     64'h63746E692D75,
     64'h70632C7663736972,
     64'h1B0000000F000000,
     64'h300000001000000,
     64'h6701000004000000,
     64'h300000000000000,
     64'h72656C6C6F72746E,
     64'h6F632D7470757272,
     64'h65746E6901000000,
     64'h5D01000000000000,
     64'h300000040420F00,
     64'h4A01000004000000,
     64'h300000000000000,
     64'h79616B6F43010000,
     64'h500000003000000,
     64'h800000032010000,
     64'h400000003000000,
     64'h40000001D010000,
     64'h400000003000000,
     64'h636466616D69,
     64'h3436767213010000,
     64'hB00000003000000,
     64'h40000000F010000,
     64'h400000003000000,
     64'h1000000FE000000,
     64'h400000003000000,
     64'h393376732C76,
     64'h63736972F5000000,
     64'hB00000003000000,
     64'h20000000EA000000,
     64'h400000003000000,
     64'h1000000DF000000,
     64'h400000003000000,
     64'h800000D2000000,
     64'h400000003000000,
     64'h40000000C5000000,
     64'h400000003000000,
     64'h40000000B2000000,
     64'h400000003000000,
     64'h93000000,
     64'h400000003000000,
     64'h75706387000000,
     64'h400000003000000,
     64'h100000007C000000,
     64'h400000003000000,
     64'h100000071000000,
     64'h400000003000000,
     64'h80000064000000,
     64'h400000003000000,
     64'h4000000057000000,
     64'h400000003000000,
     64'h4000000044000000,
     64'h400000003000000,
     64'h76637369720030,
     64'h6D6F6F622C726162,
     64'h2D6263751B000000,
     64'h1400000003000000,
     64'h34000000,
     64'h400000003000000,
     64'h3440757063,
     64'h100000002000000,
     64'h200000008000000,
     64'h9301000004000000,
     64'h300000008000000,
     64'h8D01000004000000,
     64'h300000078010000,
     64'h3000000,
     64'h63746E692D75,
     64'h70632C7663736972,
     64'h1B0000000F000000,
     64'h300000001000000,
     64'h6701000004000000,
     64'h300000000000000,
     64'h72656C6C6F72746E,
     64'h6F632D7470757272,
     64'h65746E6901000000,
     64'h5D01000000000000,
     64'h300000040420F00,
     64'h4A01000004000000,
     64'h300000000000000,
     64'h79616B6F43010000,
     64'h500000003000000,
     64'h800000032010000,
     64'h400000003000000,
     64'h40000001D010000,
     64'h400000003000000,
     64'h636466616D69,
     64'h3436767213010000,
     64'hB00000003000000,
     64'h30000000F010000,
     64'h400000003000000,
     64'h1000000FE000000,
     64'h400000003000000,
     64'h393376732C76,
     64'h63736972F5000000,
     64'hB00000003000000,
     64'h20000000EA000000,
     64'h400000003000000,
     64'h1000000DF000000,
     64'h400000003000000,
     64'h800000D2000000,
     64'h400000003000000,
     64'h40000000C5000000,
     64'h400000003000000,
     64'h40000000B2000000,
     64'h400000003000000,
     64'h93000000,
     64'h400000003000000,
     64'h75706387000000,
     64'h400000003000000,
     64'h200000007C000000,
     64'h400000003000000,
     64'h100000071000000,
     64'h400000003000000,
     64'h80000064000000,
     64'h400000003000000,
     64'h4000000057000000,
     64'h400000003000000,
     64'h4000000044000000,
     64'h400000003000000,
     64'h76637369720030,
     64'h6D6F6F622C726162,
     64'h2D6263751B000000,
     64'h1400000003000000,
     64'h34000000,
     64'h400000003000000,
     64'h3340757063,
     64'h100000002000000,
     64'h200000007000000,
     64'h9301000004000000,
     64'h300000007000000,
     64'h8D01000004000000,
     64'h300000078010000,
     64'h3000000,
     64'h63746E692D75,
     64'h70632C7663736972,
     64'h1B0000000F000000,
     64'h300000001000000,
     64'h6701000004000000,
     64'h300000000000000,
     64'h72656C6C6F72746E,
     64'h6F632D7470757272,
     64'h65746E6901000000,
     64'h40420F004A010000,
     64'h400000003000000,
     64'h79616B6F,
     64'h4301000005000000,
     64'h300000008000000,
     64'h3201000004000000,
     64'h300000004000000,
     64'h1D01000004000000,
     64'h300000000000000,
     64'h63616D6934367672,
     64'h1301000009000000,
     64'h300000002000000,
     64'hF01000004000000,
     64'h300000001000000,
     64'hFE00000004000000,
     64'h300000000100000,
     64'hD200000004000000,
     64'h300000040000000,
     64'hC500000004000000,
     64'h300000040000000,
     64'hB200000004000000,
     64'h300000001000000,
     64'h9300000004000000,
     64'h300000000757063,
     64'h8700000004000000,
     64'h300000000100000,
     64'h6400000004000000,
     64'h300000040000000,
     64'h5700000004000000,
     64'h300000040000000,
     64'h4400000004000000,
     64'h300000000000000,
     64'h7663736972003074,
     64'h656B636F722C6576,
     64'h696669731B000000,
     64'h1500000003000000,
     64'h34000000,
     64'h400000003000000,
     64'h3240757063,
     64'h100000002000000,
     64'h200000006000000,
     64'h9301000004000000,
     64'h300000006000000,
     64'h8D01000004000000,
     64'h300000078010000,
     64'h3000000,
     64'h63746E692D75,
     64'h70632C7663736972,
     64'h1B0000000F000000,
     64'h300000001000000,
     64'h6701000004000000,
     64'h300000000000000,
     64'h72656C6C6F72746E,
     64'h6F632D7470757272,
     64'h65746E6901000000,
     64'h5D01000000000000,
     64'h300000040420F00,
     64'h4A01000004000000,
     64'h300000000000000,
     64'h79616B6F43010000,
     64'h500000003000000,
     64'h800000032010000,
     64'h400000003000000,
     64'h40000001D010000,
     64'h400000003000000,
     64'h63616D69,
     64'h3436767213010000,
     64'h900000003000000,
     64'h10000000F010000,
     64'h400000003000000,
     64'h1000000FE000000,
     64'h400000003000000,
     64'h393376732C76,
     64'h63736972F5000000,
     64'hB00000003000000,
     64'h4000000EA000000,
     64'h400000003000000,
     64'h1000000DF000000,
     64'h400000003000000,
     64'h100000D2000000,
     64'h400000003000000,
     64'h40000000C5000000,
     64'h400000003000000,
     64'h40000000B2000000,
     64'h400000003000000,
     64'h100000093000000,
     64'h400000003000000,
     64'h75706387000000,
     64'h400000003000000,
     64'h40000007C000000,
     64'h400000003000000,
     64'h100000071000000,
     64'h400000003000000,
     64'h10000064000000,
     64'h400000003000000,
     64'h4000000057000000,
     64'h400000003000000,
     64'h4000000044000000,
     64'h400000003000000,
     64'h76637369,
     64'h72003074656B636F,
     64'h722C657669666973,
     64'h1B00000015000000,
     64'h300000000000000,
     64'h3400000004000000,
     64'h300000000000031,
     64'h4075706301000000,
     64'h200000002000000,
     64'h500000093010000,
     64'h400000003000000,
     64'h50000008D010000,
     64'h400000003000000,
     64'h7801000000000000,
     64'h300000000006374,
     64'h6E692D7570632C76,
     64'h637369721B000000,
     64'hF00000003000000,
     64'h100000067010000,
     64'h400000003000000,
     64'h72656C6C,
     64'h6F72746E6F632D74,
     64'h7075727265746E69,
     64'h10000005D010000,
     64'h3000000,
     64'h40420F004A010000,
     64'h400000003000000,
     64'h79616B6F,
     64'h4301000005000000,
     64'h300000008000000,
     64'h3201000004000000,
     64'h300000004000000,
     64'h1D01000004000000,
     64'h300000000006364,
     64'h66616D6934367672,
     64'h130100000B000000,
     64'h300000000000000,
     64'hF01000004000000,
     64'h300000001000000,
     64'hFE00000004000000,
     64'h300000000003933,
     64'h76732C7663736972,
     64'hF50000000B000000,
     64'h300000020000000,
     64'hEA00000004000000,
     64'h300000001000000,
     64'hDF00000004000000,
     64'h300000000400000,
     64'hD200000004000000,
     64'h300000040000000,
     64'hC500000004000000,
     64'h300000040000000,
     64'hB200000004000000,
     64'h300000001000000,
     64'h9300000004000000,
     64'h300000000757063,
     64'h8700000004000000,
     64'h300000020000000,
     64'h7C00000004000000,
     64'h300000001000000,
     64'h7100000004000000,
     64'h300000000400000,
     64'h6400000004000000,
     64'h300000040000000,
     64'h5700000004000000,
     64'h300000040000000,
     64'h4400000004000000,
     64'h300000000000000,
     64'h7663736972003074,
     64'h656B636F722C6576,
     64'h696669731B000000,
     64'h1500000003000000,
     64'h34000000,
     64'h400000003000000,
     64'h3040757063,
     64'h100000000000000,
     64'hF00000004000000,
     64'h300000001000000,
     64'h4000000,
     64'h300000000000000,
     64'h7375706301000000,
     64'h200000000000000,
     64'h3030303030303435,
     64'h406C61697265732F,
     64'h636F732F2C000000,
     64'h1500000003000000,
     64'h73657361696C61,
     64'h100000000000000,
     64'h6E776F6E6B6E752D,
     64'h7069686374656B63,
     64'h6F722C7370696863,
     64'h6565726626000000,
     64'h1D00000003000000,
     64'h7665642D,
     64'h6E776F6E6B6E752D,
     64'h7069686374656B63,
     64'h6F722C7370696863,
     64'h656572661B000000,
     64'h2100000003000000,
     64'h10000000F000000,
     64'h400000003000000,
     64'h100000000000000,
     64'h400000003000000,
     64'h1000000,
     64'h0,
     64'h0,
     64'h4C1500005A020000,
     64'h10000000,
     64'h1100000028000000,
     64'h8415000038000000,
     64'hDE170000EDFE0DD0,
     64'h1330200073,
     64'h3006307308000613,
     64'h185859300000597,
     64'hF140257334151073,
     64'h5650300004537,
     64'h5A02300B505B3,
     64'h251513FE029EE3,
     64'h5A283FFDFF06F,
     64'h1050007330052073,
     64'h3045107300800513,
     64'h3030107300028463,
     64'h12F2934122D293,
     64'h301022F330551073,
     64'hFC05051300000517,
     64'h0,
     64'h0,
     64'h5C0006F,
     64'hFE069AE3FFC62683,
     64'h46061300D62023,
     64'h10069300458613,
     64'h680006F00050463,
     64'hF1402573020005B7};	// BootROM.scala:51:47
  TLMonitor_77 monitor (	// Nodes.scala:24:25
    .clock                (clock),
    .reset                (reset),
    .io_in_a_ready        (auto_in_d_ready),
    .io_in_a_valid        (auto_in_a_valid),
    .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
    .io_in_a_bits_param   (auto_in_a_bits_param),
    .io_in_a_bits_size    (auto_in_a_bits_size),
    .io_in_a_bits_source  (auto_in_a_bits_source),
    .io_in_a_bits_address (auto_in_a_bits_address),
    .io_in_a_bits_mask    (auto_in_a_bits_mask),
    .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
    .io_in_d_ready        (auto_in_d_ready),
    .io_in_d_valid        (auto_in_a_valid),
    .io_in_d_bits_size    (auto_in_a_bits_size),
    .io_in_d_bits_source  (auto_in_a_bits_source)
  );
  assign auto_in_a_ready = auto_in_d_ready;
  assign auto_in_d_valid = auto_in_a_valid;
  assign auto_in_d_bits_size = auto_in_a_bits_size;
  assign auto_in_d_bits_source = auto_in_a_bits_source;
  assign auto_in_d_bits_data =
    (|(auto_in_a_bits_address[15:13])) ? 64'h0 : _GEN[auto_in_a_bits_address[12:3]];	// BootROM.scala:44:18, :49:34, :50:68, :51:{47,53}
endmodule

