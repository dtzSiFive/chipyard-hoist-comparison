// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module FetchBuffer_1(
  input         clock,
                reset,
                io_enq_valid,
  input  [39:0] io_enq_bits_pc,
  input         io_enq_bits_edge_inst_0,
                io_enq_bits_edge_inst_1,
  input  [31:0] io_enq_bits_insts_0,
                io_enq_bits_insts_1,
                io_enq_bits_insts_2,
                io_enq_bits_insts_3,
                io_enq_bits_insts_4,
                io_enq_bits_insts_5,
                io_enq_bits_insts_6,
                io_enq_bits_insts_7,
                io_enq_bits_exp_insts_0,
                io_enq_bits_exp_insts_1,
                io_enq_bits_exp_insts_2,
                io_enq_bits_exp_insts_3,
                io_enq_bits_exp_insts_4,
                io_enq_bits_exp_insts_5,
                io_enq_bits_exp_insts_6,
                io_enq_bits_exp_insts_7,
  input         io_enq_bits_shadowed_mask_0,
                io_enq_bits_shadowed_mask_1,
                io_enq_bits_shadowed_mask_2,
                io_enq_bits_shadowed_mask_3,
                io_enq_bits_shadowed_mask_4,
                io_enq_bits_shadowed_mask_5,
                io_enq_bits_shadowed_mask_6,
                io_enq_bits_shadowed_mask_7,
                io_enq_bits_cfi_idx_valid,
  input  [2:0]  io_enq_bits_cfi_idx_bits,
  input  [4:0]  io_enq_bits_ftq_idx,
  input  [7:0]  io_enq_bits_mask,
  input         io_enq_bits_xcpt_pf_if,
                io_enq_bits_xcpt_ae_if,
                io_enq_bits_bp_debug_if_oh_0,
                io_enq_bits_bp_debug_if_oh_1,
                io_enq_bits_bp_debug_if_oh_2,
                io_enq_bits_bp_debug_if_oh_3,
                io_enq_bits_bp_debug_if_oh_4,
                io_enq_bits_bp_debug_if_oh_5,
                io_enq_bits_bp_debug_if_oh_6,
                io_enq_bits_bp_debug_if_oh_7,
                io_enq_bits_bp_xcpt_if_oh_0,
                io_enq_bits_bp_xcpt_if_oh_1,
                io_enq_bits_bp_xcpt_if_oh_2,
                io_enq_bits_bp_xcpt_if_oh_3,
                io_enq_bits_bp_xcpt_if_oh_4,
                io_enq_bits_bp_xcpt_if_oh_5,
                io_enq_bits_bp_xcpt_if_oh_6,
                io_enq_bits_bp_xcpt_if_oh_7,
  input  [1:0]  io_enq_bits_fsrc,
  input         io_deq_ready,
                io_clear,
  output        io_enq_ready,
                io_deq_valid,
                io_deq_bits_uops_0_valid,
  output [31:0] io_deq_bits_uops_0_bits_inst,
                io_deq_bits_uops_0_bits_debug_inst,
  output        io_deq_bits_uops_0_bits_is_rvc,
  output [39:0] io_deq_bits_uops_0_bits_debug_pc,
  output [3:0]  io_deq_bits_uops_0_bits_ctrl_br_type,
  output [1:0]  io_deq_bits_uops_0_bits_ctrl_op1_sel,
  output [2:0]  io_deq_bits_uops_0_bits_ctrl_op2_sel,
                io_deq_bits_uops_0_bits_ctrl_imm_sel,
  output [3:0]  io_deq_bits_uops_0_bits_ctrl_op_fcn,
  output        io_deq_bits_uops_0_bits_ctrl_fcn_dw,
  output [2:0]  io_deq_bits_uops_0_bits_ctrl_csr_cmd,
  output        io_deq_bits_uops_0_bits_ctrl_is_load,
                io_deq_bits_uops_0_bits_ctrl_is_sta,
                io_deq_bits_uops_0_bits_ctrl_is_std,
  output [1:0]  io_deq_bits_uops_0_bits_iw_state,
  output        io_deq_bits_uops_0_bits_iw_p1_poisoned,
                io_deq_bits_uops_0_bits_iw_p2_poisoned,
                io_deq_bits_uops_0_bits_is_sfb,
  output [4:0]  io_deq_bits_uops_0_bits_ftq_idx,
  output        io_deq_bits_uops_0_bits_edge_inst,
  output [5:0]  io_deq_bits_uops_0_bits_pc_lob,
  output        io_deq_bits_uops_0_bits_taken,
  output [11:0] io_deq_bits_uops_0_bits_csr_addr,
  output [1:0]  io_deq_bits_uops_0_bits_rxq_idx,
  output        io_deq_bits_uops_0_bits_xcpt_pf_if,
                io_deq_bits_uops_0_bits_xcpt_ae_if,
                io_deq_bits_uops_0_bits_xcpt_ma_if,
                io_deq_bits_uops_0_bits_bp_debug_if,
                io_deq_bits_uops_0_bits_bp_xcpt_if,
  output [1:0]  io_deq_bits_uops_0_bits_debug_fsrc,
                io_deq_bits_uops_0_bits_debug_tsrc,
  output        io_deq_bits_uops_1_valid,
  output [31:0] io_deq_bits_uops_1_bits_inst,
                io_deq_bits_uops_1_bits_debug_inst,
  output        io_deq_bits_uops_1_bits_is_rvc,
  output [39:0] io_deq_bits_uops_1_bits_debug_pc,
  output [3:0]  io_deq_bits_uops_1_bits_ctrl_br_type,
  output [1:0]  io_deq_bits_uops_1_bits_ctrl_op1_sel,
  output [2:0]  io_deq_bits_uops_1_bits_ctrl_op2_sel,
                io_deq_bits_uops_1_bits_ctrl_imm_sel,
  output [3:0]  io_deq_bits_uops_1_bits_ctrl_op_fcn,
  output        io_deq_bits_uops_1_bits_ctrl_fcn_dw,
  output [2:0]  io_deq_bits_uops_1_bits_ctrl_csr_cmd,
  output        io_deq_bits_uops_1_bits_ctrl_is_load,
                io_deq_bits_uops_1_bits_ctrl_is_sta,
                io_deq_bits_uops_1_bits_ctrl_is_std,
  output [1:0]  io_deq_bits_uops_1_bits_iw_state,
  output        io_deq_bits_uops_1_bits_iw_p1_poisoned,
                io_deq_bits_uops_1_bits_iw_p2_poisoned,
                io_deq_bits_uops_1_bits_is_sfb,
  output [4:0]  io_deq_bits_uops_1_bits_ftq_idx,
  output        io_deq_bits_uops_1_bits_edge_inst,
  output [5:0]  io_deq_bits_uops_1_bits_pc_lob,
  output        io_deq_bits_uops_1_bits_taken,
  output [11:0] io_deq_bits_uops_1_bits_csr_addr,
  output [1:0]  io_deq_bits_uops_1_bits_rxq_idx,
  output        io_deq_bits_uops_1_bits_xcpt_pf_if,
                io_deq_bits_uops_1_bits_xcpt_ae_if,
                io_deq_bits_uops_1_bits_xcpt_ma_if,
                io_deq_bits_uops_1_bits_bp_debug_if,
                io_deq_bits_uops_1_bits_bp_xcpt_if,
  output [1:0]  io_deq_bits_uops_1_bits_debug_fsrc,
                io_deq_bits_uops_1_bits_debug_tsrc,
  output        io_deq_bits_uops_2_valid,
  output [31:0] io_deq_bits_uops_2_bits_inst,
                io_deq_bits_uops_2_bits_debug_inst,
  output        io_deq_bits_uops_2_bits_is_rvc,
  output [39:0] io_deq_bits_uops_2_bits_debug_pc,
  output [3:0]  io_deq_bits_uops_2_bits_ctrl_br_type,
  output [1:0]  io_deq_bits_uops_2_bits_ctrl_op1_sel,
  output [2:0]  io_deq_bits_uops_2_bits_ctrl_op2_sel,
                io_deq_bits_uops_2_bits_ctrl_imm_sel,
  output [3:0]  io_deq_bits_uops_2_bits_ctrl_op_fcn,
  output        io_deq_bits_uops_2_bits_ctrl_fcn_dw,
  output [2:0]  io_deq_bits_uops_2_bits_ctrl_csr_cmd,
  output        io_deq_bits_uops_2_bits_ctrl_is_load,
                io_deq_bits_uops_2_bits_ctrl_is_sta,
                io_deq_bits_uops_2_bits_ctrl_is_std,
  output [1:0]  io_deq_bits_uops_2_bits_iw_state,
  output        io_deq_bits_uops_2_bits_iw_p1_poisoned,
                io_deq_bits_uops_2_bits_iw_p2_poisoned,
                io_deq_bits_uops_2_bits_is_sfb,
  output [4:0]  io_deq_bits_uops_2_bits_ftq_idx,
  output        io_deq_bits_uops_2_bits_edge_inst,
  output [5:0]  io_deq_bits_uops_2_bits_pc_lob,
  output        io_deq_bits_uops_2_bits_taken,
  output [11:0] io_deq_bits_uops_2_bits_csr_addr,
  output [1:0]  io_deq_bits_uops_2_bits_rxq_idx,
  output        io_deq_bits_uops_2_bits_xcpt_pf_if,
                io_deq_bits_uops_2_bits_xcpt_ae_if,
                io_deq_bits_uops_2_bits_xcpt_ma_if,
                io_deq_bits_uops_2_bits_bp_debug_if,
                io_deq_bits_uops_2_bits_bp_xcpt_if,
  output [1:0]  io_deq_bits_uops_2_bits_debug_fsrc,
                io_deq_bits_uops_2_bits_debug_tsrc
);

  reg  [31:0] fb_uop_ram_0_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_0_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_0_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_0_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_0_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_0_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_0_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_0_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_0_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_0_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_0_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_0_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_0_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_0_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_0_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_0_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_0_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_1_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_1_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_1_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_1_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_1_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_1_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_1_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_1_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_1_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_1_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_1_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_1_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_1_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_1_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_1_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_1_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_1_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_2_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_2_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_2_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_2_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_2_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_2_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_2_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_2_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_2_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_2_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_2_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_2_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_2_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_2_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_2_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_2_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_2_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_3_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_3_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_3_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_3_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_3_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_3_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_3_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_3_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_3_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_3_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_3_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_3_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_3_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_3_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_3_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_3_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_3_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_4_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_4_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_4_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_4_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_4_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_4_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_4_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_4_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_4_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_4_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_4_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_4_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_4_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_4_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_4_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_4_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_4_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_5_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_5_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_5_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_5_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_5_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_5_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_5_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_5_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_5_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_5_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_5_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_5_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_5_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_5_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_5_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_5_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_5_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_6_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_6_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_6_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_6_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_6_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_6_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_6_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_6_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_6_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_6_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_6_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_6_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_6_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_6_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_6_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_6_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_6_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_7_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_7_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_7_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_7_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_7_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_7_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_7_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_7_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_7_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_7_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_7_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_7_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_7_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_7_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_7_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_7_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_7_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_8_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_8_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_8_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_8_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_8_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_8_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_8_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_8_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_8_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_8_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_8_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_8_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_8_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_8_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_8_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_8_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_8_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_9_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_9_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_9_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_9_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_9_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_9_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_9_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_9_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_9_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_9_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_9_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_9_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_9_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_9_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_9_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_9_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_9_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_10_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_10_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_10_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_10_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_10_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_10_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_10_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_10_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_10_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_10_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_10_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_10_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_10_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_10_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_10_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_10_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_10_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_11_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_11_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_11_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_11_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_11_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_11_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_11_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_11_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_11_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_11_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_11_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_11_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_11_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_11_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_11_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_11_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_11_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_12_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_12_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_12_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_12_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_12_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_12_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_12_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_12_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_12_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_12_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_12_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_12_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_12_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_12_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_12_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_12_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_12_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_13_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_13_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_13_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_13_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_13_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_13_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_13_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_13_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_13_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_13_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_13_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_13_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_13_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_13_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_13_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_13_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_13_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_14_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_14_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_14_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_14_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_14_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_14_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_14_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_14_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_14_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_14_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_14_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_14_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_14_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_14_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_14_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_14_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_14_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_15_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_15_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_15_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_15_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_15_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_15_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_15_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_15_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_15_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_15_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_15_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_15_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_15_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_15_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_15_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_15_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_15_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_16_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_16_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_16_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_16_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_16_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_16_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_16_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_16_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_16_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_16_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_16_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_16_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_16_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_16_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_16_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_16_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_16_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_17_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_17_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_17_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_17_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_17_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_17_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_17_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_17_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_17_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_17_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_17_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_17_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_17_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_17_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_17_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_17_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_17_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_18_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_18_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_18_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_18_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_18_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_18_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_18_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_18_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_18_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_18_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_18_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_18_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_18_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_18_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_18_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_18_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_18_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_19_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_19_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_19_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_19_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_19_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_19_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_19_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_19_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_19_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_19_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_19_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_19_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_19_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_19_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_19_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_19_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_19_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_20_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_20_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_20_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_20_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_20_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_20_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_20_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_20_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_20_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_20_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_20_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_20_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_20_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_20_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_20_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_20_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_20_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_21_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_21_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_21_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_21_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_21_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_21_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_21_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_21_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_21_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_21_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_21_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_21_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_21_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_21_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_21_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_21_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_21_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_22_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_22_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_22_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_22_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_22_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_22_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_22_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_22_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_22_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_22_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_22_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_22_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_22_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_22_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_22_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_22_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_22_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_23_inst;	// fetch-buffer.scala:57:16
  reg  [31:0] fb_uop_ram_23_debug_inst;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_is_rvc;	// fetch-buffer.scala:57:16
  reg  [39:0] fb_uop_ram_23_debug_pc;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_23_ctrl_br_type;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_23_ctrl_op1_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_23_ctrl_op2_sel;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_23_ctrl_imm_sel;	// fetch-buffer.scala:57:16
  reg  [3:0]  fb_uop_ram_23_ctrl_op_fcn;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_ctrl_fcn_dw;	// fetch-buffer.scala:57:16
  reg  [2:0]  fb_uop_ram_23_ctrl_csr_cmd;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_ctrl_is_load;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_ctrl_is_sta;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_ctrl_is_std;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_23_iw_state;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_iw_p1_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_iw_p2_poisoned;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_is_sfb;	// fetch-buffer.scala:57:16
  reg  [4:0]  fb_uop_ram_23_ftq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_edge_inst;	// fetch-buffer.scala:57:16
  reg  [5:0]  fb_uop_ram_23_pc_lob;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_taken;	// fetch-buffer.scala:57:16
  reg  [11:0] fb_uop_ram_23_csr_addr;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_23_rxq_idx;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_xcpt_pf_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_xcpt_ae_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_xcpt_ma_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_bp_debug_if;	// fetch-buffer.scala:57:16
  reg         fb_uop_ram_23_bp_xcpt_if;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_23_debug_fsrc;	// fetch-buffer.scala:57:16
  reg  [1:0]  fb_uop_ram_23_debug_tsrc;	// fetch-buffer.scala:57:16
  reg  [7:0]  head;	// fetch-buffer.scala:61:21
  reg  [23:0] tail;	// fetch-buffer.scala:62:21
  reg         maybe_full;	// fetch-buffer.scala:64:27
  wire        _do_enq_T_1 =
    (|({tail[21], tail[18], tail[15], tail[12], tail[9], tail[6], tail[3], tail[0]}
       & head)) & maybe_full
    | (|(head
         & {tail[20], tail[17], tail[14], tail[11], tail[8], tail[5], tail[2], tail[23]}
         | head
         & {tail[19], tail[16], tail[13], tail[10], tail[7], tail[4], tail[1], tail[22]}
         | head
         & {tail[18], tail[15], tail[12], tail[9], tail[6], tail[3], tail[0], tail[21]}
         | head
         & {tail[17], tail[14], tail[11], tail[8], tail[5], tail[2], tail[23], tail[20]}
         | head
         & {tail[16], tail[13], tail[10], tail[7], tail[4], tail[1], tail[22], tail[19]}
         | head
         & {tail[15], tail[12], tail[9], tail[6], tail[3], tail[0], tail[21], tail[18]}
         | head
         & {tail[14],
            tail[11],
            tail[8],
            tail[5],
            tail[2],
            tail[23],
            tail[20],
            tail[17]}));	// fetch-buffer.scala:61:21, :62:21, :64:27, :75:24, :78:82, :79:{63,88,104,108}, :80:31, :81:{29,36,44}, :82:{26,40}
  wire [2:0]  slot_will_hit_tail =
    {{2{head[0]}}, head[0] & ~maybe_full} & tail[2:0]
    | {{2{head[1]}}, head[1] & ~maybe_full} & tail[5:3]
    | {{2{head[2]}}, head[2] & ~maybe_full} & tail[8:6]
    | {{2{head[3]}}, head[3] & ~maybe_full} & tail[11:9]
    | {{2{head[4]}}, head[4] & ~maybe_full} & tail[14:12]
    | {{2{head[5]}}, head[5] & ~maybe_full} & tail[17:15]
    | {{2{head[6]}}, head[6] & ~maybe_full} & tail[20:18]
    | {{2{head[7]}}, head[7] & ~maybe_full} & tail[23:21];	// fetch-buffer.scala:61:21, :62:21, :64:27, :155:{31,45,49,90,97}, :156:{70,112}
  wire [2:0]  _deq_valids_T_7 =
    slot_will_hit_tail
    | {slot_will_hit_tail[1] | slot_will_hit_tail[0], slot_will_hit_tail[0], 1'h0};	// fetch-buffer.scala:156:112, util.scala:384:{37,54}
  wire [2:0]  _deq_valids_T_8 = ~_deq_valids_T_7;	// fetch-buffer.scala:161:21, util.scala:384:54
  always @(posedge clock) begin
    automatic logic [39:0] pc;	// frontend.scala:161:39
    automatic logic        in_mask_0;	// fetch-buffer.scala:98:49
    automatic logic [39:0] _GEN = {io_enq_bits_pc[39:3], 3'h0};	// fetch-buffer.scala:97:33, :107:81
    automatic logic [39:0] _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:107:81
    automatic logic [5:0]  in_uops_0_pc_lob;	// fetch-buffer.scala:101:33, :106:41, :108:32
    automatic logic        in_uops_0_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_0_taken;	// fetch-buffer.scala:116:69
    automatic logic [39:0] _pc_T_7;	// fetch-buffer.scala:95:43
    automatic logic        in_mask_1;	// fetch-buffer.scala:98:49
    automatic logic        in_uops_1_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_1_taken;	// fetch-buffer.scala:116:69
    automatic logic [39:0] _pc_T_11;	// fetch-buffer.scala:95:43
    automatic logic        in_mask_2;	// fetch-buffer.scala:98:49
    automatic logic        in_uops_2_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_2_taken;	// fetch-buffer.scala:116:69
    automatic logic [39:0] _pc_T_15;	// fetch-buffer.scala:95:43
    automatic logic        in_mask_3;	// fetch-buffer.scala:98:49
    automatic logic        in_uops_3_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_3_taken;	// fetch-buffer.scala:116:69
    automatic logic [39:0] _pc_T_19;	// fetch-buffer.scala:95:43
    automatic logic        in_mask_4;	// fetch-buffer.scala:98:49
    automatic logic [39:0] _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:107:81
    automatic logic [5:0]  _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:108:61
    automatic logic        in_uops_4_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_4_taken;	// fetch-buffer.scala:116:69
    automatic logic [39:0] _pc_T_23;	// fetch-buffer.scala:95:43
    automatic logic        in_mask_5;	// fetch-buffer.scala:98:49
    automatic logic        in_uops_5_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_5_taken;	// fetch-buffer.scala:116:69
    automatic logic [39:0] _pc_T_27;	// fetch-buffer.scala:95:43
    automatic logic        in_mask_6;	// fetch-buffer.scala:98:49
    automatic logic        in_uops_6_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_6_taken;	// fetch-buffer.scala:116:69
    automatic logic [39:0] _pc_T_31;	// fetch-buffer.scala:95:43
    automatic logic        in_mask_7;	// fetch-buffer.scala:98:49
    automatic logic        in_uops_7_is_rvc;	// fetch-buffer.scala:115:62
    automatic logic        in_uops_7_taken;	// fetch-buffer.scala:116:69
    automatic logic [23:0] _GEN_0;	// Cat.scala:30:58
    automatic logic [23:0] enq_idxs_1;	// fetch-buffer.scala:138:18
    automatic logic [23:0] _GEN_1;	// Cat.scala:30:58
    automatic logic [23:0] enq_idxs_2;	// fetch-buffer.scala:138:18
    automatic logic [23:0] _GEN_2;	// Cat.scala:30:58
    automatic logic [23:0] enq_idxs_3;	// fetch-buffer.scala:138:18
    automatic logic [23:0] _GEN_3;	// Cat.scala:30:58
    automatic logic [23:0] enq_idxs_4;	// fetch-buffer.scala:138:18
    automatic logic [23:0] _GEN_4;	// Cat.scala:30:58
    automatic logic [23:0] enq_idxs_5;	// fetch-buffer.scala:138:18
    automatic logic [23:0] _GEN_5;	// Cat.scala:30:58
    automatic logic [23:0] enq_idxs_6;	// fetch-buffer.scala:138:18
    automatic logic [23:0] _GEN_6;	// Cat.scala:30:58
    automatic logic [23:0] enq_idxs_7;	// fetch-buffer.scala:138:18
    automatic logic        _GEN_7;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_8;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_9;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_10;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_11;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_12;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_13;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_14;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_15;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_16;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_17;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_18;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_19;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_20;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_21;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_22;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_23;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_24;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_25;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_26;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_27;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_28;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_29;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_30;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_31;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_32;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_33;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_34;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_35;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_36;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_37;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_38;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_39;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_40;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_41;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_42;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_43;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_44;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_45;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_46;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_47;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_48;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_49;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_50;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_51;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_52;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_53;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_54;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_55;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_56;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_57;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_58;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_59;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_60;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_61;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_62;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_63;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_64;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_65;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_66;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_67;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_68;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_69;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_70;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_71;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_72;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_73;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_74;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_75;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_76;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_77;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_78;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_79;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_80;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_81;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_82;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_83;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_84;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_85;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_86;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_87;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_88;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_89;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_90;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_91;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_92;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_93;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_94;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_95;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_96;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_97;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_98;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_99;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_100;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_101;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_102;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_103;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_104;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_105;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_106;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_107;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_108;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_109;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_110;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_111;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_112;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_113;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_114;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_115;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_116;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_117;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_118;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_119;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_120;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_121;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_122;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_123;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_124;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_125;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_126;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_127;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_128;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_129;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_130;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_131;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_132;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_133;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_134;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_135;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_136;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_137;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_138;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_139;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_140;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_141;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_142;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_143;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_144;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_145;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_146;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_147;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_148;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_149;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_150;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_151;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_152;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_153;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_154;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_155;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_156;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_157;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_158;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_159;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_160;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_161;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_162;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_163;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_164;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_165;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_166;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_167;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_168;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_169;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_170;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_171;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_172;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_173;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_174;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_175;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_176;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_177;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_178;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_179;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_180;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_181;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_182;	// fetch-buffer.scala:144:20
    automatic logic        _GEN_183;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_184;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_185;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_186;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_187;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_188;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_189;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_190;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_191;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_192;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_193;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_194;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_195;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_196;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_197;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_198;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_199;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_200;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_201;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_202;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_203;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_204;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_205;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_206;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_207;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_208;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_209;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_210;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_211;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_212;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_213;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_214;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_215;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_216;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_217;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_218;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_219;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_220;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_221;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_222;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_223;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_224;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_225;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_226;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_227;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_228;	// fetch-buffer.scala:57:16, :144:53, :145:16
    automatic logic        _GEN_229;	// fetch-buffer.scala:144:34
    automatic logic        _GEN_230;	// fetch-buffer.scala:57:16, :144:53, :145:16
    pc = {io_enq_bits_pc[39:3], 3'h0};	// fetch-buffer.scala:97:33, frontend.scala:161:39
    in_mask_0 = io_enq_valid & io_enq_bits_mask[0];	// fetch-buffer.scala:98:{49,68}
    _in_uops_0_debug_pc_T_5 = _GEN - 40'h2;	// fetch-buffer.scala:107:81
    in_uops_0_pc_lob = {io_enq_bits_pc[5:3], 3'h0};	// fetch-buffer.scala:97:33, :101:33, :106:41, :108:32
    in_uops_0_is_rvc = io_enq_bits_insts_0[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_0_taken = io_enq_bits_cfi_idx_bits == 3'h0 & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:97:33, :116:{61,69}
    _pc_T_7 = _GEN + 40'h2;	// fetch-buffer.scala:95:43, :107:81
    in_mask_1 = io_enq_valid & io_enq_bits_mask[1];	// fetch-buffer.scala:98:{49,68}
    in_uops_1_is_rvc = io_enq_bits_insts_1[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_1_taken = io_enq_bits_cfi_idx_bits == 3'h1 & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:116:{61,69}
    _pc_T_11 = _GEN + 40'h4;	// fetch-buffer.scala:95:43, :107:81
    in_mask_2 = io_enq_valid & io_enq_bits_mask[2];	// fetch-buffer.scala:98:{49,68}
    in_uops_2_is_rvc = io_enq_bits_insts_2[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_2_taken = io_enq_bits_cfi_idx_bits == 3'h2 & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:116:{61,69}
    _pc_T_15 = _GEN + 40'h6;	// fetch-buffer.scala:95:43, :107:81
    in_mask_3 = io_enq_valid & io_enq_bits_mask[3];	// fetch-buffer.scala:98:{49,68}
    in_uops_3_is_rvc = io_enq_bits_insts_3[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_3_taken = io_enq_bits_cfi_idx_bits == 3'h3 & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:116:{61,69}
    _pc_T_19 = _GEN + 40'h8;	// fetch-buffer.scala:95:43, :107:81
    in_mask_4 = io_enq_valid & io_enq_bits_mask[4];	// fetch-buffer.scala:98:{49,68}
    _in_uops_4_debug_pc_T_5 = _GEN + 40'h6;	// fetch-buffer.scala:95:43, :107:81
    _in_uops_4_pc_lob_T_3 = {io_enq_bits_pc[5:3], 3'h0} + 6'h8;	// fetch-buffer.scala:95:43, :97:33, :101:33, :108:61
    in_uops_4_is_rvc = io_enq_bits_insts_4[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_4_taken = io_enq_bits_cfi_idx_bits == 3'h4 & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:95:43, :116:{61,69}
    _pc_T_23 = _GEN + 40'hA;	// fetch-buffer.scala:95:43, :107:81
    in_mask_5 = io_enq_valid & io_enq_bits_mask[5];	// fetch-buffer.scala:98:{49,68}
    in_uops_5_is_rvc = io_enq_bits_insts_5[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_5_taken = io_enq_bits_cfi_idx_bits == 3'h5 & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:116:{61,69}
    _pc_T_27 = _GEN + 40'hC;	// fetch-buffer.scala:95:43, :107:81
    in_mask_6 = io_enq_valid & io_enq_bits_mask[6];	// fetch-buffer.scala:98:{49,68}
    in_uops_6_is_rvc = io_enq_bits_insts_6[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_6_taken = io_enq_bits_cfi_idx_bits == 3'h6 & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:95:43, :116:{61,69}
    _pc_T_31 = _GEN + 40'hE;	// fetch-buffer.scala:95:43, :107:81
    in_mask_7 = io_enq_valid & io_enq_bits_mask[7];	// fetch-buffer.scala:98:{49,68}
    in_uops_7_is_rvc = io_enq_bits_insts_7[1:0] != 2'h3;	// fetch-buffer.scala:115:{56,62}
    in_uops_7_taken = (&io_enq_bits_cfi_idx_bits) & io_enq_bits_cfi_idx_valid;	// fetch-buffer.scala:116:{61,69}
    _GEN_0 = {tail[22:0], tail[23]};	// Cat.scala:30:58, fetch-buffer.scala:62:21, :75:{11,24}
    enq_idxs_1 = in_mask_0 ? _GEN_0 : tail;	// Cat.scala:30:58, fetch-buffer.scala:62:21, :98:49, :138:18
    _GEN_1 = {enq_idxs_1[22:0], enq_idxs_1[23]};	// Cat.scala:30:58, fetch-buffer.scala:132:{12,24}, :138:18
    enq_idxs_2 = in_mask_1 ? _GEN_1 : enq_idxs_1;	// Cat.scala:30:58, fetch-buffer.scala:98:49, :138:18
    _GEN_2 = {enq_idxs_2[22:0], enq_idxs_2[23]};	// Cat.scala:30:58, fetch-buffer.scala:132:{12,24}, :138:18
    enq_idxs_3 = in_mask_2 ? _GEN_2 : enq_idxs_2;	// Cat.scala:30:58, fetch-buffer.scala:98:49, :138:18
    _GEN_3 = {enq_idxs_3[22:0], enq_idxs_3[23]};	// Cat.scala:30:58, fetch-buffer.scala:132:{12,24}, :138:18
    enq_idxs_4 = in_mask_3 ? _GEN_3 : enq_idxs_3;	// Cat.scala:30:58, fetch-buffer.scala:98:49, :138:18
    _GEN_4 = {enq_idxs_4[22:0], enq_idxs_4[23]};	// Cat.scala:30:58, fetch-buffer.scala:132:{12,24}, :138:18
    enq_idxs_5 = in_mask_4 ? _GEN_4 : enq_idxs_4;	// Cat.scala:30:58, fetch-buffer.scala:98:49, :138:18
    _GEN_5 = {enq_idxs_5[22:0], enq_idxs_5[23]};	// Cat.scala:30:58, fetch-buffer.scala:132:{12,24}, :138:18
    enq_idxs_6 = in_mask_5 ? _GEN_5 : enq_idxs_5;	// Cat.scala:30:58, fetch-buffer.scala:98:49, :138:18
    _GEN_6 = {enq_idxs_6[22:0], enq_idxs_6[23]};	// Cat.scala:30:58, fetch-buffer.scala:132:{12,24}, :138:18
    enq_idxs_7 = in_mask_6 ? _GEN_6 : enq_idxs_6;	// Cat.scala:30:58, fetch-buffer.scala:98:49, :138:18
    _GEN_7 = ~_do_enq_T_1 & in_mask_0;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_8 = _GEN_7 & tail[0];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_9 = _GEN_7 & tail[1];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_10 = _GEN_7 & tail[2];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_11 = _GEN_7 & tail[3];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_12 = _GEN_7 & tail[4];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_13 = _GEN_7 & tail[5];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_14 = _GEN_7 & tail[6];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_15 = _GEN_7 & tail[7];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_16 = _GEN_7 & tail[8];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_17 = _GEN_7 & tail[9];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_18 = _GEN_7 & tail[10];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_19 = _GEN_7 & tail[11];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_20 = _GEN_7 & tail[12];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_21 = _GEN_7 & tail[13];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_22 = _GEN_7 & tail[14];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_23 = _GEN_7 & tail[15];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_24 = _GEN_7 & tail[16];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_25 = _GEN_7 & tail[17];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_26 = _GEN_7 & tail[18];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_27 = _GEN_7 & tail[19];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_28 = _GEN_7 & tail[20];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_29 = _GEN_7 & tail[21];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_30 = _GEN_7 & tail[22];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_31 = _GEN_7 & tail[23];	// fetch-buffer.scala:62:21, :144:{20,34,48}
    _GEN_32 = ~_do_enq_T_1 & in_mask_1;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_33 = _GEN_32 & enq_idxs_1[0];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_34 = _GEN_32 & enq_idxs_1[1];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_35 = _GEN_32 & enq_idxs_1[2];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_36 = _GEN_32 & enq_idxs_1[3];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_37 = _GEN_32 & enq_idxs_1[4];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_38 = _GEN_32 & enq_idxs_1[5];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_39 = _GEN_32 & enq_idxs_1[6];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_40 = _GEN_32 & enq_idxs_1[7];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_41 = _GEN_32 & enq_idxs_1[8];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_42 = _GEN_32 & enq_idxs_1[9];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_43 = _GEN_32 & enq_idxs_1[10];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_44 = _GEN_32 & enq_idxs_1[11];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_45 = _GEN_32 & enq_idxs_1[12];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_46 = _GEN_32 & enq_idxs_1[13];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_47 = _GEN_32 & enq_idxs_1[14];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_48 = _GEN_32 & enq_idxs_1[15];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_49 = _GEN_32 & enq_idxs_1[16];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_50 = _GEN_32 & enq_idxs_1[17];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_51 = _GEN_32 & enq_idxs_1[18];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_52 = _GEN_32 & enq_idxs_1[19];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_53 = _GEN_32 & enq_idxs_1[20];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_54 = _GEN_32 & enq_idxs_1[21];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_55 = _GEN_32 & enq_idxs_1[22];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_56 = _GEN_32 & enq_idxs_1[23];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_57 = ~_do_enq_T_1 & in_mask_2;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_58 = _GEN_57 & enq_idxs_2[0];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_59 = _GEN_57 & enq_idxs_2[1];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_60 = _GEN_57 & enq_idxs_2[2];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_61 = _GEN_57 & enq_idxs_2[3];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_62 = _GEN_57 & enq_idxs_2[4];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_63 = _GEN_57 & enq_idxs_2[5];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_64 = _GEN_57 & enq_idxs_2[6];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_65 = _GEN_57 & enq_idxs_2[7];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_66 = _GEN_57 & enq_idxs_2[8];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_67 = _GEN_57 & enq_idxs_2[9];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_68 = _GEN_57 & enq_idxs_2[10];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_69 = _GEN_57 & enq_idxs_2[11];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_70 = _GEN_57 & enq_idxs_2[12];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_71 = _GEN_57 & enq_idxs_2[13];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_72 = _GEN_57 & enq_idxs_2[14];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_73 = _GEN_57 & enq_idxs_2[15];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_74 = _GEN_57 & enq_idxs_2[16];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_75 = _GEN_57 & enq_idxs_2[17];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_76 = _GEN_57 & enq_idxs_2[18];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_77 = _GEN_57 & enq_idxs_2[19];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_78 = _GEN_57 & enq_idxs_2[20];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_79 = _GEN_57 & enq_idxs_2[21];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_80 = _GEN_57 & enq_idxs_2[22];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_81 = _GEN_57 & enq_idxs_2[23];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_82 = ~_do_enq_T_1 & in_mask_3;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_83 = _GEN_82 & enq_idxs_3[0];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_84 = _GEN_82 & enq_idxs_3[1];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_85 = _GEN_82 & enq_idxs_3[2];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_86 = _GEN_82 & enq_idxs_3[3];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_87 = _GEN_82 & enq_idxs_3[4];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_88 = _GEN_82 & enq_idxs_3[5];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_89 = _GEN_82 & enq_idxs_3[6];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_90 = _GEN_82 & enq_idxs_3[7];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_91 = _GEN_82 & enq_idxs_3[8];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_92 = _GEN_82 & enq_idxs_3[9];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_93 = _GEN_82 & enq_idxs_3[10];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_94 = _GEN_82 & enq_idxs_3[11];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_95 = _GEN_82 & enq_idxs_3[12];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_96 = _GEN_82 & enq_idxs_3[13];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_97 = _GEN_82 & enq_idxs_3[14];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_98 = _GEN_82 & enq_idxs_3[15];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_99 = _GEN_82 & enq_idxs_3[16];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_100 = _GEN_82 & enq_idxs_3[17];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_101 = _GEN_82 & enq_idxs_3[18];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_102 = _GEN_82 & enq_idxs_3[19];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_103 = _GEN_82 & enq_idxs_3[20];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_104 = _GEN_82 & enq_idxs_3[21];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_105 = _GEN_82 & enq_idxs_3[22];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_106 = _GEN_82 & enq_idxs_3[23];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_107 = ~_do_enq_T_1 & in_mask_4;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_108 = _GEN_107 & enq_idxs_4[0];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_109 = _GEN_107 & enq_idxs_4[1];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_110 = _GEN_107 & enq_idxs_4[2];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_111 = _GEN_107 & enq_idxs_4[3];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_112 = _GEN_107 & enq_idxs_4[4];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_113 = _GEN_107 & enq_idxs_4[5];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_114 = _GEN_107 & enq_idxs_4[6];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_115 = _GEN_107 & enq_idxs_4[7];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_116 = _GEN_107 & enq_idxs_4[8];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_117 = _GEN_107 & enq_idxs_4[9];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_118 = _GEN_107 & enq_idxs_4[10];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_119 = _GEN_107 & enq_idxs_4[11];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_120 = _GEN_107 & enq_idxs_4[12];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_121 = _GEN_107 & enq_idxs_4[13];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_122 = _GEN_107 & enq_idxs_4[14];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_123 = _GEN_107 & enq_idxs_4[15];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_124 = _GEN_107 & enq_idxs_4[16];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_125 = _GEN_107 & enq_idxs_4[17];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_126 = _GEN_107 & enq_idxs_4[18];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_127 = _GEN_107 & enq_idxs_4[19];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_128 = _GEN_107 & enq_idxs_4[20];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_129 = _GEN_107 & enq_idxs_4[21];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_130 = _GEN_107 & enq_idxs_4[22];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_131 = _GEN_107 & enq_idxs_4[23];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_132 = ~_do_enq_T_1 & in_mask_5;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_133 = _GEN_132 & enq_idxs_5[0];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_134 = _GEN_132 & enq_idxs_5[1];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_135 = _GEN_132 & enq_idxs_5[2];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_136 = _GEN_132 & enq_idxs_5[3];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_137 = _GEN_132 & enq_idxs_5[4];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_138 = _GEN_132 & enq_idxs_5[5];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_139 = _GEN_132 & enq_idxs_5[6];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_140 = _GEN_132 & enq_idxs_5[7];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_141 = _GEN_132 & enq_idxs_5[8];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_142 = _GEN_132 & enq_idxs_5[9];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_143 = _GEN_132 & enq_idxs_5[10];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_144 = _GEN_132 & enq_idxs_5[11];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_145 = _GEN_132 & enq_idxs_5[12];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_146 = _GEN_132 & enq_idxs_5[13];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_147 = _GEN_132 & enq_idxs_5[14];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_148 = _GEN_132 & enq_idxs_5[15];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_149 = _GEN_132 & enq_idxs_5[16];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_150 = _GEN_132 & enq_idxs_5[17];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_151 = _GEN_132 & enq_idxs_5[18];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_152 = _GEN_132 & enq_idxs_5[19];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_153 = _GEN_132 & enq_idxs_5[20];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_154 = _GEN_132 & enq_idxs_5[21];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_155 = _GEN_132 & enq_idxs_5[22];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_156 = _GEN_132 & enq_idxs_5[23];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_157 = ~_do_enq_T_1 & in_mask_6;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_158 = _GEN_157 & enq_idxs_6[0];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_159 = _GEN_157 & enq_idxs_6[1];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_160 = _GEN_157 & enq_idxs_6[2];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_161 = _GEN_157 & enq_idxs_6[3];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_162 = _GEN_157 & enq_idxs_6[4];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_163 = _GEN_157 & enq_idxs_6[5];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_164 = _GEN_157 & enq_idxs_6[6];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_165 = _GEN_157 & enq_idxs_6[7];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_166 = _GEN_157 & enq_idxs_6[8];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_167 = _GEN_157 & enq_idxs_6[9];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_168 = _GEN_157 & enq_idxs_6[10];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_169 = _GEN_157 & enq_idxs_6[11];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_170 = _GEN_157 & enq_idxs_6[12];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_171 = _GEN_157 & enq_idxs_6[13];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_172 = _GEN_157 & enq_idxs_6[14];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_173 = _GEN_157 & enq_idxs_6[15];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_174 = _GEN_157 & enq_idxs_6[16];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_175 = _GEN_157 & enq_idxs_6[17];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_176 = _GEN_157 & enq_idxs_6[18];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_177 = _GEN_157 & enq_idxs_6[19];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_178 = _GEN_157 & enq_idxs_6[20];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_179 = _GEN_157 & enq_idxs_6[21];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_180 = _GEN_157 & enq_idxs_6[22];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_181 = _GEN_157 & enq_idxs_6[23];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_182 = ~_do_enq_T_1 & in_mask_7;	// fetch-buffer.scala:82:{16,40}, :98:49, :144:20
    _GEN_183 = _GEN_182 & enq_idxs_7[0];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_184 =
      _GEN_183 | _GEN_158 | _GEN_133 | _GEN_108 | _GEN_83 | _GEN_58 | _GEN_33 | _GEN_8;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_185 = _GEN_182 & enq_idxs_7[1];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_186 =
      _GEN_185 | _GEN_159 | _GEN_134 | _GEN_109 | _GEN_84 | _GEN_59 | _GEN_34 | _GEN_9;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_187 = _GEN_182 & enq_idxs_7[2];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_188 =
      _GEN_187 | _GEN_160 | _GEN_135 | _GEN_110 | _GEN_85 | _GEN_60 | _GEN_35 | _GEN_10;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_189 = _GEN_182 & enq_idxs_7[3];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_190 =
      _GEN_189 | _GEN_161 | _GEN_136 | _GEN_111 | _GEN_86 | _GEN_61 | _GEN_36 | _GEN_11;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_191 = _GEN_182 & enq_idxs_7[4];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_192 =
      _GEN_191 | _GEN_162 | _GEN_137 | _GEN_112 | _GEN_87 | _GEN_62 | _GEN_37 | _GEN_12;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_193 = _GEN_182 & enq_idxs_7[5];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_194 =
      _GEN_193 | _GEN_163 | _GEN_138 | _GEN_113 | _GEN_88 | _GEN_63 | _GEN_38 | _GEN_13;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_195 = _GEN_182 & enq_idxs_7[6];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_196 =
      _GEN_195 | _GEN_164 | _GEN_139 | _GEN_114 | _GEN_89 | _GEN_64 | _GEN_39 | _GEN_14;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_197 = _GEN_182 & enq_idxs_7[7];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_198 =
      _GEN_197 | _GEN_165 | _GEN_140 | _GEN_115 | _GEN_90 | _GEN_65 | _GEN_40 | _GEN_15;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_199 = _GEN_182 & enq_idxs_7[8];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_200 =
      _GEN_199 | _GEN_166 | _GEN_141 | _GEN_116 | _GEN_91 | _GEN_66 | _GEN_41 | _GEN_16;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_201 = _GEN_182 & enq_idxs_7[9];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_202 =
      _GEN_201 | _GEN_167 | _GEN_142 | _GEN_117 | _GEN_92 | _GEN_67 | _GEN_42 | _GEN_17;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_203 = _GEN_182 & enq_idxs_7[10];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_204 =
      _GEN_203 | _GEN_168 | _GEN_143 | _GEN_118 | _GEN_93 | _GEN_68 | _GEN_43 | _GEN_18;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_205 = _GEN_182 & enq_idxs_7[11];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_206 =
      _GEN_205 | _GEN_169 | _GEN_144 | _GEN_119 | _GEN_94 | _GEN_69 | _GEN_44 | _GEN_19;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_207 = _GEN_182 & enq_idxs_7[12];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_208 =
      _GEN_207 | _GEN_170 | _GEN_145 | _GEN_120 | _GEN_95 | _GEN_70 | _GEN_45 | _GEN_20;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_209 = _GEN_182 & enq_idxs_7[13];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_210 =
      _GEN_209 | _GEN_171 | _GEN_146 | _GEN_121 | _GEN_96 | _GEN_71 | _GEN_46 | _GEN_21;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_211 = _GEN_182 & enq_idxs_7[14];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_212 =
      _GEN_211 | _GEN_172 | _GEN_147 | _GEN_122 | _GEN_97 | _GEN_72 | _GEN_47 | _GEN_22;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_213 = _GEN_182 & enq_idxs_7[15];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_214 =
      _GEN_213 | _GEN_173 | _GEN_148 | _GEN_123 | _GEN_98 | _GEN_73 | _GEN_48 | _GEN_23;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_215 = _GEN_182 & enq_idxs_7[16];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_216 =
      _GEN_215 | _GEN_174 | _GEN_149 | _GEN_124 | _GEN_99 | _GEN_74 | _GEN_49 | _GEN_24;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_217 = _GEN_182 & enq_idxs_7[17];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_218 =
      _GEN_217 | _GEN_175 | _GEN_150 | _GEN_125 | _GEN_100 | _GEN_75 | _GEN_50 | _GEN_25;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_219 = _GEN_182 & enq_idxs_7[18];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_220 =
      _GEN_219 | _GEN_176 | _GEN_151 | _GEN_126 | _GEN_101 | _GEN_76 | _GEN_51 | _GEN_26;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_221 = _GEN_182 & enq_idxs_7[19];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_222 =
      _GEN_221 | _GEN_177 | _GEN_152 | _GEN_127 | _GEN_102 | _GEN_77 | _GEN_52 | _GEN_27;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_223 = _GEN_182 & enq_idxs_7[20];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_224 =
      _GEN_223 | _GEN_178 | _GEN_153 | _GEN_128 | _GEN_103 | _GEN_78 | _GEN_53 | _GEN_28;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_225 = _GEN_182 & enq_idxs_7[21];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_226 =
      _GEN_225 | _GEN_179 | _GEN_154 | _GEN_129 | _GEN_104 | _GEN_79 | _GEN_54 | _GEN_29;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_227 = _GEN_182 & enq_idxs_7[22];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_228 =
      _GEN_227 | _GEN_180 | _GEN_155 | _GEN_130 | _GEN_105 | _GEN_80 | _GEN_55 | _GEN_30;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    _GEN_229 = _GEN_182 & enq_idxs_7[23];	// fetch-buffer.scala:138:18, :144:{20,34,48}
    _GEN_230 =
      _GEN_229 | _GEN_181 | _GEN_156 | _GEN_131 | _GEN_106 | _GEN_81 | _GEN_56 | _GEN_31;	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    if (_GEN_183) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_0_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_0_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_158) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_0_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_0_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_133) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_0_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_0_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_108) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_0_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_0_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_0_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_0_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_83) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_0_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_0_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_58) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_0_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_0_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_33) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_0_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_0_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_8) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_0_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_0_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_0_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_0_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_0_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_0_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_184) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_0_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_0_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_0_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_0_ctrl_fcn_dw <= ~_GEN_184 & fb_uop_ram_0_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_0_ctrl_is_load <= ~_GEN_184 & fb_uop_ram_0_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_0_ctrl_is_sta <= ~_GEN_184 & fb_uop_ram_0_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_0_ctrl_is_std <= ~_GEN_184 & fb_uop_ram_0_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_0_iw_p1_poisoned <= ~_GEN_184 & fb_uop_ram_0_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_0_iw_p2_poisoned <= ~_GEN_184 & fb_uop_ram_0_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_0_edge_inst <=
      ~(_GEN_183 | _GEN_158 | _GEN_133)
      & (_GEN_108
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_83 | _GEN_58 | _GEN_33)
             & (_GEN_8 ? io_enq_bits_edge_inst_0 : fb_uop_ram_0_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_0_xcpt_ma_if <= ~_GEN_184 & fb_uop_ram_0_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_185) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_1_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_1_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_159) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_1_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_1_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_134) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_1_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_1_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_109) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_1_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_1_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_1_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_1_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_84) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_1_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_1_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_59) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_1_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_1_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_34) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_1_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_1_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_9) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_1_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_1_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_1_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_1_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_1_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_1_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_186) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_1_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_1_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_1_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_1_ctrl_fcn_dw <= ~_GEN_186 & fb_uop_ram_1_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_1_ctrl_is_load <= ~_GEN_186 & fb_uop_ram_1_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_1_ctrl_is_sta <= ~_GEN_186 & fb_uop_ram_1_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_1_ctrl_is_std <= ~_GEN_186 & fb_uop_ram_1_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_1_iw_p1_poisoned <= ~_GEN_186 & fb_uop_ram_1_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_1_iw_p2_poisoned <= ~_GEN_186 & fb_uop_ram_1_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_1_edge_inst <=
      ~(_GEN_185 | _GEN_159 | _GEN_134)
      & (_GEN_109
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_84 | _GEN_59 | _GEN_34)
             & (_GEN_9 ? io_enq_bits_edge_inst_0 : fb_uop_ram_1_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_1_xcpt_ma_if <= ~_GEN_186 & fb_uop_ram_1_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_187) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_2_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_2_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_160) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_2_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_2_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_135) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_2_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_2_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_110) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_2_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_2_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_2_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_2_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_85) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_2_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_2_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_60) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_2_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_2_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_35) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_2_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_2_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_10) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_2_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_2_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_2_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_2_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_2_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_2_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_188) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_2_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_2_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_2_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_2_ctrl_fcn_dw <= ~_GEN_188 & fb_uop_ram_2_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_2_ctrl_is_load <= ~_GEN_188 & fb_uop_ram_2_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_2_ctrl_is_sta <= ~_GEN_188 & fb_uop_ram_2_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_2_ctrl_is_std <= ~_GEN_188 & fb_uop_ram_2_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_2_iw_p1_poisoned <= ~_GEN_188 & fb_uop_ram_2_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_2_iw_p2_poisoned <= ~_GEN_188 & fb_uop_ram_2_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_2_edge_inst <=
      ~(_GEN_187 | _GEN_160 | _GEN_135)
      & (_GEN_110
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_85 | _GEN_60 | _GEN_35)
             & (_GEN_10 ? io_enq_bits_edge_inst_0 : fb_uop_ram_2_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_2_xcpt_ma_if <= ~_GEN_188 & fb_uop_ram_2_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_189) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_3_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_3_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_161) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_3_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_3_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_136) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_3_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_3_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_111) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_3_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_3_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_3_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_3_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_86) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_3_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_3_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_61) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_3_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_3_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_36) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_3_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_3_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_11) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_3_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_3_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_3_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_3_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_3_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_3_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_190) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_3_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_3_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_3_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_3_ctrl_fcn_dw <= ~_GEN_190 & fb_uop_ram_3_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_3_ctrl_is_load <= ~_GEN_190 & fb_uop_ram_3_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_3_ctrl_is_sta <= ~_GEN_190 & fb_uop_ram_3_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_3_ctrl_is_std <= ~_GEN_190 & fb_uop_ram_3_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_3_iw_p1_poisoned <= ~_GEN_190 & fb_uop_ram_3_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_3_iw_p2_poisoned <= ~_GEN_190 & fb_uop_ram_3_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_3_edge_inst <=
      ~(_GEN_189 | _GEN_161 | _GEN_136)
      & (_GEN_111
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_86 | _GEN_61 | _GEN_36)
             & (_GEN_11 ? io_enq_bits_edge_inst_0 : fb_uop_ram_3_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_3_xcpt_ma_if <= ~_GEN_190 & fb_uop_ram_3_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_191) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_4_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_4_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_162) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_4_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_4_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_137) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_4_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_4_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_112) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_4_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_4_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_4_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_4_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_87) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_4_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_4_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_62) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_4_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_4_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_37) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_4_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_4_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_12) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_4_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_4_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_4_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_4_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_4_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_4_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_192) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_4_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_4_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_4_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_4_ctrl_fcn_dw <= ~_GEN_192 & fb_uop_ram_4_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_4_ctrl_is_load <= ~_GEN_192 & fb_uop_ram_4_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_4_ctrl_is_sta <= ~_GEN_192 & fb_uop_ram_4_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_4_ctrl_is_std <= ~_GEN_192 & fb_uop_ram_4_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_4_iw_p1_poisoned <= ~_GEN_192 & fb_uop_ram_4_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_4_iw_p2_poisoned <= ~_GEN_192 & fb_uop_ram_4_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_4_edge_inst <=
      ~(_GEN_191 | _GEN_162 | _GEN_137)
      & (_GEN_112
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_87 | _GEN_62 | _GEN_37)
             & (_GEN_12 ? io_enq_bits_edge_inst_0 : fb_uop_ram_4_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_4_xcpt_ma_if <= ~_GEN_192 & fb_uop_ram_4_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_193) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_5_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_5_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_163) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_5_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_5_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_138) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_5_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_5_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_113) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_5_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_5_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_5_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_5_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_88) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_5_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_5_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_63) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_5_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_5_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_38) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_5_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_5_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_13) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_5_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_5_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_5_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_5_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_5_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_5_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_194) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_5_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_5_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_5_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_5_ctrl_fcn_dw <= ~_GEN_194 & fb_uop_ram_5_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_5_ctrl_is_load <= ~_GEN_194 & fb_uop_ram_5_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_5_ctrl_is_sta <= ~_GEN_194 & fb_uop_ram_5_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_5_ctrl_is_std <= ~_GEN_194 & fb_uop_ram_5_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_5_iw_p1_poisoned <= ~_GEN_194 & fb_uop_ram_5_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_5_iw_p2_poisoned <= ~_GEN_194 & fb_uop_ram_5_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_5_edge_inst <=
      ~(_GEN_193 | _GEN_163 | _GEN_138)
      & (_GEN_113
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_88 | _GEN_63 | _GEN_38)
             & (_GEN_13 ? io_enq_bits_edge_inst_0 : fb_uop_ram_5_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_5_xcpt_ma_if <= ~_GEN_194 & fb_uop_ram_5_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_195) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_6_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_6_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_164) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_6_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_6_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_139) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_6_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_6_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_114) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_6_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_6_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_6_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_6_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_89) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_6_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_6_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_64) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_6_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_6_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_39) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_6_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_6_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_14) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_6_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_6_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_6_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_6_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_6_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_6_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_196) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_6_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_6_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_6_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_6_ctrl_fcn_dw <= ~_GEN_196 & fb_uop_ram_6_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_6_ctrl_is_load <= ~_GEN_196 & fb_uop_ram_6_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_6_ctrl_is_sta <= ~_GEN_196 & fb_uop_ram_6_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_6_ctrl_is_std <= ~_GEN_196 & fb_uop_ram_6_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_6_iw_p1_poisoned <= ~_GEN_196 & fb_uop_ram_6_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_6_iw_p2_poisoned <= ~_GEN_196 & fb_uop_ram_6_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_6_edge_inst <=
      ~(_GEN_195 | _GEN_164 | _GEN_139)
      & (_GEN_114
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_89 | _GEN_64 | _GEN_39)
             & (_GEN_14 ? io_enq_bits_edge_inst_0 : fb_uop_ram_6_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_6_xcpt_ma_if <= ~_GEN_196 & fb_uop_ram_6_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_197) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_7_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_7_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_165) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_7_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_7_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_140) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_7_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_7_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_115) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_7_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_7_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_7_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_7_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_90) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_7_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_7_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_65) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_7_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_7_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_40) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_7_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_7_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_15) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_7_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_7_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_7_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_7_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_7_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_7_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_198) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_7_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_7_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_7_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_7_ctrl_fcn_dw <= ~_GEN_198 & fb_uop_ram_7_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_7_ctrl_is_load <= ~_GEN_198 & fb_uop_ram_7_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_7_ctrl_is_sta <= ~_GEN_198 & fb_uop_ram_7_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_7_ctrl_is_std <= ~_GEN_198 & fb_uop_ram_7_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_7_iw_p1_poisoned <= ~_GEN_198 & fb_uop_ram_7_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_7_iw_p2_poisoned <= ~_GEN_198 & fb_uop_ram_7_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_7_edge_inst <=
      ~(_GEN_197 | _GEN_165 | _GEN_140)
      & (_GEN_115
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_90 | _GEN_65 | _GEN_40)
             & (_GEN_15 ? io_enq_bits_edge_inst_0 : fb_uop_ram_7_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_7_xcpt_ma_if <= ~_GEN_198 & fb_uop_ram_7_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_199) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_8_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_8_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_166) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_8_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_8_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_141) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_8_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_8_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_116) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_8_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_8_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_8_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_8_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_91) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_8_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_8_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_66) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_8_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_8_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_41) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_8_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_8_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_16) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_8_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_8_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_8_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_8_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_8_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_8_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_200) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_8_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_8_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_8_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_8_ctrl_fcn_dw <= ~_GEN_200 & fb_uop_ram_8_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_8_ctrl_is_load <= ~_GEN_200 & fb_uop_ram_8_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_8_ctrl_is_sta <= ~_GEN_200 & fb_uop_ram_8_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_8_ctrl_is_std <= ~_GEN_200 & fb_uop_ram_8_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_8_iw_p1_poisoned <= ~_GEN_200 & fb_uop_ram_8_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_8_iw_p2_poisoned <= ~_GEN_200 & fb_uop_ram_8_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_8_edge_inst <=
      ~(_GEN_199 | _GEN_166 | _GEN_141)
      & (_GEN_116
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_91 | _GEN_66 | _GEN_41)
             & (_GEN_16 ? io_enq_bits_edge_inst_0 : fb_uop_ram_8_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_8_xcpt_ma_if <= ~_GEN_200 & fb_uop_ram_8_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_201) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_9_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_9_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_167) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_9_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_9_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_142) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_9_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_9_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_117) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_9_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_9_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_9_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_9_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_92) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_9_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_9_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_67) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_9_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_9_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_42) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_9_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_9_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_17) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_9_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_9_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_9_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_9_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_9_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_9_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_202) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_9_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_9_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_9_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_9_ctrl_fcn_dw <= ~_GEN_202 & fb_uop_ram_9_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_9_ctrl_is_load <= ~_GEN_202 & fb_uop_ram_9_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_9_ctrl_is_sta <= ~_GEN_202 & fb_uop_ram_9_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_9_ctrl_is_std <= ~_GEN_202 & fb_uop_ram_9_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_9_iw_p1_poisoned <= ~_GEN_202 & fb_uop_ram_9_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_9_iw_p2_poisoned <= ~_GEN_202 & fb_uop_ram_9_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_9_edge_inst <=
      ~(_GEN_201 | _GEN_167 | _GEN_142)
      & (_GEN_117
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_92 | _GEN_67 | _GEN_42)
             & (_GEN_17 ? io_enq_bits_edge_inst_0 : fb_uop_ram_9_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_9_xcpt_ma_if <= ~_GEN_202 & fb_uop_ram_9_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_203) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_10_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_10_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_168) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_10_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_10_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_143) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_10_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_10_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_118) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_10_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_10_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_10_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_10_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_93) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_10_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_10_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_68) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_10_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_10_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_43) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_10_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_10_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_18) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_10_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_10_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_10_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_10_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_10_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_10_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_204) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_10_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_10_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_10_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_10_ctrl_fcn_dw <= ~_GEN_204 & fb_uop_ram_10_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_10_ctrl_is_load <= ~_GEN_204 & fb_uop_ram_10_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_10_ctrl_is_sta <= ~_GEN_204 & fb_uop_ram_10_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_10_ctrl_is_std <= ~_GEN_204 & fb_uop_ram_10_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_10_iw_p1_poisoned <= ~_GEN_204 & fb_uop_ram_10_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_10_iw_p2_poisoned <= ~_GEN_204 & fb_uop_ram_10_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_10_edge_inst <=
      ~(_GEN_203 | _GEN_168 | _GEN_143)
      & (_GEN_118
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_93 | _GEN_68 | _GEN_43)
             & (_GEN_18 ? io_enq_bits_edge_inst_0 : fb_uop_ram_10_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_10_xcpt_ma_if <= ~_GEN_204 & fb_uop_ram_10_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_205) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_11_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_11_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_169) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_11_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_11_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_144) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_11_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_11_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_119) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_11_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_11_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_11_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_11_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_94) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_11_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_11_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_69) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_11_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_11_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_44) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_11_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_11_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_19) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_11_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_11_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_11_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_11_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_11_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_11_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_206) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_11_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_11_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_11_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_11_ctrl_fcn_dw <= ~_GEN_206 & fb_uop_ram_11_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_11_ctrl_is_load <= ~_GEN_206 & fb_uop_ram_11_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_11_ctrl_is_sta <= ~_GEN_206 & fb_uop_ram_11_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_11_ctrl_is_std <= ~_GEN_206 & fb_uop_ram_11_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_11_iw_p1_poisoned <= ~_GEN_206 & fb_uop_ram_11_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_11_iw_p2_poisoned <= ~_GEN_206 & fb_uop_ram_11_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_11_edge_inst <=
      ~(_GEN_205 | _GEN_169 | _GEN_144)
      & (_GEN_119
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_94 | _GEN_69 | _GEN_44)
             & (_GEN_19 ? io_enq_bits_edge_inst_0 : fb_uop_ram_11_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_11_xcpt_ma_if <= ~_GEN_206 & fb_uop_ram_11_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_207) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_12_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_12_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_170) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_12_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_12_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_145) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_12_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_12_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_120) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_12_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_12_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_12_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_12_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_95) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_12_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_12_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_70) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_12_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_12_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_45) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_12_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_12_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_20) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_12_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_12_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_12_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_12_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_12_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_12_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_208) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_12_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_12_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_12_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_12_ctrl_fcn_dw <= ~_GEN_208 & fb_uop_ram_12_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_12_ctrl_is_load <= ~_GEN_208 & fb_uop_ram_12_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_12_ctrl_is_sta <= ~_GEN_208 & fb_uop_ram_12_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_12_ctrl_is_std <= ~_GEN_208 & fb_uop_ram_12_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_12_iw_p1_poisoned <= ~_GEN_208 & fb_uop_ram_12_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_12_iw_p2_poisoned <= ~_GEN_208 & fb_uop_ram_12_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_12_edge_inst <=
      ~(_GEN_207 | _GEN_170 | _GEN_145)
      & (_GEN_120
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_95 | _GEN_70 | _GEN_45)
             & (_GEN_20 ? io_enq_bits_edge_inst_0 : fb_uop_ram_12_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_12_xcpt_ma_if <= ~_GEN_208 & fb_uop_ram_12_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_209) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_13_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_13_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_171) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_13_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_13_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_146) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_13_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_13_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_121) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_13_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_13_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_13_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_13_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_96) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_13_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_13_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_71) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_13_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_13_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_46) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_13_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_13_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_21) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_13_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_13_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_13_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_13_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_13_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_13_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_210) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_13_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_13_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_13_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_13_ctrl_fcn_dw <= ~_GEN_210 & fb_uop_ram_13_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_13_ctrl_is_load <= ~_GEN_210 & fb_uop_ram_13_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_13_ctrl_is_sta <= ~_GEN_210 & fb_uop_ram_13_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_13_ctrl_is_std <= ~_GEN_210 & fb_uop_ram_13_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_13_iw_p1_poisoned <= ~_GEN_210 & fb_uop_ram_13_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_13_iw_p2_poisoned <= ~_GEN_210 & fb_uop_ram_13_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_13_edge_inst <=
      ~(_GEN_209 | _GEN_171 | _GEN_146)
      & (_GEN_121
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_96 | _GEN_71 | _GEN_46)
             & (_GEN_21 ? io_enq_bits_edge_inst_0 : fb_uop_ram_13_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_13_xcpt_ma_if <= ~_GEN_210 & fb_uop_ram_13_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_211) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_14_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_14_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_172) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_14_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_14_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_147) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_14_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_14_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_122) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_14_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_14_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_14_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_14_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_97) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_14_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_14_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_72) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_14_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_14_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_47) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_14_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_14_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_22) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_14_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_14_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_14_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_14_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_14_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_14_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_212) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_14_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_14_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_14_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_14_ctrl_fcn_dw <= ~_GEN_212 & fb_uop_ram_14_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_14_ctrl_is_load <= ~_GEN_212 & fb_uop_ram_14_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_14_ctrl_is_sta <= ~_GEN_212 & fb_uop_ram_14_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_14_ctrl_is_std <= ~_GEN_212 & fb_uop_ram_14_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_14_iw_p1_poisoned <= ~_GEN_212 & fb_uop_ram_14_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_14_iw_p2_poisoned <= ~_GEN_212 & fb_uop_ram_14_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_14_edge_inst <=
      ~(_GEN_211 | _GEN_172 | _GEN_147)
      & (_GEN_122
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_97 | _GEN_72 | _GEN_47)
             & (_GEN_22 ? io_enq_bits_edge_inst_0 : fb_uop_ram_14_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_14_xcpt_ma_if <= ~_GEN_212 & fb_uop_ram_14_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_213) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_15_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_15_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_173) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_15_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_15_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_148) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_15_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_15_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_123) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_15_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_15_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_15_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_15_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_98) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_15_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_15_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_73) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_15_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_15_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_48) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_15_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_15_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_23) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_15_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_15_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_15_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_15_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_15_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_15_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_214) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_15_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_15_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_15_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_15_ctrl_fcn_dw <= ~_GEN_214 & fb_uop_ram_15_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_15_ctrl_is_load <= ~_GEN_214 & fb_uop_ram_15_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_15_ctrl_is_sta <= ~_GEN_214 & fb_uop_ram_15_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_15_ctrl_is_std <= ~_GEN_214 & fb_uop_ram_15_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_15_iw_p1_poisoned <= ~_GEN_214 & fb_uop_ram_15_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_15_iw_p2_poisoned <= ~_GEN_214 & fb_uop_ram_15_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_15_edge_inst <=
      ~(_GEN_213 | _GEN_173 | _GEN_148)
      & (_GEN_123
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_98 | _GEN_73 | _GEN_48)
             & (_GEN_23 ? io_enq_bits_edge_inst_0 : fb_uop_ram_15_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_15_xcpt_ma_if <= ~_GEN_214 & fb_uop_ram_15_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_215) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_16_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_16_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_174) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_16_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_16_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_149) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_16_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_16_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_124) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_16_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_16_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_16_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_16_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_99) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_16_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_16_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_74) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_16_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_16_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_49) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_16_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_16_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_24) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_16_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_16_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_16_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_16_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_16_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_16_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_216) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_16_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_16_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_16_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_16_ctrl_fcn_dw <= ~_GEN_216 & fb_uop_ram_16_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_16_ctrl_is_load <= ~_GEN_216 & fb_uop_ram_16_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_16_ctrl_is_sta <= ~_GEN_216 & fb_uop_ram_16_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_16_ctrl_is_std <= ~_GEN_216 & fb_uop_ram_16_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_16_iw_p1_poisoned <= ~_GEN_216 & fb_uop_ram_16_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_16_iw_p2_poisoned <= ~_GEN_216 & fb_uop_ram_16_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_16_edge_inst <=
      ~(_GEN_215 | _GEN_174 | _GEN_149)
      & (_GEN_124
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_99 | _GEN_74 | _GEN_49)
             & (_GEN_24 ? io_enq_bits_edge_inst_0 : fb_uop_ram_16_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_16_xcpt_ma_if <= ~_GEN_216 & fb_uop_ram_16_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_217) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_17_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_17_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_175) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_17_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_17_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_150) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_17_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_17_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_125) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_17_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_17_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_17_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_17_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_100) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_17_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_17_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_75) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_17_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_17_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_50) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_17_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_17_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_25) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_17_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_17_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_17_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_17_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_17_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_17_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_218) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_17_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_17_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_17_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_17_ctrl_fcn_dw <= ~_GEN_218 & fb_uop_ram_17_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_17_ctrl_is_load <= ~_GEN_218 & fb_uop_ram_17_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_17_ctrl_is_sta <= ~_GEN_218 & fb_uop_ram_17_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_17_ctrl_is_std <= ~_GEN_218 & fb_uop_ram_17_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_17_iw_p1_poisoned <= ~_GEN_218 & fb_uop_ram_17_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_17_iw_p2_poisoned <= ~_GEN_218 & fb_uop_ram_17_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_17_edge_inst <=
      ~(_GEN_217 | _GEN_175 | _GEN_150)
      & (_GEN_125
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_100 | _GEN_75 | _GEN_50)
             & (_GEN_25 ? io_enq_bits_edge_inst_0 : fb_uop_ram_17_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_17_xcpt_ma_if <= ~_GEN_218 & fb_uop_ram_17_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_219) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_18_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_18_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_176) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_18_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_18_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_151) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_18_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_18_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_126) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_18_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_18_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_18_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_18_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_101) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_18_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_18_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_76) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_18_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_18_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_51) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_18_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_18_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_26) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_18_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_18_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_18_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_18_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_18_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_18_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_220) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_18_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_18_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_18_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_18_ctrl_fcn_dw <= ~_GEN_220 & fb_uop_ram_18_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_18_ctrl_is_load <= ~_GEN_220 & fb_uop_ram_18_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_18_ctrl_is_sta <= ~_GEN_220 & fb_uop_ram_18_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_18_ctrl_is_std <= ~_GEN_220 & fb_uop_ram_18_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_18_iw_p1_poisoned <= ~_GEN_220 & fb_uop_ram_18_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_18_iw_p2_poisoned <= ~_GEN_220 & fb_uop_ram_18_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_18_edge_inst <=
      ~(_GEN_219 | _GEN_176 | _GEN_151)
      & (_GEN_126
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_101 | _GEN_76 | _GEN_51)
             & (_GEN_26 ? io_enq_bits_edge_inst_0 : fb_uop_ram_18_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_18_xcpt_ma_if <= ~_GEN_220 & fb_uop_ram_18_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_221) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_19_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_19_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_177) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_19_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_19_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_152) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_19_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_19_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_127) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_19_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_19_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_19_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_19_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_102) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_19_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_19_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_77) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_19_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_19_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_52) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_19_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_19_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_27) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_19_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_19_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_19_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_19_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_19_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_19_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_222) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_19_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_19_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_19_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_19_ctrl_fcn_dw <= ~_GEN_222 & fb_uop_ram_19_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_19_ctrl_is_load <= ~_GEN_222 & fb_uop_ram_19_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_19_ctrl_is_sta <= ~_GEN_222 & fb_uop_ram_19_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_19_ctrl_is_std <= ~_GEN_222 & fb_uop_ram_19_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_19_iw_p1_poisoned <= ~_GEN_222 & fb_uop_ram_19_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_19_iw_p2_poisoned <= ~_GEN_222 & fb_uop_ram_19_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_19_edge_inst <=
      ~(_GEN_221 | _GEN_177 | _GEN_152)
      & (_GEN_127
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_102 | _GEN_77 | _GEN_52)
             & (_GEN_27 ? io_enq_bits_edge_inst_0 : fb_uop_ram_19_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_19_xcpt_ma_if <= ~_GEN_222 & fb_uop_ram_19_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_223) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_20_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_20_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_178) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_20_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_20_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_153) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_20_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_20_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_128) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_20_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_20_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_20_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_20_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_103) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_20_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_20_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_78) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_20_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_20_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_53) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_20_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_20_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_28) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_20_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_20_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_20_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_20_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_20_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_20_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_224) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_20_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_20_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_20_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_20_ctrl_fcn_dw <= ~_GEN_224 & fb_uop_ram_20_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_20_ctrl_is_load <= ~_GEN_224 & fb_uop_ram_20_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_20_ctrl_is_sta <= ~_GEN_224 & fb_uop_ram_20_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_20_ctrl_is_std <= ~_GEN_224 & fb_uop_ram_20_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_20_iw_p1_poisoned <= ~_GEN_224 & fb_uop_ram_20_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_20_iw_p2_poisoned <= ~_GEN_224 & fb_uop_ram_20_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_20_edge_inst <=
      ~(_GEN_223 | _GEN_178 | _GEN_153)
      & (_GEN_128
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_103 | _GEN_78 | _GEN_53)
             & (_GEN_28 ? io_enq_bits_edge_inst_0 : fb_uop_ram_20_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_20_xcpt_ma_if <= ~_GEN_224 & fb_uop_ram_20_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_225) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_21_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_21_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_179) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_21_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_21_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_154) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_21_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_21_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_129) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_21_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_21_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_21_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_21_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_104) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_21_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_21_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_79) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_21_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_21_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_54) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_21_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_21_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_29) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_21_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_21_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_21_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_21_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_21_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_21_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_226) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_21_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_21_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_21_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_21_ctrl_fcn_dw <= ~_GEN_226 & fb_uop_ram_21_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_21_ctrl_is_load <= ~_GEN_226 & fb_uop_ram_21_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_21_ctrl_is_sta <= ~_GEN_226 & fb_uop_ram_21_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_21_ctrl_is_std <= ~_GEN_226 & fb_uop_ram_21_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_21_iw_p1_poisoned <= ~_GEN_226 & fb_uop_ram_21_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_21_iw_p2_poisoned <= ~_GEN_226 & fb_uop_ram_21_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_21_edge_inst <=
      ~(_GEN_225 | _GEN_179 | _GEN_154)
      & (_GEN_129
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_104 | _GEN_79 | _GEN_54)
             & (_GEN_29 ? io_enq_bits_edge_inst_0 : fb_uop_ram_21_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_21_xcpt_ma_if <= ~_GEN_226 & fb_uop_ram_21_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_227) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_22_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_22_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_180) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_22_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_22_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_155) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_22_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_22_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_130) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_22_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_22_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_22_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_22_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_105) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_22_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_22_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_80) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_22_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_22_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_55) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_22_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_22_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_30) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_22_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_22_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_22_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_22_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_22_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_22_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_228) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_22_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_22_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_22_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_22_ctrl_fcn_dw <= ~_GEN_228 & fb_uop_ram_22_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_22_ctrl_is_load <= ~_GEN_228 & fb_uop_ram_22_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_22_ctrl_is_sta <= ~_GEN_228 & fb_uop_ram_22_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_22_ctrl_is_std <= ~_GEN_228 & fb_uop_ram_22_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_22_iw_p1_poisoned <= ~_GEN_228 & fb_uop_ram_22_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_22_iw_p2_poisoned <= ~_GEN_228 & fb_uop_ram_22_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_22_edge_inst <=
      ~(_GEN_227 | _GEN_180 | _GEN_155)
      & (_GEN_130
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_105 | _GEN_80 | _GEN_55)
             & (_GEN_30 ? io_enq_bits_edge_inst_0 : fb_uop_ram_22_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_22_xcpt_ma_if <= ~_GEN_228 & fb_uop_ram_22_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (_GEN_229) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_7_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_23_debug_pc <= _pc_T_31;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_pc_lob <= _pc_T_31[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_23_taken <= in_uops_7_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_7;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_7;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_181) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_6_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_23_debug_pc <= _pc_T_27;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_pc_lob <= _pc_T_27[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_23_taken <= in_uops_6_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_6;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_6;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_156) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_5_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_23_debug_pc <= _pc_T_23;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_pc_lob <= _pc_T_23[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_23_taken <= in_uops_5_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_5;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_5;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_131) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_4_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_1) begin
        fb_uop_ram_23_debug_pc <= _in_uops_4_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
        fb_uop_ram_23_pc_lob <= _in_uops_4_pc_lob_T_3;	// fetch-buffer.scala:57:16, :108:61
      end
      else begin
        fb_uop_ram_23_debug_pc <= _pc_T_19;	// fetch-buffer.scala:57:16, :95:43
        fb_uop_ram_23_pc_lob <= _pc_T_19[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      end
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_taken <= in_uops_4_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_4;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_4;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_106) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_3_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_23_debug_pc <= _pc_T_15;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_pc_lob <= _pc_T_15[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_23_taken <= in_uops_3_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_3;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_3;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_81) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_2_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_23_debug_pc <= _pc_T_11;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_pc_lob <= _pc_T_11[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_23_taken <= in_uops_2_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_2;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_2;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_56) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_1_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      fb_uop_ram_23_debug_pc <= _pc_T_7;	// fetch-buffer.scala:57:16, :95:43
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_pc_lob <= _pc_T_7[5:0];	// fetch-buffer.scala:57:16, :95:43, :101:33
      fb_uop_ram_23_taken <= in_uops_1_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_1;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_1;	// fetch-buffer.scala:57:16
    end
    else if (_GEN_31) begin	// fetch-buffer.scala:144:34
      fb_uop_ram_23_inst <= io_enq_bits_exp_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_inst <= io_enq_bits_insts_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_is_rvc <= in_uops_0_is_rvc;	// fetch-buffer.scala:57:16, :115:62
      if (io_enq_bits_edge_inst_0)
        fb_uop_ram_23_debug_pc <= _in_uops_0_debug_pc_T_5;	// fetch-buffer.scala:57:16, :107:81
      else
        fb_uop_ram_23_debug_pc <= pc;	// fetch-buffer.scala:57:16, frontend.scala:161:39
      fb_uop_ram_23_is_sfb <= io_enq_bits_shadowed_mask_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_pc_lob <= in_uops_0_pc_lob;	// fetch-buffer.scala:57:16, :101:33, :106:41, :108:32
      fb_uop_ram_23_taken <= in_uops_0_taken;	// fetch-buffer.scala:57:16, :116:69
      fb_uop_ram_23_bp_debug_if <= io_enq_bits_bp_debug_if_oh_0;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_bp_xcpt_if <= io_enq_bits_bp_xcpt_if_oh_0;	// fetch-buffer.scala:57:16
    end
    if (_GEN_230) begin	// fetch-buffer.scala:57:16, :144:53, :145:16
      fb_uop_ram_23_ctrl_br_type <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_ctrl_op1_sel <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_ctrl_op2_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_ctrl_imm_sel <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_ctrl_op_fcn <= 4'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_ctrl_csr_cmd <= 3'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_iw_state <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_ftq_idx <= io_enq_bits_ftq_idx;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_csr_addr <= 12'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_rxq_idx <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
      fb_uop_ram_23_xcpt_pf_if <= io_enq_bits_xcpt_pf_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_xcpt_ae_if <= io_enq_bits_xcpt_ae_if;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_fsrc <= io_enq_bits_fsrc;	// fetch-buffer.scala:57:16
      fb_uop_ram_23_debug_tsrc <= 2'h0;	// fetch-buffer.scala:57:16, :97:33
    end
    fb_uop_ram_23_ctrl_fcn_dw <= ~_GEN_230 & fb_uop_ram_23_ctrl_fcn_dw;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_23_ctrl_is_load <= ~_GEN_230 & fb_uop_ram_23_ctrl_is_load;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_23_ctrl_is_sta <= ~_GEN_230 & fb_uop_ram_23_ctrl_is_sta;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_23_ctrl_is_std <= ~_GEN_230 & fb_uop_ram_23_ctrl_is_std;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_23_iw_p1_poisoned <= ~_GEN_230 & fb_uop_ram_23_iw_p1_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_23_iw_p2_poisoned <= ~_GEN_230 & fb_uop_ram_23_iw_p2_poisoned;	// fetch-buffer.scala:57:16, :144:53, :145:16
    fb_uop_ram_23_edge_inst <=
      ~(_GEN_229 | _GEN_181 | _GEN_156)
      & (_GEN_131
           ? io_enq_bits_edge_inst_1
           : ~(_GEN_106 | _GEN_81 | _GEN_56)
             & (_GEN_31 ? io_enq_bits_edge_inst_0 : fb_uop_ram_23_edge_inst));	// fetch-buffer.scala:57:16, :144:{34,53}, :145:16
    fb_uop_ram_23_xcpt_ma_if <= ~_GEN_230 & fb_uop_ram_23_xcpt_ma_if;	// fetch-buffer.scala:57:16, :144:53, :145:16
    if (reset) begin
      head <= 8'h1;	// fetch-buffer.scala:61:21
      tail <= 24'h1;	// fetch-buffer.scala:62:21
      maybe_full <= 1'h0;	// fetch-buffer.scala:64:27
    end
    else begin
      automatic logic do_deq;	// fetch-buffer.scala:159:29
      do_deq = io_deq_ready & slot_will_hit_tail == 3'h0;	// fetch-buffer.scala:97:33, :156:112, :157:42, :159:29
      if (io_clear) begin
        head <= 8'h1;	// fetch-buffer.scala:61:21
        tail <= 24'h1;	// fetch-buffer.scala:62:21
      end
      else begin
        if (do_deq)	// fetch-buffer.scala:159:29
          head <= {head[6:0], head[7]};	// Cat.scala:30:58, fetch-buffer.scala:61:21, :132:12, :155:31
        if (~_do_enq_T_1) begin	// fetch-buffer.scala:82:40
          if (in_mask_7)	// fetch-buffer.scala:98:49
            tail <= {enq_idxs_7[22:0], enq_idxs_7[23]};	// Cat.scala:30:58, fetch-buffer.scala:62:21, :132:{12,24}, :138:18
          else if (in_mask_6)	// fetch-buffer.scala:98:49
            tail <= _GEN_6;	// Cat.scala:30:58, fetch-buffer.scala:62:21
          else if (in_mask_5)	// fetch-buffer.scala:98:49
            tail <= _GEN_5;	// Cat.scala:30:58, fetch-buffer.scala:62:21
          else if (in_mask_4)	// fetch-buffer.scala:98:49
            tail <= _GEN_4;	// Cat.scala:30:58, fetch-buffer.scala:62:21
          else if (in_mask_3)	// fetch-buffer.scala:98:49
            tail <= _GEN_3;	// Cat.scala:30:58, fetch-buffer.scala:62:21
          else if (in_mask_2)	// fetch-buffer.scala:98:49
            tail <= _GEN_2;	// Cat.scala:30:58, fetch-buffer.scala:62:21
          else if (in_mask_1)	// fetch-buffer.scala:98:49
            tail <= _GEN_1;	// Cat.scala:30:58, fetch-buffer.scala:62:21
          else if (in_mask_0)	// fetch-buffer.scala:98:49
            tail <= _GEN_0;	// Cat.scala:30:58, fetch-buffer.scala:62:21
        end
      end
      maybe_full <=
        ~(io_clear | do_deq)
        & (~_do_enq_T_1
           & (in_mask_0 | in_mask_1 | in_mask_2 | in_mask_3 | in_mask_4 | in_mask_5
              | in_mask_6 | in_mask_7) | maybe_full);	// fetch-buffer.scala:64:27, :82:{16,40}, :98:49, :159:29, :176:17, :178:{27,33}, :179:18, :183:17, :185:16, :188:19, :191:16
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:308];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [8:0] i = 9'h0; i < 9'h135; i += 9'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        fb_uop_ram_0_inst = {_RANDOM[9'h0][31:7], _RANDOM[9'h1][6:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_0_debug_inst = {_RANDOM[9'h1][31:7], _RANDOM[9'h2][6:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_0_is_rvc = _RANDOM[9'h2][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_debug_pc = {_RANDOM[9'h2][31:8], _RANDOM[9'h3][15:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_br_type = {_RANDOM[9'h3][31:29], _RANDOM[9'h4][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_op1_sel = _RANDOM[9'h4][2:1];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_op2_sel = _RANDOM[9'h4][5:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_imm_sel = _RANDOM[9'h4][8:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_op_fcn = _RANDOM[9'h4][12:9];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_fcn_dw = _RANDOM[9'h4][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_csr_cmd = _RANDOM[9'h4][16:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_is_load = _RANDOM[9'h4][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_is_sta = _RANDOM[9'h4][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ctrl_is_std = _RANDOM[9'h4][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_iw_state = _RANDOM[9'h4][21:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_iw_p1_poisoned = _RANDOM[9'h4][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_iw_p2_poisoned = _RANDOM[9'h4][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_is_sfb = _RANDOM[9'h4][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_ftq_idx = _RANDOM[9'h5][20:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_edge_inst = _RANDOM[9'h5][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_pc_lob = _RANDOM[9'h5][27:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_taken = _RANDOM[9'h5][28];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_csr_addr = _RANDOM[9'h6][28:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_rxq_idx = _RANDOM[9'h7][15:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_xcpt_pf_if = _RANDOM[9'hC][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_xcpt_ae_if = _RANDOM[9'hC][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_xcpt_ma_if = _RANDOM[9'hC][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_bp_debug_if = _RANDOM[9'hC][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_bp_xcpt_if = _RANDOM[9'hC][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_debug_fsrc = _RANDOM[9'hC][23:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_0_debug_tsrc = _RANDOM[9'hC][25:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_inst = {_RANDOM[9'hD][31:1], _RANDOM[9'hE][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_1_debug_inst = {_RANDOM[9'hE][31:1], _RANDOM[9'hF][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_1_is_rvc = _RANDOM[9'hF][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_debug_pc = {_RANDOM[9'hF][31:2], _RANDOM[9'h10][9:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_br_type = _RANDOM[9'h10][26:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_op1_sel = _RANDOM[9'h10][28:27];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_op2_sel = _RANDOM[9'h10][31:29];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_imm_sel = _RANDOM[9'h11][2:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_op_fcn = _RANDOM[9'h11][6:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_fcn_dw = _RANDOM[9'h11][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_csr_cmd = _RANDOM[9'h11][10:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_is_load = _RANDOM[9'h11][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_is_sta = _RANDOM[9'h11][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ctrl_is_std = _RANDOM[9'h11][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_iw_state = _RANDOM[9'h11][15:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_iw_p1_poisoned = _RANDOM[9'h11][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_iw_p2_poisoned = _RANDOM[9'h11][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_is_sfb = _RANDOM[9'h11][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_ftq_idx = _RANDOM[9'h12][14:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_edge_inst = _RANDOM[9'h12][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_pc_lob = _RANDOM[9'h12][21:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_taken = _RANDOM[9'h12][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_csr_addr = _RANDOM[9'h13][22:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_rxq_idx = _RANDOM[9'h14][9:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_xcpt_pf_if = _RANDOM[9'h19][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_xcpt_ae_if = _RANDOM[9'h19][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_xcpt_ma_if = _RANDOM[9'h19][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_bp_debug_if = _RANDOM[9'h19][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_bp_xcpt_if = _RANDOM[9'h19][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_debug_fsrc = _RANDOM[9'h19][17:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_1_debug_tsrc = _RANDOM[9'h19][19:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_inst = {_RANDOM[9'h19][31:27], _RANDOM[9'h1A][26:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_2_debug_inst = {_RANDOM[9'h1A][31:27], _RANDOM[9'h1B][26:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_2_is_rvc = _RANDOM[9'h1B][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_debug_pc =
          {_RANDOM[9'h1B][31:28], _RANDOM[9'h1C], _RANDOM[9'h1D][3:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_br_type = _RANDOM[9'h1D][20:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_op1_sel = _RANDOM[9'h1D][22:21];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_op2_sel = _RANDOM[9'h1D][25:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_imm_sel = _RANDOM[9'h1D][28:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_op_fcn = {_RANDOM[9'h1D][31:29], _RANDOM[9'h1E][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_fcn_dw = _RANDOM[9'h1E][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_csr_cmd = _RANDOM[9'h1E][4:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_is_load = _RANDOM[9'h1E][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_is_sta = _RANDOM[9'h1E][6];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ctrl_is_std = _RANDOM[9'h1E][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_iw_state = _RANDOM[9'h1E][9:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_iw_p1_poisoned = _RANDOM[9'h1E][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_iw_p2_poisoned = _RANDOM[9'h1E][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_is_sfb = _RANDOM[9'h1E][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_ftq_idx = _RANDOM[9'h1F][8:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_edge_inst = _RANDOM[9'h1F][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_pc_lob = _RANDOM[9'h1F][15:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_taken = _RANDOM[9'h1F][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_csr_addr = _RANDOM[9'h20][16:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_rxq_idx = _RANDOM[9'h21][3:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_xcpt_pf_if = _RANDOM[9'h26][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_xcpt_ae_if = _RANDOM[9'h26][6];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_xcpt_ma_if = _RANDOM[9'h26][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_bp_debug_if = _RANDOM[9'h26][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_bp_xcpt_if = _RANDOM[9'h26][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_debug_fsrc = _RANDOM[9'h26][11:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_2_debug_tsrc = _RANDOM[9'h26][13:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_inst = {_RANDOM[9'h26][31:21], _RANDOM[9'h27][20:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_3_debug_inst = {_RANDOM[9'h27][31:21], _RANDOM[9'h28][20:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_3_is_rvc = _RANDOM[9'h28][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_debug_pc = {_RANDOM[9'h28][31:22], _RANDOM[9'h29][29:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_br_type = _RANDOM[9'h2A][14:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_op1_sel = _RANDOM[9'h2A][16:15];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_op2_sel = _RANDOM[9'h2A][19:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_imm_sel = _RANDOM[9'h2A][22:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_op_fcn = _RANDOM[9'h2A][26:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_fcn_dw = _RANDOM[9'h2A][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_csr_cmd = _RANDOM[9'h2A][30:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_is_load = _RANDOM[9'h2A][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_is_sta = _RANDOM[9'h2B][0];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ctrl_is_std = _RANDOM[9'h2B][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_iw_state = _RANDOM[9'h2B][3:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_iw_p1_poisoned = _RANDOM[9'h2B][4];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_iw_p2_poisoned = _RANDOM[9'h2B][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_is_sfb = _RANDOM[9'h2B][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_ftq_idx = {_RANDOM[9'h2B][31:30], _RANDOM[9'h2C][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_3_edge_inst = _RANDOM[9'h2C][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_pc_lob = _RANDOM[9'h2C][9:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_taken = _RANDOM[9'h2C][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_csr_addr = {_RANDOM[9'h2C][31], _RANDOM[9'h2D][10:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_3_rxq_idx = _RANDOM[9'h2D][29:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_xcpt_pf_if = _RANDOM[9'h32][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_xcpt_ae_if = _RANDOM[9'h33][0];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_xcpt_ma_if = _RANDOM[9'h33][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_bp_debug_if = _RANDOM[9'h33][2];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_bp_xcpt_if = _RANDOM[9'h33][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_debug_fsrc = _RANDOM[9'h33][5:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_3_debug_tsrc = _RANDOM[9'h33][7:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_inst = {_RANDOM[9'h33][31:15], _RANDOM[9'h34][14:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_4_debug_inst = {_RANDOM[9'h34][31:15], _RANDOM[9'h35][14:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_4_is_rvc = _RANDOM[9'h35][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_debug_pc = {_RANDOM[9'h35][31:16], _RANDOM[9'h36][23:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_br_type = _RANDOM[9'h37][8:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_op1_sel = _RANDOM[9'h37][10:9];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_op2_sel = _RANDOM[9'h37][13:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_imm_sel = _RANDOM[9'h37][16:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_op_fcn = _RANDOM[9'h37][20:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_fcn_dw = _RANDOM[9'h37][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_csr_cmd = _RANDOM[9'h37][24:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_is_load = _RANDOM[9'h37][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_is_sta = _RANDOM[9'h37][26];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ctrl_is_std = _RANDOM[9'h37][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_iw_state = _RANDOM[9'h37][29:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_iw_p1_poisoned = _RANDOM[9'h37][30];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_iw_p2_poisoned = _RANDOM[9'h37][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_is_sfb = _RANDOM[9'h38][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_ftq_idx = _RANDOM[9'h38][28:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_edge_inst = _RANDOM[9'h38][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_pc_lob = {_RANDOM[9'h38][31:30], _RANDOM[9'h39][3:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_4_taken = _RANDOM[9'h39][4];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_csr_addr = {_RANDOM[9'h39][31:25], _RANDOM[9'h3A][4:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_4_rxq_idx = _RANDOM[9'h3A][23:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_xcpt_pf_if = _RANDOM[9'h3F][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_xcpt_ae_if = _RANDOM[9'h3F][26];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_xcpt_ma_if = _RANDOM[9'h3F][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_bp_debug_if = _RANDOM[9'h3F][28];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_bp_xcpt_if = _RANDOM[9'h3F][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_debug_fsrc = _RANDOM[9'h3F][31:30];	// fetch-buffer.scala:57:16
        fb_uop_ram_4_debug_tsrc = _RANDOM[9'h40][1:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_inst = {_RANDOM[9'h40][31:9], _RANDOM[9'h41][8:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_5_debug_inst = {_RANDOM[9'h41][31:9], _RANDOM[9'h42][8:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_5_is_rvc = _RANDOM[9'h42][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_debug_pc = {_RANDOM[9'h42][31:10], _RANDOM[9'h43][17:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_br_type = {_RANDOM[9'h43][31], _RANDOM[9'h44][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_op1_sel = _RANDOM[9'h44][4:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_op2_sel = _RANDOM[9'h44][7:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_imm_sel = _RANDOM[9'h44][10:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_op_fcn = _RANDOM[9'h44][14:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_fcn_dw = _RANDOM[9'h44][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_csr_cmd = _RANDOM[9'h44][18:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_is_load = _RANDOM[9'h44][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_is_sta = _RANDOM[9'h44][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ctrl_is_std = _RANDOM[9'h44][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_iw_state = _RANDOM[9'h44][23:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_iw_p1_poisoned = _RANDOM[9'h44][24];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_iw_p2_poisoned = _RANDOM[9'h44][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_is_sfb = _RANDOM[9'h44][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_ftq_idx = _RANDOM[9'h45][22:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_edge_inst = _RANDOM[9'h45][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_pc_lob = _RANDOM[9'h45][29:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_taken = _RANDOM[9'h45][30];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_csr_addr = _RANDOM[9'h46][30:19];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_rxq_idx = _RANDOM[9'h47][17:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_xcpt_pf_if = _RANDOM[9'h4C][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_xcpt_ae_if = _RANDOM[9'h4C][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_xcpt_ma_if = _RANDOM[9'h4C][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_bp_debug_if = _RANDOM[9'h4C][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_bp_xcpt_if = _RANDOM[9'h4C][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_debug_fsrc = _RANDOM[9'h4C][25:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_5_debug_tsrc = _RANDOM[9'h4C][27:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_inst = {_RANDOM[9'h4D][31:3], _RANDOM[9'h4E][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_6_debug_inst = {_RANDOM[9'h4E][31:3], _RANDOM[9'h4F][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_6_is_rvc = _RANDOM[9'h4F][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_debug_pc = {_RANDOM[9'h4F][31:4], _RANDOM[9'h50][11:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_br_type = _RANDOM[9'h50][28:25];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_op1_sel = _RANDOM[9'h50][30:29];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_op2_sel = {_RANDOM[9'h50][31], _RANDOM[9'h51][1:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_imm_sel = _RANDOM[9'h51][4:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_op_fcn = _RANDOM[9'h51][8:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_fcn_dw = _RANDOM[9'h51][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_csr_cmd = _RANDOM[9'h51][12:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_is_load = _RANDOM[9'h51][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_is_sta = _RANDOM[9'h51][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ctrl_is_std = _RANDOM[9'h51][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_iw_state = _RANDOM[9'h51][17:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_iw_p1_poisoned = _RANDOM[9'h51][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_iw_p2_poisoned = _RANDOM[9'h51][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_is_sfb = _RANDOM[9'h51][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_ftq_idx = _RANDOM[9'h52][16:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_edge_inst = _RANDOM[9'h52][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_pc_lob = _RANDOM[9'h52][23:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_taken = _RANDOM[9'h52][24];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_csr_addr = _RANDOM[9'h53][24:13];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_rxq_idx = _RANDOM[9'h54][11:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_xcpt_pf_if = _RANDOM[9'h59][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_xcpt_ae_if = _RANDOM[9'h59][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_xcpt_ma_if = _RANDOM[9'h59][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_bp_debug_if = _RANDOM[9'h59][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_bp_xcpt_if = _RANDOM[9'h59][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_debug_fsrc = _RANDOM[9'h59][19:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_6_debug_tsrc = _RANDOM[9'h59][21:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_inst = {_RANDOM[9'h59][31:29], _RANDOM[9'h5A][28:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_7_debug_inst = {_RANDOM[9'h5A][31:29], _RANDOM[9'h5B][28:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_7_is_rvc = _RANDOM[9'h5B][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_debug_pc =
          {_RANDOM[9'h5B][31:30], _RANDOM[9'h5C], _RANDOM[9'h5D][5:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_br_type = _RANDOM[9'h5D][22:19];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_op1_sel = _RANDOM[9'h5D][24:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_op2_sel = _RANDOM[9'h5D][27:25];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_imm_sel = _RANDOM[9'h5D][30:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_op_fcn = {_RANDOM[9'h5D][31], _RANDOM[9'h5E][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_fcn_dw = _RANDOM[9'h5E][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_csr_cmd = _RANDOM[9'h5E][6:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_is_load = _RANDOM[9'h5E][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_is_sta = _RANDOM[9'h5E][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ctrl_is_std = _RANDOM[9'h5E][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_iw_state = _RANDOM[9'h5E][11:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_iw_p1_poisoned = _RANDOM[9'h5E][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_iw_p2_poisoned = _RANDOM[9'h5E][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_is_sfb = _RANDOM[9'h5E][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_ftq_idx = _RANDOM[9'h5F][10:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_edge_inst = _RANDOM[9'h5F][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_pc_lob = _RANDOM[9'h5F][17:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_taken = _RANDOM[9'h5F][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_csr_addr = _RANDOM[9'h60][18:7];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_rxq_idx = _RANDOM[9'h61][5:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_xcpt_pf_if = _RANDOM[9'h66][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_xcpt_ae_if = _RANDOM[9'h66][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_xcpt_ma_if = _RANDOM[9'h66][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_bp_debug_if = _RANDOM[9'h66][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_bp_xcpt_if = _RANDOM[9'h66][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_debug_fsrc = _RANDOM[9'h66][13:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_7_debug_tsrc = _RANDOM[9'h66][15:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_inst = {_RANDOM[9'h66][31:23], _RANDOM[9'h67][22:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_8_debug_inst = {_RANDOM[9'h67][31:23], _RANDOM[9'h68][22:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_8_is_rvc = _RANDOM[9'h68][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_debug_pc = {_RANDOM[9'h68][31:24], _RANDOM[9'h69]};	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_br_type = _RANDOM[9'h6A][16:13];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_op1_sel = _RANDOM[9'h6A][18:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_op2_sel = _RANDOM[9'h6A][21:19];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_imm_sel = _RANDOM[9'h6A][24:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_op_fcn = _RANDOM[9'h6A][28:25];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_fcn_dw = _RANDOM[9'h6A][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_csr_cmd = {_RANDOM[9'h6A][31:30], _RANDOM[9'h6B][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_is_load = _RANDOM[9'h6B][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_is_sta = _RANDOM[9'h6B][2];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ctrl_is_std = _RANDOM[9'h6B][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_iw_state = _RANDOM[9'h6B][5:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_iw_p1_poisoned = _RANDOM[9'h6B][6];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_iw_p2_poisoned = _RANDOM[9'h6B][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_is_sfb = _RANDOM[9'h6B][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_ftq_idx = _RANDOM[9'h6C][4:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_edge_inst = _RANDOM[9'h6C][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_pc_lob = _RANDOM[9'h6C][11:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_taken = _RANDOM[9'h6C][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_csr_addr = _RANDOM[9'h6D][12:1];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_rxq_idx = _RANDOM[9'h6D][31:30];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_xcpt_pf_if = _RANDOM[9'h73][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_xcpt_ae_if = _RANDOM[9'h73][2];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_xcpt_ma_if = _RANDOM[9'h73][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_bp_debug_if = _RANDOM[9'h73][4];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_bp_xcpt_if = _RANDOM[9'h73][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_debug_fsrc = _RANDOM[9'h73][7:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_8_debug_tsrc = _RANDOM[9'h73][9:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_inst = {_RANDOM[9'h73][31:17], _RANDOM[9'h74][16:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_9_debug_inst = {_RANDOM[9'h74][31:17], _RANDOM[9'h75][16:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_9_is_rvc = _RANDOM[9'h75][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_debug_pc = {_RANDOM[9'h75][31:18], _RANDOM[9'h76][25:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_br_type = _RANDOM[9'h77][10:7];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_op1_sel = _RANDOM[9'h77][12:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_op2_sel = _RANDOM[9'h77][15:13];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_imm_sel = _RANDOM[9'h77][18:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_op_fcn = _RANDOM[9'h77][22:19];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_fcn_dw = _RANDOM[9'h77][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_csr_cmd = _RANDOM[9'h77][26:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_is_load = _RANDOM[9'h77][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_is_sta = _RANDOM[9'h77][28];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ctrl_is_std = _RANDOM[9'h77][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_iw_state = _RANDOM[9'h77][31:30];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_iw_p1_poisoned = _RANDOM[9'h78][0];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_iw_p2_poisoned = _RANDOM[9'h78][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_is_sfb = _RANDOM[9'h78][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_ftq_idx = _RANDOM[9'h78][30:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_edge_inst = _RANDOM[9'h78][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_pc_lob = _RANDOM[9'h79][5:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_taken = _RANDOM[9'h79][6];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_csr_addr = {_RANDOM[9'h79][31:27], _RANDOM[9'h7A][6:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_9_rxq_idx = _RANDOM[9'h7A][25:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_xcpt_pf_if = _RANDOM[9'h7F][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_xcpt_ae_if = _RANDOM[9'h7F][28];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_xcpt_ma_if = _RANDOM[9'h7F][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_bp_debug_if = _RANDOM[9'h7F][30];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_bp_xcpt_if = _RANDOM[9'h7F][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_debug_fsrc = _RANDOM[9'h80][1:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_9_debug_tsrc = _RANDOM[9'h80][3:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_inst = {_RANDOM[9'h80][31:11], _RANDOM[9'h81][10:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_10_debug_inst = {_RANDOM[9'h81][31:11], _RANDOM[9'h82][10:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_10_is_rvc = _RANDOM[9'h82][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_debug_pc = {_RANDOM[9'h82][31:12], _RANDOM[9'h83][19:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_br_type = _RANDOM[9'h84][4:1];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_op1_sel = _RANDOM[9'h84][6:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_op2_sel = _RANDOM[9'h84][9:7];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_imm_sel = _RANDOM[9'h84][12:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_op_fcn = _RANDOM[9'h84][16:13];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_fcn_dw = _RANDOM[9'h84][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_csr_cmd = _RANDOM[9'h84][20:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_is_load = _RANDOM[9'h84][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_is_sta = _RANDOM[9'h84][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ctrl_is_std = _RANDOM[9'h84][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_iw_state = _RANDOM[9'h84][25:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_iw_p1_poisoned = _RANDOM[9'h84][26];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_iw_p2_poisoned = _RANDOM[9'h84][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_is_sfb = _RANDOM[9'h84][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_ftq_idx = _RANDOM[9'h85][24:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_edge_inst = _RANDOM[9'h85][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_pc_lob = _RANDOM[9'h85][31:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_taken = _RANDOM[9'h86][0];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_csr_addr = {_RANDOM[9'h86][31:21], _RANDOM[9'h87][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_10_rxq_idx = _RANDOM[9'h87][19:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_xcpt_pf_if = _RANDOM[9'h8C][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_xcpt_ae_if = _RANDOM[9'h8C][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_xcpt_ma_if = _RANDOM[9'h8C][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_bp_debug_if = _RANDOM[9'h8C][24];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_bp_xcpt_if = _RANDOM[9'h8C][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_debug_fsrc = _RANDOM[9'h8C][27:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_10_debug_tsrc = _RANDOM[9'h8C][29:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_inst = {_RANDOM[9'h8D][31:5], _RANDOM[9'h8E][4:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_11_debug_inst = {_RANDOM[9'h8E][31:5], _RANDOM[9'h8F][4:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_11_is_rvc = _RANDOM[9'h8F][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_debug_pc = {_RANDOM[9'h8F][31:6], _RANDOM[9'h90][13:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_br_type = _RANDOM[9'h90][30:27];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_op1_sel = {_RANDOM[9'h90][31], _RANDOM[9'h91][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_op2_sel = _RANDOM[9'h91][3:1];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_imm_sel = _RANDOM[9'h91][6:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_op_fcn = _RANDOM[9'h91][10:7];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_fcn_dw = _RANDOM[9'h91][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_csr_cmd = _RANDOM[9'h91][14:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_is_load = _RANDOM[9'h91][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_is_sta = _RANDOM[9'h91][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ctrl_is_std = _RANDOM[9'h91][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_iw_state = _RANDOM[9'h91][19:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_iw_p1_poisoned = _RANDOM[9'h91][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_iw_p2_poisoned = _RANDOM[9'h91][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_is_sfb = _RANDOM[9'h91][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_ftq_idx = _RANDOM[9'h92][18:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_edge_inst = _RANDOM[9'h92][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_pc_lob = _RANDOM[9'h92][25:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_taken = _RANDOM[9'h92][26];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_csr_addr = _RANDOM[9'h93][26:15];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_rxq_idx = _RANDOM[9'h94][13:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_xcpt_pf_if = _RANDOM[9'h99][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_xcpt_ae_if = _RANDOM[9'h99][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_xcpt_ma_if = _RANDOM[9'h99][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_bp_debug_if = _RANDOM[9'h99][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_bp_xcpt_if = _RANDOM[9'h99][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_debug_fsrc = _RANDOM[9'h99][21:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_11_debug_tsrc = _RANDOM[9'h99][23:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_inst = {_RANDOM[9'h99][31], _RANDOM[9'h9A][30:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_12_debug_inst = {_RANDOM[9'h9A][31], _RANDOM[9'h9B][30:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_12_is_rvc = _RANDOM[9'h9B][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_debug_pc = {_RANDOM[9'h9C], _RANDOM[9'h9D][7:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_br_type = _RANDOM[9'h9D][24:21];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_op1_sel = _RANDOM[9'h9D][26:25];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_op2_sel = _RANDOM[9'h9D][29:27];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_imm_sel = {_RANDOM[9'h9D][31:30], _RANDOM[9'h9E][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_op_fcn = _RANDOM[9'h9E][4:1];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_fcn_dw = _RANDOM[9'h9E][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_csr_cmd = _RANDOM[9'h9E][8:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_is_load = _RANDOM[9'h9E][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_is_sta = _RANDOM[9'h9E][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ctrl_is_std = _RANDOM[9'h9E][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_iw_state = _RANDOM[9'h9E][13:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_iw_p1_poisoned = _RANDOM[9'h9E][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_iw_p2_poisoned = _RANDOM[9'h9E][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_is_sfb = _RANDOM[9'h9E][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_ftq_idx = _RANDOM[9'h9F][12:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_edge_inst = _RANDOM[9'h9F][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_pc_lob = _RANDOM[9'h9F][19:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_taken = _RANDOM[9'h9F][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_csr_addr = _RANDOM[9'hA0][20:9];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_rxq_idx = _RANDOM[9'hA1][7:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_xcpt_pf_if = _RANDOM[9'hA6][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_xcpt_ae_if = _RANDOM[9'hA6][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_xcpt_ma_if = _RANDOM[9'hA6][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_bp_debug_if = _RANDOM[9'hA6][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_bp_xcpt_if = _RANDOM[9'hA6][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_debug_fsrc = _RANDOM[9'hA6][15:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_12_debug_tsrc = _RANDOM[9'hA6][17:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_inst = {_RANDOM[9'hA6][31:25], _RANDOM[9'hA7][24:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_13_debug_inst = {_RANDOM[9'hA7][31:25], _RANDOM[9'hA8][24:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_13_is_rvc = _RANDOM[9'hA8][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_debug_pc =
          {_RANDOM[9'hA8][31:26], _RANDOM[9'hA9], _RANDOM[9'hAA][1:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_br_type = _RANDOM[9'hAA][18:15];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_op1_sel = _RANDOM[9'hAA][20:19];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_op2_sel = _RANDOM[9'hAA][23:21];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_imm_sel = _RANDOM[9'hAA][26:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_op_fcn = _RANDOM[9'hAA][30:27];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_fcn_dw = _RANDOM[9'hAA][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_csr_cmd = _RANDOM[9'hAB][2:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_is_load = _RANDOM[9'hAB][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_is_sta = _RANDOM[9'hAB][4];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ctrl_is_std = _RANDOM[9'hAB][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_iw_state = _RANDOM[9'hAB][7:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_iw_p1_poisoned = _RANDOM[9'hAB][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_iw_p2_poisoned = _RANDOM[9'hAB][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_is_sfb = _RANDOM[9'hAB][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_ftq_idx = _RANDOM[9'hAC][6:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_edge_inst = _RANDOM[9'hAC][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_pc_lob = _RANDOM[9'hAC][13:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_taken = _RANDOM[9'hAC][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_csr_addr = _RANDOM[9'hAD][14:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_rxq_idx = _RANDOM[9'hAE][1:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_xcpt_pf_if = _RANDOM[9'hB3][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_xcpt_ae_if = _RANDOM[9'hB3][4];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_xcpt_ma_if = _RANDOM[9'hB3][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_bp_debug_if = _RANDOM[9'hB3][6];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_bp_xcpt_if = _RANDOM[9'hB3][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_debug_fsrc = _RANDOM[9'hB3][9:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_13_debug_tsrc = _RANDOM[9'hB3][11:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_inst = {_RANDOM[9'hB3][31:19], _RANDOM[9'hB4][18:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_14_debug_inst = {_RANDOM[9'hB4][31:19], _RANDOM[9'hB5][18:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_14_is_rvc = _RANDOM[9'hB5][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_debug_pc = {_RANDOM[9'hB5][31:20], _RANDOM[9'hB6][27:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_br_type = _RANDOM[9'hB7][12:9];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_op1_sel = _RANDOM[9'hB7][14:13];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_op2_sel = _RANDOM[9'hB7][17:15];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_imm_sel = _RANDOM[9'hB7][20:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_op_fcn = _RANDOM[9'hB7][24:21];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_fcn_dw = _RANDOM[9'hB7][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_csr_cmd = _RANDOM[9'hB7][28:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_is_load = _RANDOM[9'hB7][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_is_sta = _RANDOM[9'hB7][30];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ctrl_is_std = _RANDOM[9'hB7][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_iw_state = _RANDOM[9'hB8][1:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_iw_p1_poisoned = _RANDOM[9'hB8][2];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_iw_p2_poisoned = _RANDOM[9'hB8][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_is_sfb = _RANDOM[9'hB8][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_ftq_idx = {_RANDOM[9'hB8][31:28], _RANDOM[9'hB9][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_14_edge_inst = _RANDOM[9'hB9][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_pc_lob = _RANDOM[9'hB9][7:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_taken = _RANDOM[9'hB9][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_csr_addr = {_RANDOM[9'hB9][31:29], _RANDOM[9'hBA][8:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_14_rxq_idx = _RANDOM[9'hBA][27:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_xcpt_pf_if = _RANDOM[9'hBF][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_xcpt_ae_if = _RANDOM[9'hBF][30];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_xcpt_ma_if = _RANDOM[9'hBF][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_bp_debug_if = _RANDOM[9'hC0][0];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_bp_xcpt_if = _RANDOM[9'hC0][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_debug_fsrc = _RANDOM[9'hC0][3:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_14_debug_tsrc = _RANDOM[9'hC0][5:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_inst = {_RANDOM[9'hC0][31:13], _RANDOM[9'hC1][12:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_15_debug_inst = {_RANDOM[9'hC1][31:13], _RANDOM[9'hC2][12:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_15_is_rvc = _RANDOM[9'hC2][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_debug_pc = {_RANDOM[9'hC2][31:14], _RANDOM[9'hC3][21:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_br_type = _RANDOM[9'hC4][6:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_op1_sel = _RANDOM[9'hC4][8:7];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_op2_sel = _RANDOM[9'hC4][11:9];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_imm_sel = _RANDOM[9'hC4][14:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_op_fcn = _RANDOM[9'hC4][18:15];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_fcn_dw = _RANDOM[9'hC4][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_csr_cmd = _RANDOM[9'hC4][22:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_is_load = _RANDOM[9'hC4][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_is_sta = _RANDOM[9'hC4][24];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ctrl_is_std = _RANDOM[9'hC4][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_iw_state = _RANDOM[9'hC4][27:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_iw_p1_poisoned = _RANDOM[9'hC4][28];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_iw_p2_poisoned = _RANDOM[9'hC4][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_is_sfb = _RANDOM[9'hC5][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_ftq_idx = _RANDOM[9'hC5][26:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_edge_inst = _RANDOM[9'hC5][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_pc_lob = {_RANDOM[9'hC5][31:28], _RANDOM[9'hC6][1:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_15_taken = _RANDOM[9'hC6][2];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_csr_addr = {_RANDOM[9'hC6][31:23], _RANDOM[9'hC7][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_15_rxq_idx = _RANDOM[9'hC7][21:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_xcpt_pf_if = _RANDOM[9'hCC][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_xcpt_ae_if = _RANDOM[9'hCC][24];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_xcpt_ma_if = _RANDOM[9'hCC][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_bp_debug_if = _RANDOM[9'hCC][26];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_bp_xcpt_if = _RANDOM[9'hCC][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_debug_fsrc = _RANDOM[9'hCC][29:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_15_debug_tsrc = _RANDOM[9'hCC][31:30];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_inst = {_RANDOM[9'hCD][31:7], _RANDOM[9'hCE][6:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_16_debug_inst = {_RANDOM[9'hCE][31:7], _RANDOM[9'hCF][6:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_16_is_rvc = _RANDOM[9'hCF][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_debug_pc = {_RANDOM[9'hCF][31:8], _RANDOM[9'hD0][15:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_br_type = {_RANDOM[9'hD0][31:29], _RANDOM[9'hD1][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_op1_sel = _RANDOM[9'hD1][2:1];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_op2_sel = _RANDOM[9'hD1][5:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_imm_sel = _RANDOM[9'hD1][8:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_op_fcn = _RANDOM[9'hD1][12:9];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_fcn_dw = _RANDOM[9'hD1][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_csr_cmd = _RANDOM[9'hD1][16:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_is_load = _RANDOM[9'hD1][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_is_sta = _RANDOM[9'hD1][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ctrl_is_std = _RANDOM[9'hD1][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_iw_state = _RANDOM[9'hD1][21:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_iw_p1_poisoned = _RANDOM[9'hD1][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_iw_p2_poisoned = _RANDOM[9'hD1][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_is_sfb = _RANDOM[9'hD1][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_ftq_idx = _RANDOM[9'hD2][20:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_edge_inst = _RANDOM[9'hD2][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_pc_lob = _RANDOM[9'hD2][27:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_taken = _RANDOM[9'hD2][28];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_csr_addr = _RANDOM[9'hD3][28:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_rxq_idx = _RANDOM[9'hD4][15:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_xcpt_pf_if = _RANDOM[9'hD9][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_xcpt_ae_if = _RANDOM[9'hD9][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_xcpt_ma_if = _RANDOM[9'hD9][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_bp_debug_if = _RANDOM[9'hD9][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_bp_xcpt_if = _RANDOM[9'hD9][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_debug_fsrc = _RANDOM[9'hD9][23:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_16_debug_tsrc = _RANDOM[9'hD9][25:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_inst = {_RANDOM[9'hDA][31:1], _RANDOM[9'hDB][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_17_debug_inst = {_RANDOM[9'hDB][31:1], _RANDOM[9'hDC][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_17_is_rvc = _RANDOM[9'hDC][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_debug_pc = {_RANDOM[9'hDC][31:2], _RANDOM[9'hDD][9:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_br_type = _RANDOM[9'hDD][26:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_op1_sel = _RANDOM[9'hDD][28:27];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_op2_sel = _RANDOM[9'hDD][31:29];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_imm_sel = _RANDOM[9'hDE][2:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_op_fcn = _RANDOM[9'hDE][6:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_fcn_dw = _RANDOM[9'hDE][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_csr_cmd = _RANDOM[9'hDE][10:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_is_load = _RANDOM[9'hDE][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_is_sta = _RANDOM[9'hDE][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ctrl_is_std = _RANDOM[9'hDE][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_iw_state = _RANDOM[9'hDE][15:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_iw_p1_poisoned = _RANDOM[9'hDE][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_iw_p2_poisoned = _RANDOM[9'hDE][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_is_sfb = _RANDOM[9'hDE][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_ftq_idx = _RANDOM[9'hDF][14:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_edge_inst = _RANDOM[9'hDF][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_pc_lob = _RANDOM[9'hDF][21:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_taken = _RANDOM[9'hDF][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_csr_addr = _RANDOM[9'hE0][22:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_rxq_idx = _RANDOM[9'hE1][9:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_xcpt_pf_if = _RANDOM[9'hE6][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_xcpt_ae_if = _RANDOM[9'hE6][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_xcpt_ma_if = _RANDOM[9'hE6][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_bp_debug_if = _RANDOM[9'hE6][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_bp_xcpt_if = _RANDOM[9'hE6][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_debug_fsrc = _RANDOM[9'hE6][17:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_17_debug_tsrc = _RANDOM[9'hE6][19:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_inst = {_RANDOM[9'hE6][31:27], _RANDOM[9'hE7][26:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_18_debug_inst = {_RANDOM[9'hE7][31:27], _RANDOM[9'hE8][26:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_18_is_rvc = _RANDOM[9'hE8][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_debug_pc =
          {_RANDOM[9'hE8][31:28], _RANDOM[9'hE9], _RANDOM[9'hEA][3:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_br_type = _RANDOM[9'hEA][20:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_op1_sel = _RANDOM[9'hEA][22:21];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_op2_sel = _RANDOM[9'hEA][25:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_imm_sel = _RANDOM[9'hEA][28:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_op_fcn = {_RANDOM[9'hEA][31:29], _RANDOM[9'hEB][0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_fcn_dw = _RANDOM[9'hEB][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_csr_cmd = _RANDOM[9'hEB][4:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_is_load = _RANDOM[9'hEB][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_is_sta = _RANDOM[9'hEB][6];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ctrl_is_std = _RANDOM[9'hEB][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_iw_state = _RANDOM[9'hEB][9:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_iw_p1_poisoned = _RANDOM[9'hEB][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_iw_p2_poisoned = _RANDOM[9'hEB][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_is_sfb = _RANDOM[9'hEB][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_ftq_idx = _RANDOM[9'hEC][8:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_edge_inst = _RANDOM[9'hEC][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_pc_lob = _RANDOM[9'hEC][15:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_taken = _RANDOM[9'hEC][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_csr_addr = _RANDOM[9'hED][16:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_rxq_idx = _RANDOM[9'hEE][3:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_xcpt_pf_if = _RANDOM[9'hF3][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_xcpt_ae_if = _RANDOM[9'hF3][6];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_xcpt_ma_if = _RANDOM[9'hF3][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_bp_debug_if = _RANDOM[9'hF3][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_bp_xcpt_if = _RANDOM[9'hF3][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_debug_fsrc = _RANDOM[9'hF3][11:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_18_debug_tsrc = _RANDOM[9'hF3][13:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_inst = {_RANDOM[9'hF3][31:21], _RANDOM[9'hF4][20:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_19_debug_inst = {_RANDOM[9'hF4][31:21], _RANDOM[9'hF5][20:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_19_is_rvc = _RANDOM[9'hF5][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_debug_pc = {_RANDOM[9'hF5][31:22], _RANDOM[9'hF6][29:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_br_type = _RANDOM[9'hF7][14:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_op1_sel = _RANDOM[9'hF7][16:15];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_op2_sel = _RANDOM[9'hF7][19:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_imm_sel = _RANDOM[9'hF7][22:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_op_fcn = _RANDOM[9'hF7][26:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_fcn_dw = _RANDOM[9'hF7][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_csr_cmd = _RANDOM[9'hF7][30:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_is_load = _RANDOM[9'hF7][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_is_sta = _RANDOM[9'hF8][0];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ctrl_is_std = _RANDOM[9'hF8][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_iw_state = _RANDOM[9'hF8][3:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_iw_p1_poisoned = _RANDOM[9'hF8][4];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_iw_p2_poisoned = _RANDOM[9'hF8][5];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_is_sfb = _RANDOM[9'hF8][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_ftq_idx = {_RANDOM[9'hF8][31:30], _RANDOM[9'hF9][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_19_edge_inst = _RANDOM[9'hF9][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_pc_lob = _RANDOM[9'hF9][9:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_taken = _RANDOM[9'hF9][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_csr_addr = {_RANDOM[9'hF9][31], _RANDOM[9'hFA][10:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_19_rxq_idx = _RANDOM[9'hFA][29:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_xcpt_pf_if = _RANDOM[9'hFF][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_xcpt_ae_if = _RANDOM[9'h100][0];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_xcpt_ma_if = _RANDOM[9'h100][1];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_bp_debug_if = _RANDOM[9'h100][2];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_bp_xcpt_if = _RANDOM[9'h100][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_debug_fsrc = _RANDOM[9'h100][5:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_19_debug_tsrc = _RANDOM[9'h100][7:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_inst = {_RANDOM[9'h100][31:15], _RANDOM[9'h101][14:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_20_debug_inst = {_RANDOM[9'h101][31:15], _RANDOM[9'h102][14:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_20_is_rvc = _RANDOM[9'h102][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_debug_pc = {_RANDOM[9'h102][31:16], _RANDOM[9'h103][23:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_br_type = _RANDOM[9'h104][8:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_op1_sel = _RANDOM[9'h104][10:9];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_op2_sel = _RANDOM[9'h104][13:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_imm_sel = _RANDOM[9'h104][16:14];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_op_fcn = _RANDOM[9'h104][20:17];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_fcn_dw = _RANDOM[9'h104][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_csr_cmd = _RANDOM[9'h104][24:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_is_load = _RANDOM[9'h104][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_is_sta = _RANDOM[9'h104][26];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ctrl_is_std = _RANDOM[9'h104][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_iw_state = _RANDOM[9'h104][29:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_iw_p1_poisoned = _RANDOM[9'h104][30];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_iw_p2_poisoned = _RANDOM[9'h104][31];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_is_sfb = _RANDOM[9'h105][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_ftq_idx = _RANDOM[9'h105][28:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_edge_inst = _RANDOM[9'h105][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_pc_lob = {_RANDOM[9'h105][31:30], _RANDOM[9'h106][3:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_20_taken = _RANDOM[9'h106][4];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_csr_addr = {_RANDOM[9'h106][31:25], _RANDOM[9'h107][4:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_20_rxq_idx = _RANDOM[9'h107][23:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_xcpt_pf_if = _RANDOM[9'h10C][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_xcpt_ae_if = _RANDOM[9'h10C][26];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_xcpt_ma_if = _RANDOM[9'h10C][27];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_bp_debug_if = _RANDOM[9'h10C][28];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_bp_xcpt_if = _RANDOM[9'h10C][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_debug_fsrc = _RANDOM[9'h10C][31:30];	// fetch-buffer.scala:57:16
        fb_uop_ram_20_debug_tsrc = _RANDOM[9'h10D][1:0];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_inst = {_RANDOM[9'h10D][31:9], _RANDOM[9'h10E][8:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_21_debug_inst = {_RANDOM[9'h10E][31:9], _RANDOM[9'h10F][8:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_21_is_rvc = _RANDOM[9'h10F][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_debug_pc = {_RANDOM[9'h10F][31:10], _RANDOM[9'h110][17:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_br_type = {_RANDOM[9'h110][31], _RANDOM[9'h111][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_op1_sel = _RANDOM[9'h111][4:3];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_op2_sel = _RANDOM[9'h111][7:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_imm_sel = _RANDOM[9'h111][10:8];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_op_fcn = _RANDOM[9'h111][14:11];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_fcn_dw = _RANDOM[9'h111][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_csr_cmd = _RANDOM[9'h111][18:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_is_load = _RANDOM[9'h111][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_is_sta = _RANDOM[9'h111][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ctrl_is_std = _RANDOM[9'h111][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_iw_state = _RANDOM[9'h111][23:22];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_iw_p1_poisoned = _RANDOM[9'h111][24];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_iw_p2_poisoned = _RANDOM[9'h111][25];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_is_sfb = _RANDOM[9'h111][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_ftq_idx = _RANDOM[9'h112][22:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_edge_inst = _RANDOM[9'h112][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_pc_lob = _RANDOM[9'h112][29:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_taken = _RANDOM[9'h112][30];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_csr_addr = _RANDOM[9'h113][30:19];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_rxq_idx = _RANDOM[9'h114][17:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_xcpt_pf_if = _RANDOM[9'h119][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_xcpt_ae_if = _RANDOM[9'h119][20];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_xcpt_ma_if = _RANDOM[9'h119][21];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_bp_debug_if = _RANDOM[9'h119][22];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_bp_xcpt_if = _RANDOM[9'h119][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_debug_fsrc = _RANDOM[9'h119][25:24];	// fetch-buffer.scala:57:16
        fb_uop_ram_21_debug_tsrc = _RANDOM[9'h119][27:26];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_inst = {_RANDOM[9'h11A][31:3], _RANDOM[9'h11B][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_22_debug_inst = {_RANDOM[9'h11B][31:3], _RANDOM[9'h11C][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_22_is_rvc = _RANDOM[9'h11C][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_debug_pc = {_RANDOM[9'h11C][31:4], _RANDOM[9'h11D][11:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_br_type = _RANDOM[9'h11D][28:25];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_op1_sel = _RANDOM[9'h11D][30:29];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_op2_sel = {_RANDOM[9'h11D][31], _RANDOM[9'h11E][1:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_imm_sel = _RANDOM[9'h11E][4:2];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_op_fcn = _RANDOM[9'h11E][8:5];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_fcn_dw = _RANDOM[9'h11E][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_csr_cmd = _RANDOM[9'h11E][12:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_is_load = _RANDOM[9'h11E][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_is_sta = _RANDOM[9'h11E][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ctrl_is_std = _RANDOM[9'h11E][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_iw_state = _RANDOM[9'h11E][17:16];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_iw_p1_poisoned = _RANDOM[9'h11E][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_iw_p2_poisoned = _RANDOM[9'h11E][19];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_is_sfb = _RANDOM[9'h11E][23];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_ftq_idx = _RANDOM[9'h11F][16:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_edge_inst = _RANDOM[9'h11F][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_pc_lob = _RANDOM[9'h11F][23:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_taken = _RANDOM[9'h11F][24];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_csr_addr = _RANDOM[9'h120][24:13];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_rxq_idx = _RANDOM[9'h121][11:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_xcpt_pf_if = _RANDOM[9'h126][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_xcpt_ae_if = _RANDOM[9'h126][14];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_xcpt_ma_if = _RANDOM[9'h126][15];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_bp_debug_if = _RANDOM[9'h126][16];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_bp_xcpt_if = _RANDOM[9'h126][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_debug_fsrc = _RANDOM[9'h126][19:18];	// fetch-buffer.scala:57:16
        fb_uop_ram_22_debug_tsrc = _RANDOM[9'h126][21:20];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_inst = {_RANDOM[9'h126][31:29], _RANDOM[9'h127][28:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_23_debug_inst = {_RANDOM[9'h127][31:29], _RANDOM[9'h128][28:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_23_is_rvc = _RANDOM[9'h128][29];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_debug_pc =
          {_RANDOM[9'h128][31:30], _RANDOM[9'h129], _RANDOM[9'h12A][5:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_br_type = _RANDOM[9'h12A][22:19];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_op1_sel = _RANDOM[9'h12A][24:23];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_op2_sel = _RANDOM[9'h12A][27:25];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_imm_sel = _RANDOM[9'h12A][30:28];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_op_fcn = {_RANDOM[9'h12A][31], _RANDOM[9'h12B][2:0]};	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_fcn_dw = _RANDOM[9'h12B][3];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_csr_cmd = _RANDOM[9'h12B][6:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_is_load = _RANDOM[9'h12B][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_is_sta = _RANDOM[9'h12B][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ctrl_is_std = _RANDOM[9'h12B][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_iw_state = _RANDOM[9'h12B][11:10];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_iw_p1_poisoned = _RANDOM[9'h12B][12];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_iw_p2_poisoned = _RANDOM[9'h12B][13];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_is_sfb = _RANDOM[9'h12B][17];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_ftq_idx = _RANDOM[9'h12C][10:6];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_edge_inst = _RANDOM[9'h12C][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_pc_lob = _RANDOM[9'h12C][17:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_taken = _RANDOM[9'h12C][18];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_csr_addr = _RANDOM[9'h12D][18:7];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_rxq_idx = _RANDOM[9'h12E][5:4];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_xcpt_pf_if = _RANDOM[9'h133][7];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_xcpt_ae_if = _RANDOM[9'h133][8];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_xcpt_ma_if = _RANDOM[9'h133][9];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_bp_debug_if = _RANDOM[9'h133][10];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_bp_xcpt_if = _RANDOM[9'h133][11];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_debug_fsrc = _RANDOM[9'h133][13:12];	// fetch-buffer.scala:57:16
        fb_uop_ram_23_debug_tsrc = _RANDOM[9'h133][15:14];	// fetch-buffer.scala:57:16
        head = _RANDOM[9'h133][23:16];	// fetch-buffer.scala:57:16, :61:21
        tail = {_RANDOM[9'h133][31:24], _RANDOM[9'h134][15:0]};	// fetch-buffer.scala:57:16, :62:21
        maybe_full = _RANDOM[9'h134][16];	// fetch-buffer.scala:62:21, :64:27
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign io_enq_ready = ~_do_enq_T_1;	// fetch-buffer.scala:82:{16,40}
  assign io_deq_valid = _deq_valids_T_7 != 3'h7;	// fetch-buffer.scala:170:38, frontend.scala:161:39, util.scala:384:54
  assign io_deq_bits_uops_0_valid = ~reset & _deq_valids_T_8[0];	// fetch-buffer.scala:161:{21,53}, :168:72, :195:23, :196:41
  assign io_deq_bits_uops_0_bits_inst =
    (head[0] ? fb_uop_ram_0_inst : 32'h0) | (head[1] ? fb_uop_ram_3_inst : 32'h0)
    | (head[2] ? fb_uop_ram_6_inst : 32'h0) | (head[3] ? fb_uop_ram_9_inst : 32'h0)
    | (head[4] ? fb_uop_ram_12_inst : 32'h0) | (head[5] ? fb_uop_ram_15_inst : 32'h0)
    | (head[6] ? fb_uop_ram_18_inst : 32'h0) | (head[7] ? fb_uop_ram_21_inst : 32'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_debug_inst =
    (head[0] ? fb_uop_ram_0_debug_inst : 32'h0)
    | (head[1] ? fb_uop_ram_3_debug_inst : 32'h0)
    | (head[2] ? fb_uop_ram_6_debug_inst : 32'h0)
    | (head[3] ? fb_uop_ram_9_debug_inst : 32'h0)
    | (head[4] ? fb_uop_ram_12_debug_inst : 32'h0)
    | (head[5] ? fb_uop_ram_15_debug_inst : 32'h0)
    | (head[6] ? fb_uop_ram_18_debug_inst : 32'h0)
    | (head[7] ? fb_uop_ram_21_debug_inst : 32'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_is_rvc =
    head[0] & fb_uop_ram_0_is_rvc | head[1] & fb_uop_ram_3_is_rvc | head[2]
    & fb_uop_ram_6_is_rvc | head[3] & fb_uop_ram_9_is_rvc | head[4] & fb_uop_ram_12_is_rvc
    | head[5] & fb_uop_ram_15_is_rvc | head[6] & fb_uop_ram_18_is_rvc | head[7]
    & fb_uop_ram_21_is_rvc;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_debug_pc =
    (head[0] ? fb_uop_ram_0_debug_pc : 40'h0) | (head[1] ? fb_uop_ram_3_debug_pc : 40'h0)
    | (head[2] ? fb_uop_ram_6_debug_pc : 40'h0)
    | (head[3] ? fb_uop_ram_9_debug_pc : 40'h0)
    | (head[4] ? fb_uop_ram_12_debug_pc : 40'h0)
    | (head[5] ? fb_uop_ram_15_debug_pc : 40'h0)
    | (head[6] ? fb_uop_ram_18_debug_pc : 40'h0)
    | (head[7] ? fb_uop_ram_21_debug_pc : 40'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_br_type =
    (head[0] ? fb_uop_ram_0_ctrl_br_type : 4'h0)
    | (head[1] ? fb_uop_ram_3_ctrl_br_type : 4'h0)
    | (head[2] ? fb_uop_ram_6_ctrl_br_type : 4'h0)
    | (head[3] ? fb_uop_ram_9_ctrl_br_type : 4'h0)
    | (head[4] ? fb_uop_ram_12_ctrl_br_type : 4'h0)
    | (head[5] ? fb_uop_ram_15_ctrl_br_type : 4'h0)
    | (head[6] ? fb_uop_ram_18_ctrl_br_type : 4'h0)
    | (head[7] ? fb_uop_ram_21_ctrl_br_type : 4'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_op1_sel =
    (head[0] ? fb_uop_ram_0_ctrl_op1_sel : 2'h0)
    | (head[1] ? fb_uop_ram_3_ctrl_op1_sel : 2'h0)
    | (head[2] ? fb_uop_ram_6_ctrl_op1_sel : 2'h0)
    | (head[3] ? fb_uop_ram_9_ctrl_op1_sel : 2'h0)
    | (head[4] ? fb_uop_ram_12_ctrl_op1_sel : 2'h0)
    | (head[5] ? fb_uop_ram_15_ctrl_op1_sel : 2'h0)
    | (head[6] ? fb_uop_ram_18_ctrl_op1_sel : 2'h0)
    | (head[7] ? fb_uop_ram_21_ctrl_op1_sel : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_op2_sel =
    (head[0] ? fb_uop_ram_0_ctrl_op2_sel : 3'h0)
    | (head[1] ? fb_uop_ram_3_ctrl_op2_sel : 3'h0)
    | (head[2] ? fb_uop_ram_6_ctrl_op2_sel : 3'h0)
    | (head[3] ? fb_uop_ram_9_ctrl_op2_sel : 3'h0)
    | (head[4] ? fb_uop_ram_12_ctrl_op2_sel : 3'h0)
    | (head[5] ? fb_uop_ram_15_ctrl_op2_sel : 3'h0)
    | (head[6] ? fb_uop_ram_18_ctrl_op2_sel : 3'h0)
    | (head[7] ? fb_uop_ram_21_ctrl_op2_sel : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_imm_sel =
    (head[0] ? fb_uop_ram_0_ctrl_imm_sel : 3'h0)
    | (head[1] ? fb_uop_ram_3_ctrl_imm_sel : 3'h0)
    | (head[2] ? fb_uop_ram_6_ctrl_imm_sel : 3'h0)
    | (head[3] ? fb_uop_ram_9_ctrl_imm_sel : 3'h0)
    | (head[4] ? fb_uop_ram_12_ctrl_imm_sel : 3'h0)
    | (head[5] ? fb_uop_ram_15_ctrl_imm_sel : 3'h0)
    | (head[6] ? fb_uop_ram_18_ctrl_imm_sel : 3'h0)
    | (head[7] ? fb_uop_ram_21_ctrl_imm_sel : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_op_fcn =
    (head[0] ? fb_uop_ram_0_ctrl_op_fcn : 4'h0)
    | (head[1] ? fb_uop_ram_3_ctrl_op_fcn : 4'h0)
    | (head[2] ? fb_uop_ram_6_ctrl_op_fcn : 4'h0)
    | (head[3] ? fb_uop_ram_9_ctrl_op_fcn : 4'h0)
    | (head[4] ? fb_uop_ram_12_ctrl_op_fcn : 4'h0)
    | (head[5] ? fb_uop_ram_15_ctrl_op_fcn : 4'h0)
    | (head[6] ? fb_uop_ram_18_ctrl_op_fcn : 4'h0)
    | (head[7] ? fb_uop_ram_21_ctrl_op_fcn : 4'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_fcn_dw =
    head[0] & fb_uop_ram_0_ctrl_fcn_dw | head[1] & fb_uop_ram_3_ctrl_fcn_dw | head[2]
    & fb_uop_ram_6_ctrl_fcn_dw | head[3] & fb_uop_ram_9_ctrl_fcn_dw | head[4]
    & fb_uop_ram_12_ctrl_fcn_dw | head[5] & fb_uop_ram_15_ctrl_fcn_dw | head[6]
    & fb_uop_ram_18_ctrl_fcn_dw | head[7] & fb_uop_ram_21_ctrl_fcn_dw;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_csr_cmd =
    (head[0] ? fb_uop_ram_0_ctrl_csr_cmd : 3'h0)
    | (head[1] ? fb_uop_ram_3_ctrl_csr_cmd : 3'h0)
    | (head[2] ? fb_uop_ram_6_ctrl_csr_cmd : 3'h0)
    | (head[3] ? fb_uop_ram_9_ctrl_csr_cmd : 3'h0)
    | (head[4] ? fb_uop_ram_12_ctrl_csr_cmd : 3'h0)
    | (head[5] ? fb_uop_ram_15_ctrl_csr_cmd : 3'h0)
    | (head[6] ? fb_uop_ram_18_ctrl_csr_cmd : 3'h0)
    | (head[7] ? fb_uop_ram_21_ctrl_csr_cmd : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_is_load =
    head[0] & fb_uop_ram_0_ctrl_is_load | head[1] & fb_uop_ram_3_ctrl_is_load | head[2]
    & fb_uop_ram_6_ctrl_is_load | head[3] & fb_uop_ram_9_ctrl_is_load | head[4]
    & fb_uop_ram_12_ctrl_is_load | head[5] & fb_uop_ram_15_ctrl_is_load | head[6]
    & fb_uop_ram_18_ctrl_is_load | head[7] & fb_uop_ram_21_ctrl_is_load;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_is_sta =
    head[0] & fb_uop_ram_0_ctrl_is_sta | head[1] & fb_uop_ram_3_ctrl_is_sta | head[2]
    & fb_uop_ram_6_ctrl_is_sta | head[3] & fb_uop_ram_9_ctrl_is_sta | head[4]
    & fb_uop_ram_12_ctrl_is_sta | head[5] & fb_uop_ram_15_ctrl_is_sta | head[6]
    & fb_uop_ram_18_ctrl_is_sta | head[7] & fb_uop_ram_21_ctrl_is_sta;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_ctrl_is_std =
    head[0] & fb_uop_ram_0_ctrl_is_std | head[1] & fb_uop_ram_3_ctrl_is_std | head[2]
    & fb_uop_ram_6_ctrl_is_std | head[3] & fb_uop_ram_9_ctrl_is_std | head[4]
    & fb_uop_ram_12_ctrl_is_std | head[5] & fb_uop_ram_15_ctrl_is_std | head[6]
    & fb_uop_ram_18_ctrl_is_std | head[7] & fb_uop_ram_21_ctrl_is_std;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_iw_state =
    (head[0] ? fb_uop_ram_0_iw_state : 2'h0) | (head[1] ? fb_uop_ram_3_iw_state : 2'h0)
    | (head[2] ? fb_uop_ram_6_iw_state : 2'h0) | (head[3] ? fb_uop_ram_9_iw_state : 2'h0)
    | (head[4] ? fb_uop_ram_12_iw_state : 2'h0)
    | (head[5] ? fb_uop_ram_15_iw_state : 2'h0)
    | (head[6] ? fb_uop_ram_18_iw_state : 2'h0)
    | (head[7] ? fb_uop_ram_21_iw_state : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_iw_p1_poisoned =
    head[0] & fb_uop_ram_0_iw_p1_poisoned | head[1] & fb_uop_ram_3_iw_p1_poisoned
    | head[2] & fb_uop_ram_6_iw_p1_poisoned | head[3] & fb_uop_ram_9_iw_p1_poisoned
    | head[4] & fb_uop_ram_12_iw_p1_poisoned | head[5] & fb_uop_ram_15_iw_p1_poisoned
    | head[6] & fb_uop_ram_18_iw_p1_poisoned | head[7] & fb_uop_ram_21_iw_p1_poisoned;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_iw_p2_poisoned =
    head[0] & fb_uop_ram_0_iw_p2_poisoned | head[1] & fb_uop_ram_3_iw_p2_poisoned
    | head[2] & fb_uop_ram_6_iw_p2_poisoned | head[3] & fb_uop_ram_9_iw_p2_poisoned
    | head[4] & fb_uop_ram_12_iw_p2_poisoned | head[5] & fb_uop_ram_15_iw_p2_poisoned
    | head[6] & fb_uop_ram_18_iw_p2_poisoned | head[7] & fb_uop_ram_21_iw_p2_poisoned;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_is_sfb =
    head[0] & fb_uop_ram_0_is_sfb | head[1] & fb_uop_ram_3_is_sfb | head[2]
    & fb_uop_ram_6_is_sfb | head[3] & fb_uop_ram_9_is_sfb | head[4] & fb_uop_ram_12_is_sfb
    | head[5] & fb_uop_ram_15_is_sfb | head[6] & fb_uop_ram_18_is_sfb | head[7]
    & fb_uop_ram_21_is_sfb;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_ftq_idx =
    (head[0] ? fb_uop_ram_0_ftq_idx : 5'h0) | (head[1] ? fb_uop_ram_3_ftq_idx : 5'h0)
    | (head[2] ? fb_uop_ram_6_ftq_idx : 5'h0) | (head[3] ? fb_uop_ram_9_ftq_idx : 5'h0)
    | (head[4] ? fb_uop_ram_12_ftq_idx : 5'h0) | (head[5] ? fb_uop_ram_15_ftq_idx : 5'h0)
    | (head[6] ? fb_uop_ram_18_ftq_idx : 5'h0) | (head[7] ? fb_uop_ram_21_ftq_idx : 5'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_edge_inst =
    head[0] & fb_uop_ram_0_edge_inst | head[1] & fb_uop_ram_3_edge_inst | head[2]
    & fb_uop_ram_6_edge_inst | head[3] & fb_uop_ram_9_edge_inst | head[4]
    & fb_uop_ram_12_edge_inst | head[5] & fb_uop_ram_15_edge_inst | head[6]
    & fb_uop_ram_18_edge_inst | head[7] & fb_uop_ram_21_edge_inst;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_pc_lob =
    (head[0] ? fb_uop_ram_0_pc_lob : 6'h0) | (head[1] ? fb_uop_ram_3_pc_lob : 6'h0)
    | (head[2] ? fb_uop_ram_6_pc_lob : 6'h0) | (head[3] ? fb_uop_ram_9_pc_lob : 6'h0)
    | (head[4] ? fb_uop_ram_12_pc_lob : 6'h0) | (head[5] ? fb_uop_ram_15_pc_lob : 6'h0)
    | (head[6] ? fb_uop_ram_18_pc_lob : 6'h0) | (head[7] ? fb_uop_ram_21_pc_lob : 6'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_taken =
    head[0] & fb_uop_ram_0_taken | head[1] & fb_uop_ram_3_taken | head[2]
    & fb_uop_ram_6_taken | head[3] & fb_uop_ram_9_taken | head[4] & fb_uop_ram_12_taken
    | head[5] & fb_uop_ram_15_taken | head[6] & fb_uop_ram_18_taken | head[7]
    & fb_uop_ram_21_taken;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_csr_addr =
    (head[0] ? fb_uop_ram_0_csr_addr : 12'h0) | (head[1] ? fb_uop_ram_3_csr_addr : 12'h0)
    | (head[2] ? fb_uop_ram_6_csr_addr : 12'h0)
    | (head[3] ? fb_uop_ram_9_csr_addr : 12'h0)
    | (head[4] ? fb_uop_ram_12_csr_addr : 12'h0)
    | (head[5] ? fb_uop_ram_15_csr_addr : 12'h0)
    | (head[6] ? fb_uop_ram_18_csr_addr : 12'h0)
    | (head[7] ? fb_uop_ram_21_csr_addr : 12'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_rxq_idx =
    (head[0] ? fb_uop_ram_0_rxq_idx : 2'h0) | (head[1] ? fb_uop_ram_3_rxq_idx : 2'h0)
    | (head[2] ? fb_uop_ram_6_rxq_idx : 2'h0) | (head[3] ? fb_uop_ram_9_rxq_idx : 2'h0)
    | (head[4] ? fb_uop_ram_12_rxq_idx : 2'h0) | (head[5] ? fb_uop_ram_15_rxq_idx : 2'h0)
    | (head[6] ? fb_uop_ram_18_rxq_idx : 2'h0) | (head[7] ? fb_uop_ram_21_rxq_idx : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_xcpt_pf_if =
    head[0] & fb_uop_ram_0_xcpt_pf_if | head[1] & fb_uop_ram_3_xcpt_pf_if | head[2]
    & fb_uop_ram_6_xcpt_pf_if | head[3] & fb_uop_ram_9_xcpt_pf_if | head[4]
    & fb_uop_ram_12_xcpt_pf_if | head[5] & fb_uop_ram_15_xcpt_pf_if | head[6]
    & fb_uop_ram_18_xcpt_pf_if | head[7] & fb_uop_ram_21_xcpt_pf_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_xcpt_ae_if =
    head[0] & fb_uop_ram_0_xcpt_ae_if | head[1] & fb_uop_ram_3_xcpt_ae_if | head[2]
    & fb_uop_ram_6_xcpt_ae_if | head[3] & fb_uop_ram_9_xcpt_ae_if | head[4]
    & fb_uop_ram_12_xcpt_ae_if | head[5] & fb_uop_ram_15_xcpt_ae_if | head[6]
    & fb_uop_ram_18_xcpt_ae_if | head[7] & fb_uop_ram_21_xcpt_ae_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_xcpt_ma_if =
    head[0] & fb_uop_ram_0_xcpt_ma_if | head[1] & fb_uop_ram_3_xcpt_ma_if | head[2]
    & fb_uop_ram_6_xcpt_ma_if | head[3] & fb_uop_ram_9_xcpt_ma_if | head[4]
    & fb_uop_ram_12_xcpt_ma_if | head[5] & fb_uop_ram_15_xcpt_ma_if | head[6]
    & fb_uop_ram_18_xcpt_ma_if | head[7] & fb_uop_ram_21_xcpt_ma_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_bp_debug_if =
    head[0] & fb_uop_ram_0_bp_debug_if | head[1] & fb_uop_ram_3_bp_debug_if | head[2]
    & fb_uop_ram_6_bp_debug_if | head[3] & fb_uop_ram_9_bp_debug_if | head[4]
    & fb_uop_ram_12_bp_debug_if | head[5] & fb_uop_ram_15_bp_debug_if | head[6]
    & fb_uop_ram_18_bp_debug_if | head[7] & fb_uop_ram_21_bp_debug_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_bp_xcpt_if =
    head[0] & fb_uop_ram_0_bp_xcpt_if | head[1] & fb_uop_ram_3_bp_xcpt_if | head[2]
    & fb_uop_ram_6_bp_xcpt_if | head[3] & fb_uop_ram_9_bp_xcpt_if | head[4]
    & fb_uop_ram_12_bp_xcpt_if | head[5] & fb_uop_ram_15_bp_xcpt_if | head[6]
    & fb_uop_ram_18_bp_xcpt_if | head[7] & fb_uop_ram_21_bp_xcpt_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_0_bits_debug_fsrc =
    (head[0] ? fb_uop_ram_0_debug_fsrc : 2'h0)
    | (head[1] ? fb_uop_ram_3_debug_fsrc : 2'h0)
    | (head[2] ? fb_uop_ram_6_debug_fsrc : 2'h0)
    | (head[3] ? fb_uop_ram_9_debug_fsrc : 2'h0)
    | (head[4] ? fb_uop_ram_12_debug_fsrc : 2'h0)
    | (head[5] ? fb_uop_ram_15_debug_fsrc : 2'h0)
    | (head[6] ? fb_uop_ram_18_debug_fsrc : 2'h0)
    | (head[7] ? fb_uop_ram_21_debug_fsrc : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_0_bits_debug_tsrc =
    (head[0] ? fb_uop_ram_0_debug_tsrc : 2'h0)
    | (head[1] ? fb_uop_ram_3_debug_tsrc : 2'h0)
    | (head[2] ? fb_uop_ram_6_debug_tsrc : 2'h0)
    | (head[3] ? fb_uop_ram_9_debug_tsrc : 2'h0)
    | (head[4] ? fb_uop_ram_12_debug_tsrc : 2'h0)
    | (head[5] ? fb_uop_ram_15_debug_tsrc : 2'h0)
    | (head[6] ? fb_uop_ram_18_debug_tsrc : 2'h0)
    | (head[7] ? fb_uop_ram_21_debug_tsrc : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_valid = ~reset & _deq_valids_T_8[1];	// fetch-buffer.scala:161:{21,53}, :168:72, :195:23, :196:41
  assign io_deq_bits_uops_1_bits_inst =
    (head[0] ? fb_uop_ram_1_inst : 32'h0) | (head[1] ? fb_uop_ram_4_inst : 32'h0)
    | (head[2] ? fb_uop_ram_7_inst : 32'h0) | (head[3] ? fb_uop_ram_10_inst : 32'h0)
    | (head[4] ? fb_uop_ram_13_inst : 32'h0) | (head[5] ? fb_uop_ram_16_inst : 32'h0)
    | (head[6] ? fb_uop_ram_19_inst : 32'h0) | (head[7] ? fb_uop_ram_22_inst : 32'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_debug_inst =
    (head[0] ? fb_uop_ram_1_debug_inst : 32'h0)
    | (head[1] ? fb_uop_ram_4_debug_inst : 32'h0)
    | (head[2] ? fb_uop_ram_7_debug_inst : 32'h0)
    | (head[3] ? fb_uop_ram_10_debug_inst : 32'h0)
    | (head[4] ? fb_uop_ram_13_debug_inst : 32'h0)
    | (head[5] ? fb_uop_ram_16_debug_inst : 32'h0)
    | (head[6] ? fb_uop_ram_19_debug_inst : 32'h0)
    | (head[7] ? fb_uop_ram_22_debug_inst : 32'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_is_rvc =
    head[0] & fb_uop_ram_1_is_rvc | head[1] & fb_uop_ram_4_is_rvc | head[2]
    & fb_uop_ram_7_is_rvc | head[3] & fb_uop_ram_10_is_rvc | head[4]
    & fb_uop_ram_13_is_rvc | head[5] & fb_uop_ram_16_is_rvc | head[6]
    & fb_uop_ram_19_is_rvc | head[7] & fb_uop_ram_22_is_rvc;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_debug_pc =
    (head[0] ? fb_uop_ram_1_debug_pc : 40'h0) | (head[1] ? fb_uop_ram_4_debug_pc : 40'h0)
    | (head[2] ? fb_uop_ram_7_debug_pc : 40'h0)
    | (head[3] ? fb_uop_ram_10_debug_pc : 40'h0)
    | (head[4] ? fb_uop_ram_13_debug_pc : 40'h0)
    | (head[5] ? fb_uop_ram_16_debug_pc : 40'h0)
    | (head[6] ? fb_uop_ram_19_debug_pc : 40'h0)
    | (head[7] ? fb_uop_ram_22_debug_pc : 40'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_br_type =
    (head[0] ? fb_uop_ram_1_ctrl_br_type : 4'h0)
    | (head[1] ? fb_uop_ram_4_ctrl_br_type : 4'h0)
    | (head[2] ? fb_uop_ram_7_ctrl_br_type : 4'h0)
    | (head[3] ? fb_uop_ram_10_ctrl_br_type : 4'h0)
    | (head[4] ? fb_uop_ram_13_ctrl_br_type : 4'h0)
    | (head[5] ? fb_uop_ram_16_ctrl_br_type : 4'h0)
    | (head[6] ? fb_uop_ram_19_ctrl_br_type : 4'h0)
    | (head[7] ? fb_uop_ram_22_ctrl_br_type : 4'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_op1_sel =
    (head[0] ? fb_uop_ram_1_ctrl_op1_sel : 2'h0)
    | (head[1] ? fb_uop_ram_4_ctrl_op1_sel : 2'h0)
    | (head[2] ? fb_uop_ram_7_ctrl_op1_sel : 2'h0)
    | (head[3] ? fb_uop_ram_10_ctrl_op1_sel : 2'h0)
    | (head[4] ? fb_uop_ram_13_ctrl_op1_sel : 2'h0)
    | (head[5] ? fb_uop_ram_16_ctrl_op1_sel : 2'h0)
    | (head[6] ? fb_uop_ram_19_ctrl_op1_sel : 2'h0)
    | (head[7] ? fb_uop_ram_22_ctrl_op1_sel : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_op2_sel =
    (head[0] ? fb_uop_ram_1_ctrl_op2_sel : 3'h0)
    | (head[1] ? fb_uop_ram_4_ctrl_op2_sel : 3'h0)
    | (head[2] ? fb_uop_ram_7_ctrl_op2_sel : 3'h0)
    | (head[3] ? fb_uop_ram_10_ctrl_op2_sel : 3'h0)
    | (head[4] ? fb_uop_ram_13_ctrl_op2_sel : 3'h0)
    | (head[5] ? fb_uop_ram_16_ctrl_op2_sel : 3'h0)
    | (head[6] ? fb_uop_ram_19_ctrl_op2_sel : 3'h0)
    | (head[7] ? fb_uop_ram_22_ctrl_op2_sel : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_imm_sel =
    (head[0] ? fb_uop_ram_1_ctrl_imm_sel : 3'h0)
    | (head[1] ? fb_uop_ram_4_ctrl_imm_sel : 3'h0)
    | (head[2] ? fb_uop_ram_7_ctrl_imm_sel : 3'h0)
    | (head[3] ? fb_uop_ram_10_ctrl_imm_sel : 3'h0)
    | (head[4] ? fb_uop_ram_13_ctrl_imm_sel : 3'h0)
    | (head[5] ? fb_uop_ram_16_ctrl_imm_sel : 3'h0)
    | (head[6] ? fb_uop_ram_19_ctrl_imm_sel : 3'h0)
    | (head[7] ? fb_uop_ram_22_ctrl_imm_sel : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_op_fcn =
    (head[0] ? fb_uop_ram_1_ctrl_op_fcn : 4'h0)
    | (head[1] ? fb_uop_ram_4_ctrl_op_fcn : 4'h0)
    | (head[2] ? fb_uop_ram_7_ctrl_op_fcn : 4'h0)
    | (head[3] ? fb_uop_ram_10_ctrl_op_fcn : 4'h0)
    | (head[4] ? fb_uop_ram_13_ctrl_op_fcn : 4'h0)
    | (head[5] ? fb_uop_ram_16_ctrl_op_fcn : 4'h0)
    | (head[6] ? fb_uop_ram_19_ctrl_op_fcn : 4'h0)
    | (head[7] ? fb_uop_ram_22_ctrl_op_fcn : 4'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_fcn_dw =
    head[0] & fb_uop_ram_1_ctrl_fcn_dw | head[1] & fb_uop_ram_4_ctrl_fcn_dw | head[2]
    & fb_uop_ram_7_ctrl_fcn_dw | head[3] & fb_uop_ram_10_ctrl_fcn_dw | head[4]
    & fb_uop_ram_13_ctrl_fcn_dw | head[5] & fb_uop_ram_16_ctrl_fcn_dw | head[6]
    & fb_uop_ram_19_ctrl_fcn_dw | head[7] & fb_uop_ram_22_ctrl_fcn_dw;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_csr_cmd =
    (head[0] ? fb_uop_ram_1_ctrl_csr_cmd : 3'h0)
    | (head[1] ? fb_uop_ram_4_ctrl_csr_cmd : 3'h0)
    | (head[2] ? fb_uop_ram_7_ctrl_csr_cmd : 3'h0)
    | (head[3] ? fb_uop_ram_10_ctrl_csr_cmd : 3'h0)
    | (head[4] ? fb_uop_ram_13_ctrl_csr_cmd : 3'h0)
    | (head[5] ? fb_uop_ram_16_ctrl_csr_cmd : 3'h0)
    | (head[6] ? fb_uop_ram_19_ctrl_csr_cmd : 3'h0)
    | (head[7] ? fb_uop_ram_22_ctrl_csr_cmd : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_is_load =
    head[0] & fb_uop_ram_1_ctrl_is_load | head[1] & fb_uop_ram_4_ctrl_is_load | head[2]
    & fb_uop_ram_7_ctrl_is_load | head[3] & fb_uop_ram_10_ctrl_is_load | head[4]
    & fb_uop_ram_13_ctrl_is_load | head[5] & fb_uop_ram_16_ctrl_is_load | head[6]
    & fb_uop_ram_19_ctrl_is_load | head[7] & fb_uop_ram_22_ctrl_is_load;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_is_sta =
    head[0] & fb_uop_ram_1_ctrl_is_sta | head[1] & fb_uop_ram_4_ctrl_is_sta | head[2]
    & fb_uop_ram_7_ctrl_is_sta | head[3] & fb_uop_ram_10_ctrl_is_sta | head[4]
    & fb_uop_ram_13_ctrl_is_sta | head[5] & fb_uop_ram_16_ctrl_is_sta | head[6]
    & fb_uop_ram_19_ctrl_is_sta | head[7] & fb_uop_ram_22_ctrl_is_sta;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_ctrl_is_std =
    head[0] & fb_uop_ram_1_ctrl_is_std | head[1] & fb_uop_ram_4_ctrl_is_std | head[2]
    & fb_uop_ram_7_ctrl_is_std | head[3] & fb_uop_ram_10_ctrl_is_std | head[4]
    & fb_uop_ram_13_ctrl_is_std | head[5] & fb_uop_ram_16_ctrl_is_std | head[6]
    & fb_uop_ram_19_ctrl_is_std | head[7] & fb_uop_ram_22_ctrl_is_std;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_iw_state =
    (head[0] ? fb_uop_ram_1_iw_state : 2'h0) | (head[1] ? fb_uop_ram_4_iw_state : 2'h0)
    | (head[2] ? fb_uop_ram_7_iw_state : 2'h0) | (head[3] ? fb_uop_ram_10_iw_state : 2'h0)
    | (head[4] ? fb_uop_ram_13_iw_state : 2'h0)
    | (head[5] ? fb_uop_ram_16_iw_state : 2'h0)
    | (head[6] ? fb_uop_ram_19_iw_state : 2'h0)
    | (head[7] ? fb_uop_ram_22_iw_state : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_iw_p1_poisoned =
    head[0] & fb_uop_ram_1_iw_p1_poisoned | head[1] & fb_uop_ram_4_iw_p1_poisoned
    | head[2] & fb_uop_ram_7_iw_p1_poisoned | head[3] & fb_uop_ram_10_iw_p1_poisoned
    | head[4] & fb_uop_ram_13_iw_p1_poisoned | head[5] & fb_uop_ram_16_iw_p1_poisoned
    | head[6] & fb_uop_ram_19_iw_p1_poisoned | head[7] & fb_uop_ram_22_iw_p1_poisoned;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_iw_p2_poisoned =
    head[0] & fb_uop_ram_1_iw_p2_poisoned | head[1] & fb_uop_ram_4_iw_p2_poisoned
    | head[2] & fb_uop_ram_7_iw_p2_poisoned | head[3] & fb_uop_ram_10_iw_p2_poisoned
    | head[4] & fb_uop_ram_13_iw_p2_poisoned | head[5] & fb_uop_ram_16_iw_p2_poisoned
    | head[6] & fb_uop_ram_19_iw_p2_poisoned | head[7] & fb_uop_ram_22_iw_p2_poisoned;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_is_sfb =
    head[0] & fb_uop_ram_1_is_sfb | head[1] & fb_uop_ram_4_is_sfb | head[2]
    & fb_uop_ram_7_is_sfb | head[3] & fb_uop_ram_10_is_sfb | head[4]
    & fb_uop_ram_13_is_sfb | head[5] & fb_uop_ram_16_is_sfb | head[6]
    & fb_uop_ram_19_is_sfb | head[7] & fb_uop_ram_22_is_sfb;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_ftq_idx =
    (head[0] ? fb_uop_ram_1_ftq_idx : 5'h0) | (head[1] ? fb_uop_ram_4_ftq_idx : 5'h0)
    | (head[2] ? fb_uop_ram_7_ftq_idx : 5'h0) | (head[3] ? fb_uop_ram_10_ftq_idx : 5'h0)
    | (head[4] ? fb_uop_ram_13_ftq_idx : 5'h0) | (head[5] ? fb_uop_ram_16_ftq_idx : 5'h0)
    | (head[6] ? fb_uop_ram_19_ftq_idx : 5'h0) | (head[7] ? fb_uop_ram_22_ftq_idx : 5'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_edge_inst =
    head[0] & fb_uop_ram_1_edge_inst | head[1] & fb_uop_ram_4_edge_inst | head[2]
    & fb_uop_ram_7_edge_inst | head[3] & fb_uop_ram_10_edge_inst | head[4]
    & fb_uop_ram_13_edge_inst | head[5] & fb_uop_ram_16_edge_inst | head[6]
    & fb_uop_ram_19_edge_inst | head[7] & fb_uop_ram_22_edge_inst;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_pc_lob =
    (head[0] ? fb_uop_ram_1_pc_lob : 6'h0) | (head[1] ? fb_uop_ram_4_pc_lob : 6'h0)
    | (head[2] ? fb_uop_ram_7_pc_lob : 6'h0) | (head[3] ? fb_uop_ram_10_pc_lob : 6'h0)
    | (head[4] ? fb_uop_ram_13_pc_lob : 6'h0) | (head[5] ? fb_uop_ram_16_pc_lob : 6'h0)
    | (head[6] ? fb_uop_ram_19_pc_lob : 6'h0) | (head[7] ? fb_uop_ram_22_pc_lob : 6'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_taken =
    head[0] & fb_uop_ram_1_taken | head[1] & fb_uop_ram_4_taken | head[2]
    & fb_uop_ram_7_taken | head[3] & fb_uop_ram_10_taken | head[4] & fb_uop_ram_13_taken
    | head[5] & fb_uop_ram_16_taken | head[6] & fb_uop_ram_19_taken | head[7]
    & fb_uop_ram_22_taken;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_csr_addr =
    (head[0] ? fb_uop_ram_1_csr_addr : 12'h0) | (head[1] ? fb_uop_ram_4_csr_addr : 12'h0)
    | (head[2] ? fb_uop_ram_7_csr_addr : 12'h0)
    | (head[3] ? fb_uop_ram_10_csr_addr : 12'h0)
    | (head[4] ? fb_uop_ram_13_csr_addr : 12'h0)
    | (head[5] ? fb_uop_ram_16_csr_addr : 12'h0)
    | (head[6] ? fb_uop_ram_19_csr_addr : 12'h0)
    | (head[7] ? fb_uop_ram_22_csr_addr : 12'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_rxq_idx =
    (head[0] ? fb_uop_ram_1_rxq_idx : 2'h0) | (head[1] ? fb_uop_ram_4_rxq_idx : 2'h0)
    | (head[2] ? fb_uop_ram_7_rxq_idx : 2'h0) | (head[3] ? fb_uop_ram_10_rxq_idx : 2'h0)
    | (head[4] ? fb_uop_ram_13_rxq_idx : 2'h0) | (head[5] ? fb_uop_ram_16_rxq_idx : 2'h0)
    | (head[6] ? fb_uop_ram_19_rxq_idx : 2'h0) | (head[7] ? fb_uop_ram_22_rxq_idx : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_xcpt_pf_if =
    head[0] & fb_uop_ram_1_xcpt_pf_if | head[1] & fb_uop_ram_4_xcpt_pf_if | head[2]
    & fb_uop_ram_7_xcpt_pf_if | head[3] & fb_uop_ram_10_xcpt_pf_if | head[4]
    & fb_uop_ram_13_xcpt_pf_if | head[5] & fb_uop_ram_16_xcpt_pf_if | head[6]
    & fb_uop_ram_19_xcpt_pf_if | head[7] & fb_uop_ram_22_xcpt_pf_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_xcpt_ae_if =
    head[0] & fb_uop_ram_1_xcpt_ae_if | head[1] & fb_uop_ram_4_xcpt_ae_if | head[2]
    & fb_uop_ram_7_xcpt_ae_if | head[3] & fb_uop_ram_10_xcpt_ae_if | head[4]
    & fb_uop_ram_13_xcpt_ae_if | head[5] & fb_uop_ram_16_xcpt_ae_if | head[6]
    & fb_uop_ram_19_xcpt_ae_if | head[7] & fb_uop_ram_22_xcpt_ae_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_xcpt_ma_if =
    head[0] & fb_uop_ram_1_xcpt_ma_if | head[1] & fb_uop_ram_4_xcpt_ma_if | head[2]
    & fb_uop_ram_7_xcpt_ma_if | head[3] & fb_uop_ram_10_xcpt_ma_if | head[4]
    & fb_uop_ram_13_xcpt_ma_if | head[5] & fb_uop_ram_16_xcpt_ma_if | head[6]
    & fb_uop_ram_19_xcpt_ma_if | head[7] & fb_uop_ram_22_xcpt_ma_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_bp_debug_if =
    head[0] & fb_uop_ram_1_bp_debug_if | head[1] & fb_uop_ram_4_bp_debug_if | head[2]
    & fb_uop_ram_7_bp_debug_if | head[3] & fb_uop_ram_10_bp_debug_if | head[4]
    & fb_uop_ram_13_bp_debug_if | head[5] & fb_uop_ram_16_bp_debug_if | head[6]
    & fb_uop_ram_19_bp_debug_if | head[7] & fb_uop_ram_22_bp_debug_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_bp_xcpt_if =
    head[0] & fb_uop_ram_1_bp_xcpt_if | head[1] & fb_uop_ram_4_bp_xcpt_if | head[2]
    & fb_uop_ram_7_bp_xcpt_if | head[3] & fb_uop_ram_10_bp_xcpt_if | head[4]
    & fb_uop_ram_13_bp_xcpt_if | head[5] & fb_uop_ram_16_bp_xcpt_if | head[6]
    & fb_uop_ram_19_bp_xcpt_if | head[7] & fb_uop_ram_22_bp_xcpt_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_1_bits_debug_fsrc =
    (head[0] ? fb_uop_ram_1_debug_fsrc : 2'h0)
    | (head[1] ? fb_uop_ram_4_debug_fsrc : 2'h0)
    | (head[2] ? fb_uop_ram_7_debug_fsrc : 2'h0)
    | (head[3] ? fb_uop_ram_10_debug_fsrc : 2'h0)
    | (head[4] ? fb_uop_ram_13_debug_fsrc : 2'h0)
    | (head[5] ? fb_uop_ram_16_debug_fsrc : 2'h0)
    | (head[6] ? fb_uop_ram_19_debug_fsrc : 2'h0)
    | (head[7] ? fb_uop_ram_22_debug_fsrc : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_1_bits_debug_tsrc =
    (head[0] ? fb_uop_ram_1_debug_tsrc : 2'h0)
    | (head[1] ? fb_uop_ram_4_debug_tsrc : 2'h0)
    | (head[2] ? fb_uop_ram_7_debug_tsrc : 2'h0)
    | (head[3] ? fb_uop_ram_10_debug_tsrc : 2'h0)
    | (head[4] ? fb_uop_ram_13_debug_tsrc : 2'h0)
    | (head[5] ? fb_uop_ram_16_debug_tsrc : 2'h0)
    | (head[6] ? fb_uop_ram_19_debug_tsrc : 2'h0)
    | (head[7] ? fb_uop_ram_22_debug_tsrc : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_valid = ~reset & _deq_valids_T_8[2];	// fetch-buffer.scala:161:{21,53}, :168:72, :195:23, :196:41
  assign io_deq_bits_uops_2_bits_inst =
    (head[0] ? fb_uop_ram_2_inst : 32'h0) | (head[1] ? fb_uop_ram_5_inst : 32'h0)
    | (head[2] ? fb_uop_ram_8_inst : 32'h0) | (head[3] ? fb_uop_ram_11_inst : 32'h0)
    | (head[4] ? fb_uop_ram_14_inst : 32'h0) | (head[5] ? fb_uop_ram_17_inst : 32'h0)
    | (head[6] ? fb_uop_ram_20_inst : 32'h0) | (head[7] ? fb_uop_ram_23_inst : 32'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_debug_inst =
    (head[0] ? fb_uop_ram_2_debug_inst : 32'h0)
    | (head[1] ? fb_uop_ram_5_debug_inst : 32'h0)
    | (head[2] ? fb_uop_ram_8_debug_inst : 32'h0)
    | (head[3] ? fb_uop_ram_11_debug_inst : 32'h0)
    | (head[4] ? fb_uop_ram_14_debug_inst : 32'h0)
    | (head[5] ? fb_uop_ram_17_debug_inst : 32'h0)
    | (head[6] ? fb_uop_ram_20_debug_inst : 32'h0)
    | (head[7] ? fb_uop_ram_23_debug_inst : 32'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_is_rvc =
    head[0] & fb_uop_ram_2_is_rvc | head[1] & fb_uop_ram_5_is_rvc | head[2]
    & fb_uop_ram_8_is_rvc | head[3] & fb_uop_ram_11_is_rvc | head[4]
    & fb_uop_ram_14_is_rvc | head[5] & fb_uop_ram_17_is_rvc | head[6]
    & fb_uop_ram_20_is_rvc | head[7] & fb_uop_ram_23_is_rvc;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_debug_pc =
    (head[0] ? fb_uop_ram_2_debug_pc : 40'h0) | (head[1] ? fb_uop_ram_5_debug_pc : 40'h0)
    | (head[2] ? fb_uop_ram_8_debug_pc : 40'h0)
    | (head[3] ? fb_uop_ram_11_debug_pc : 40'h0)
    | (head[4] ? fb_uop_ram_14_debug_pc : 40'h0)
    | (head[5] ? fb_uop_ram_17_debug_pc : 40'h0)
    | (head[6] ? fb_uop_ram_20_debug_pc : 40'h0)
    | (head[7] ? fb_uop_ram_23_debug_pc : 40'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_br_type =
    (head[0] ? fb_uop_ram_2_ctrl_br_type : 4'h0)
    | (head[1] ? fb_uop_ram_5_ctrl_br_type : 4'h0)
    | (head[2] ? fb_uop_ram_8_ctrl_br_type : 4'h0)
    | (head[3] ? fb_uop_ram_11_ctrl_br_type : 4'h0)
    | (head[4] ? fb_uop_ram_14_ctrl_br_type : 4'h0)
    | (head[5] ? fb_uop_ram_17_ctrl_br_type : 4'h0)
    | (head[6] ? fb_uop_ram_20_ctrl_br_type : 4'h0)
    | (head[7] ? fb_uop_ram_23_ctrl_br_type : 4'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_op1_sel =
    (head[0] ? fb_uop_ram_2_ctrl_op1_sel : 2'h0)
    | (head[1] ? fb_uop_ram_5_ctrl_op1_sel : 2'h0)
    | (head[2] ? fb_uop_ram_8_ctrl_op1_sel : 2'h0)
    | (head[3] ? fb_uop_ram_11_ctrl_op1_sel : 2'h0)
    | (head[4] ? fb_uop_ram_14_ctrl_op1_sel : 2'h0)
    | (head[5] ? fb_uop_ram_17_ctrl_op1_sel : 2'h0)
    | (head[6] ? fb_uop_ram_20_ctrl_op1_sel : 2'h0)
    | (head[7] ? fb_uop_ram_23_ctrl_op1_sel : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_op2_sel =
    (head[0] ? fb_uop_ram_2_ctrl_op2_sel : 3'h0)
    | (head[1] ? fb_uop_ram_5_ctrl_op2_sel : 3'h0)
    | (head[2] ? fb_uop_ram_8_ctrl_op2_sel : 3'h0)
    | (head[3] ? fb_uop_ram_11_ctrl_op2_sel : 3'h0)
    | (head[4] ? fb_uop_ram_14_ctrl_op2_sel : 3'h0)
    | (head[5] ? fb_uop_ram_17_ctrl_op2_sel : 3'h0)
    | (head[6] ? fb_uop_ram_20_ctrl_op2_sel : 3'h0)
    | (head[7] ? fb_uop_ram_23_ctrl_op2_sel : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_imm_sel =
    (head[0] ? fb_uop_ram_2_ctrl_imm_sel : 3'h0)
    | (head[1] ? fb_uop_ram_5_ctrl_imm_sel : 3'h0)
    | (head[2] ? fb_uop_ram_8_ctrl_imm_sel : 3'h0)
    | (head[3] ? fb_uop_ram_11_ctrl_imm_sel : 3'h0)
    | (head[4] ? fb_uop_ram_14_ctrl_imm_sel : 3'h0)
    | (head[5] ? fb_uop_ram_17_ctrl_imm_sel : 3'h0)
    | (head[6] ? fb_uop_ram_20_ctrl_imm_sel : 3'h0)
    | (head[7] ? fb_uop_ram_23_ctrl_imm_sel : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_op_fcn =
    (head[0] ? fb_uop_ram_2_ctrl_op_fcn : 4'h0)
    | (head[1] ? fb_uop_ram_5_ctrl_op_fcn : 4'h0)
    | (head[2] ? fb_uop_ram_8_ctrl_op_fcn : 4'h0)
    | (head[3] ? fb_uop_ram_11_ctrl_op_fcn : 4'h0)
    | (head[4] ? fb_uop_ram_14_ctrl_op_fcn : 4'h0)
    | (head[5] ? fb_uop_ram_17_ctrl_op_fcn : 4'h0)
    | (head[6] ? fb_uop_ram_20_ctrl_op_fcn : 4'h0)
    | (head[7] ? fb_uop_ram_23_ctrl_op_fcn : 4'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_fcn_dw =
    head[0] & fb_uop_ram_2_ctrl_fcn_dw | head[1] & fb_uop_ram_5_ctrl_fcn_dw | head[2]
    & fb_uop_ram_8_ctrl_fcn_dw | head[3] & fb_uop_ram_11_ctrl_fcn_dw | head[4]
    & fb_uop_ram_14_ctrl_fcn_dw | head[5] & fb_uop_ram_17_ctrl_fcn_dw | head[6]
    & fb_uop_ram_20_ctrl_fcn_dw | head[7] & fb_uop_ram_23_ctrl_fcn_dw;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_csr_cmd =
    (head[0] ? fb_uop_ram_2_ctrl_csr_cmd : 3'h0)
    | (head[1] ? fb_uop_ram_5_ctrl_csr_cmd : 3'h0)
    | (head[2] ? fb_uop_ram_8_ctrl_csr_cmd : 3'h0)
    | (head[3] ? fb_uop_ram_11_ctrl_csr_cmd : 3'h0)
    | (head[4] ? fb_uop_ram_14_ctrl_csr_cmd : 3'h0)
    | (head[5] ? fb_uop_ram_17_ctrl_csr_cmd : 3'h0)
    | (head[6] ? fb_uop_ram_20_ctrl_csr_cmd : 3'h0)
    | (head[7] ? fb_uop_ram_23_ctrl_csr_cmd : 3'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_is_load =
    head[0] & fb_uop_ram_2_ctrl_is_load | head[1] & fb_uop_ram_5_ctrl_is_load | head[2]
    & fb_uop_ram_8_ctrl_is_load | head[3] & fb_uop_ram_11_ctrl_is_load | head[4]
    & fb_uop_ram_14_ctrl_is_load | head[5] & fb_uop_ram_17_ctrl_is_load | head[6]
    & fb_uop_ram_20_ctrl_is_load | head[7] & fb_uop_ram_23_ctrl_is_load;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_is_sta =
    head[0] & fb_uop_ram_2_ctrl_is_sta | head[1] & fb_uop_ram_5_ctrl_is_sta | head[2]
    & fb_uop_ram_8_ctrl_is_sta | head[3] & fb_uop_ram_11_ctrl_is_sta | head[4]
    & fb_uop_ram_14_ctrl_is_sta | head[5] & fb_uop_ram_17_ctrl_is_sta | head[6]
    & fb_uop_ram_20_ctrl_is_sta | head[7] & fb_uop_ram_23_ctrl_is_sta;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_ctrl_is_std =
    head[0] & fb_uop_ram_2_ctrl_is_std | head[1] & fb_uop_ram_5_ctrl_is_std | head[2]
    & fb_uop_ram_8_ctrl_is_std | head[3] & fb_uop_ram_11_ctrl_is_std | head[4]
    & fb_uop_ram_14_ctrl_is_std | head[5] & fb_uop_ram_17_ctrl_is_std | head[6]
    & fb_uop_ram_20_ctrl_is_std | head[7] & fb_uop_ram_23_ctrl_is_std;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_iw_state =
    (head[0] ? fb_uop_ram_2_iw_state : 2'h0) | (head[1] ? fb_uop_ram_5_iw_state : 2'h0)
    | (head[2] ? fb_uop_ram_8_iw_state : 2'h0) | (head[3] ? fb_uop_ram_11_iw_state : 2'h0)
    | (head[4] ? fb_uop_ram_14_iw_state : 2'h0)
    | (head[5] ? fb_uop_ram_17_iw_state : 2'h0)
    | (head[6] ? fb_uop_ram_20_iw_state : 2'h0)
    | (head[7] ? fb_uop_ram_23_iw_state : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_iw_p1_poisoned =
    head[0] & fb_uop_ram_2_iw_p1_poisoned | head[1] & fb_uop_ram_5_iw_p1_poisoned
    | head[2] & fb_uop_ram_8_iw_p1_poisoned | head[3] & fb_uop_ram_11_iw_p1_poisoned
    | head[4] & fb_uop_ram_14_iw_p1_poisoned | head[5] & fb_uop_ram_17_iw_p1_poisoned
    | head[6] & fb_uop_ram_20_iw_p1_poisoned | head[7] & fb_uop_ram_23_iw_p1_poisoned;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_iw_p2_poisoned =
    head[0] & fb_uop_ram_2_iw_p2_poisoned | head[1] & fb_uop_ram_5_iw_p2_poisoned
    | head[2] & fb_uop_ram_8_iw_p2_poisoned | head[3] & fb_uop_ram_11_iw_p2_poisoned
    | head[4] & fb_uop_ram_14_iw_p2_poisoned | head[5] & fb_uop_ram_17_iw_p2_poisoned
    | head[6] & fb_uop_ram_20_iw_p2_poisoned | head[7] & fb_uop_ram_23_iw_p2_poisoned;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_is_sfb =
    head[0] & fb_uop_ram_2_is_sfb | head[1] & fb_uop_ram_5_is_sfb | head[2]
    & fb_uop_ram_8_is_sfb | head[3] & fb_uop_ram_11_is_sfb | head[4]
    & fb_uop_ram_14_is_sfb | head[5] & fb_uop_ram_17_is_sfb | head[6]
    & fb_uop_ram_20_is_sfb | head[7] & fb_uop_ram_23_is_sfb;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_ftq_idx =
    (head[0] ? fb_uop_ram_2_ftq_idx : 5'h0) | (head[1] ? fb_uop_ram_5_ftq_idx : 5'h0)
    | (head[2] ? fb_uop_ram_8_ftq_idx : 5'h0) | (head[3] ? fb_uop_ram_11_ftq_idx : 5'h0)
    | (head[4] ? fb_uop_ram_14_ftq_idx : 5'h0) | (head[5] ? fb_uop_ram_17_ftq_idx : 5'h0)
    | (head[6] ? fb_uop_ram_20_ftq_idx : 5'h0) | (head[7] ? fb_uop_ram_23_ftq_idx : 5'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_edge_inst =
    head[0] & fb_uop_ram_2_edge_inst | head[1] & fb_uop_ram_5_edge_inst | head[2]
    & fb_uop_ram_8_edge_inst | head[3] & fb_uop_ram_11_edge_inst | head[4]
    & fb_uop_ram_14_edge_inst | head[5] & fb_uop_ram_17_edge_inst | head[6]
    & fb_uop_ram_20_edge_inst | head[7] & fb_uop_ram_23_edge_inst;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_pc_lob =
    (head[0] ? fb_uop_ram_2_pc_lob : 6'h0) | (head[1] ? fb_uop_ram_5_pc_lob : 6'h0)
    | (head[2] ? fb_uop_ram_8_pc_lob : 6'h0) | (head[3] ? fb_uop_ram_11_pc_lob : 6'h0)
    | (head[4] ? fb_uop_ram_14_pc_lob : 6'h0) | (head[5] ? fb_uop_ram_17_pc_lob : 6'h0)
    | (head[6] ? fb_uop_ram_20_pc_lob : 6'h0) | (head[7] ? fb_uop_ram_23_pc_lob : 6'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_taken =
    head[0] & fb_uop_ram_2_taken | head[1] & fb_uop_ram_5_taken | head[2]
    & fb_uop_ram_8_taken | head[3] & fb_uop_ram_11_taken | head[4] & fb_uop_ram_14_taken
    | head[5] & fb_uop_ram_17_taken | head[6] & fb_uop_ram_20_taken | head[7]
    & fb_uop_ram_23_taken;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_csr_addr =
    (head[0] ? fb_uop_ram_2_csr_addr : 12'h0) | (head[1] ? fb_uop_ram_5_csr_addr : 12'h0)
    | (head[2] ? fb_uop_ram_8_csr_addr : 12'h0)
    | (head[3] ? fb_uop_ram_11_csr_addr : 12'h0)
    | (head[4] ? fb_uop_ram_14_csr_addr : 12'h0)
    | (head[5] ? fb_uop_ram_17_csr_addr : 12'h0)
    | (head[6] ? fb_uop_ram_20_csr_addr : 12'h0)
    | (head[7] ? fb_uop_ram_23_csr_addr : 12'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_rxq_idx =
    (head[0] ? fb_uop_ram_2_rxq_idx : 2'h0) | (head[1] ? fb_uop_ram_5_rxq_idx : 2'h0)
    | (head[2] ? fb_uop_ram_8_rxq_idx : 2'h0) | (head[3] ? fb_uop_ram_11_rxq_idx : 2'h0)
    | (head[4] ? fb_uop_ram_14_rxq_idx : 2'h0) | (head[5] ? fb_uop_ram_17_rxq_idx : 2'h0)
    | (head[6] ? fb_uop_ram_20_rxq_idx : 2'h0) | (head[7] ? fb_uop_ram_23_rxq_idx : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_xcpt_pf_if =
    head[0] & fb_uop_ram_2_xcpt_pf_if | head[1] & fb_uop_ram_5_xcpt_pf_if | head[2]
    & fb_uop_ram_8_xcpt_pf_if | head[3] & fb_uop_ram_11_xcpt_pf_if | head[4]
    & fb_uop_ram_14_xcpt_pf_if | head[5] & fb_uop_ram_17_xcpt_pf_if | head[6]
    & fb_uop_ram_20_xcpt_pf_if | head[7] & fb_uop_ram_23_xcpt_pf_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_xcpt_ae_if =
    head[0] & fb_uop_ram_2_xcpt_ae_if | head[1] & fb_uop_ram_5_xcpt_ae_if | head[2]
    & fb_uop_ram_8_xcpt_ae_if | head[3] & fb_uop_ram_11_xcpt_ae_if | head[4]
    & fb_uop_ram_14_xcpt_ae_if | head[5] & fb_uop_ram_17_xcpt_ae_if | head[6]
    & fb_uop_ram_20_xcpt_ae_if | head[7] & fb_uop_ram_23_xcpt_ae_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_xcpt_ma_if =
    head[0] & fb_uop_ram_2_xcpt_ma_if | head[1] & fb_uop_ram_5_xcpt_ma_if | head[2]
    & fb_uop_ram_8_xcpt_ma_if | head[3] & fb_uop_ram_11_xcpt_ma_if | head[4]
    & fb_uop_ram_14_xcpt_ma_if | head[5] & fb_uop_ram_17_xcpt_ma_if | head[6]
    & fb_uop_ram_20_xcpt_ma_if | head[7] & fb_uop_ram_23_xcpt_ma_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_bp_debug_if =
    head[0] & fb_uop_ram_2_bp_debug_if | head[1] & fb_uop_ram_5_bp_debug_if | head[2]
    & fb_uop_ram_8_bp_debug_if | head[3] & fb_uop_ram_11_bp_debug_if | head[4]
    & fb_uop_ram_14_bp_debug_if | head[5] & fb_uop_ram_17_bp_debug_if | head[6]
    & fb_uop_ram_20_bp_debug_if | head[7] & fb_uop_ram_23_bp_debug_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_bp_xcpt_if =
    head[0] & fb_uop_ram_2_bp_xcpt_if | head[1] & fb_uop_ram_5_bp_xcpt_if | head[2]
    & fb_uop_ram_8_bp_xcpt_if | head[3] & fb_uop_ram_11_bp_xcpt_if | head[4]
    & fb_uop_ram_14_bp_xcpt_if | head[5] & fb_uop_ram_17_bp_xcpt_if | head[6]
    & fb_uop_ram_20_bp_xcpt_if | head[7] & fb_uop_ram_23_bp_xcpt_if;	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :155:31
  assign io_deq_bits_uops_2_bits_debug_fsrc =
    (head[0] ? fb_uop_ram_2_debug_fsrc : 2'h0)
    | (head[1] ? fb_uop_ram_5_debug_fsrc : 2'h0)
    | (head[2] ? fb_uop_ram_8_debug_fsrc : 2'h0)
    | (head[3] ? fb_uop_ram_11_debug_fsrc : 2'h0)
    | (head[4] ? fb_uop_ram_14_debug_fsrc : 2'h0)
    | (head[5] ? fb_uop_ram_17_debug_fsrc : 2'h0)
    | (head[6] ? fb_uop_ram_20_debug_fsrc : 2'h0)
    | (head[7] ? fb_uop_ram_23_debug_fsrc : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
  assign io_deq_bits_uops_2_bits_debug_tsrc =
    (head[0] ? fb_uop_ram_2_debug_tsrc : 2'h0)
    | (head[1] ? fb_uop_ram_5_debug_tsrc : 2'h0)
    | (head[2] ? fb_uop_ram_8_debug_tsrc : 2'h0)
    | (head[3] ? fb_uop_ram_11_debug_tsrc : 2'h0)
    | (head[4] ? fb_uop_ram_14_debug_tsrc : 2'h0)
    | (head[5] ? fb_uop_ram_17_debug_tsrc : 2'h0)
    | (head[6] ? fb_uop_ram_20_debug_tsrc : 2'h0)
    | (head[7] ? fb_uop_ram_23_debug_tsrc : 2'h0);	// Mux.scala:27:72, fetch-buffer.scala:57:16, :61:21, :97:33, :155:31
endmodule

