// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module RoundAnyRawFNToRecFN_2(
  input         io_in_isZero,
                io_in_sign,
  input  [8:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags
);

  wire        roundingMode_near_even = io_roundingMode == 3'h0;	// RoundAnyRawFNToRecFN.scala:88:53
  wire        common_inexact = io_in_sig[10] | (|(io_in_sig[9:0]));	// RoundAnyRawFNToRecFN.scala:115:{26,60}, :162:40, :164:36
  wire [54:0] roundedSig =
    (roundingMode_near_even | io_roundingMode == 3'h4) & io_in_sig[10]
    | (io_roundingMode == 3'h2 & io_in_sign | io_roundingMode == 3'h3 & ~io_in_sign)
    & common_inexact
      ? {1'h0, io_in_sig[64:11]} + 55'h1
        & {54'h3FFFFFFFFFFFFF,
           ~(roundingMode_near_even & io_in_sig[10] & ~(|(io_in_sig[9:0])))}
      : {1'h0,
         io_in_sig[64:12],
         io_in_sig[11] | io_roundingMode == 3'h6 & common_inexact};	// Cat.scala:30:58, RoundAnyRawFNToRecFN.scala:88:53, :90:53, :91:53, :92:53, :93:53, :96:{27,42,63,66}, :104:31, :115:{26,60}, :160:57, :162:40, :164:36, :167:{38,67}, :168:31, :169:29, :171:16, :172:{49,61}, :173:{21,25,64}, :174:30, :178:47, :179:42
  assign io_out =
    {io_in_sign,
     {{3{io_in_sExp[8]}}, io_in_sExp} + {10'h0, roundedSig[54:53]} + 12'h780
       & ~(io_in_isZero ? 12'hE00 : 12'h0),
     io_in_isZero ? 52'h0 : roundedSig[51:0]};	// Cat.scala:30:58, RoundAnyRawFNToRecFN.scala:102:25, :115:60, :171:16, :183:{40,54}, :189:27, :250:24, :251:{14,18}, :275:16, :276:16, :278:12, :279:16
  assign io_exceptionFlags = {4'h0, ~io_in_isZero & common_inexact};	// Cat.scala:30:58, RoundAnyRawFNToRecFN.scala:164:36, :235:64, :238:43
endmodule

