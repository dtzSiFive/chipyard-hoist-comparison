// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module Rob(
  input         clock,
                reset,
                io_enq_valids_0,
                io_enq_valids_1,
                io_enq_valids_2,
                io_enq_valids_3,
  input  [6:0]  io_enq_uops_0_uopc,
  input         io_enq_uops_0_is_rvc,
                io_enq_uops_0_is_br,
                io_enq_uops_0_is_jalr,
  input  [19:0] io_enq_uops_0_br_mask,
  input  [5:0]  io_enq_uops_0_ftq_idx,
  input         io_enq_uops_0_edge_inst,
  input  [5:0]  io_enq_uops_0_pc_lob,
  input  [6:0]  io_enq_uops_0_rob_idx,
                io_enq_uops_0_pdst,
                io_enq_uops_0_stale_pdst,
  input         io_enq_uops_0_exception,
  input  [63:0] io_enq_uops_0_exc_cause,
  input         io_enq_uops_0_is_fence,
                io_enq_uops_0_is_fencei,
                io_enq_uops_0_uses_ldq,
                io_enq_uops_0_uses_stq,
                io_enq_uops_0_is_sys_pc2epc,
                io_enq_uops_0_is_unique,
                io_enq_uops_0_flush_on_commit,
  input  [5:0]  io_enq_uops_0_ldst,
  input         io_enq_uops_0_ldst_val,
  input  [1:0]  io_enq_uops_0_dst_rtype,
  input         io_enq_uops_0_fp_val,
  input  [6:0]  io_enq_uops_1_uopc,
  input         io_enq_uops_1_is_rvc,
                io_enq_uops_1_is_br,
                io_enq_uops_1_is_jalr,
  input  [19:0] io_enq_uops_1_br_mask,
  input  [5:0]  io_enq_uops_1_ftq_idx,
  input         io_enq_uops_1_edge_inst,
  input  [5:0]  io_enq_uops_1_pc_lob,
  input  [6:0]  io_enq_uops_1_rob_idx,
                io_enq_uops_1_pdst,
                io_enq_uops_1_stale_pdst,
  input         io_enq_uops_1_exception,
  input  [63:0] io_enq_uops_1_exc_cause,
  input         io_enq_uops_1_is_fence,
                io_enq_uops_1_is_fencei,
                io_enq_uops_1_uses_ldq,
                io_enq_uops_1_uses_stq,
                io_enq_uops_1_is_sys_pc2epc,
                io_enq_uops_1_is_unique,
                io_enq_uops_1_flush_on_commit,
  input  [5:0]  io_enq_uops_1_ldst,
  input         io_enq_uops_1_ldst_val,
  input  [1:0]  io_enq_uops_1_dst_rtype,
  input         io_enq_uops_1_fp_val,
  input  [6:0]  io_enq_uops_2_uopc,
  input         io_enq_uops_2_is_rvc,
                io_enq_uops_2_is_br,
                io_enq_uops_2_is_jalr,
  input  [19:0] io_enq_uops_2_br_mask,
  input  [5:0]  io_enq_uops_2_ftq_idx,
  input         io_enq_uops_2_edge_inst,
  input  [5:0]  io_enq_uops_2_pc_lob,
  input  [6:0]  io_enq_uops_2_rob_idx,
                io_enq_uops_2_pdst,
                io_enq_uops_2_stale_pdst,
  input         io_enq_uops_2_exception,
  input  [63:0] io_enq_uops_2_exc_cause,
  input         io_enq_uops_2_is_fence,
                io_enq_uops_2_is_fencei,
                io_enq_uops_2_uses_ldq,
                io_enq_uops_2_uses_stq,
                io_enq_uops_2_is_sys_pc2epc,
                io_enq_uops_2_is_unique,
                io_enq_uops_2_flush_on_commit,
  input  [5:0]  io_enq_uops_2_ldst,
  input         io_enq_uops_2_ldst_val,
  input  [1:0]  io_enq_uops_2_dst_rtype,
  input         io_enq_uops_2_fp_val,
  input  [6:0]  io_enq_uops_3_uopc,
  input         io_enq_uops_3_is_rvc,
                io_enq_uops_3_is_br,
                io_enq_uops_3_is_jalr,
  input  [19:0] io_enq_uops_3_br_mask,
  input  [5:0]  io_enq_uops_3_ftq_idx,
  input         io_enq_uops_3_edge_inst,
  input  [5:0]  io_enq_uops_3_pc_lob,
  input  [6:0]  io_enq_uops_3_rob_idx,
                io_enq_uops_3_pdst,
                io_enq_uops_3_stale_pdst,
  input         io_enq_uops_3_exception,
  input  [63:0] io_enq_uops_3_exc_cause,
  input         io_enq_uops_3_is_fence,
                io_enq_uops_3_is_fencei,
                io_enq_uops_3_uses_ldq,
                io_enq_uops_3_uses_stq,
                io_enq_uops_3_is_sys_pc2epc,
                io_enq_uops_3_is_unique,
                io_enq_uops_3_flush_on_commit,
  input  [5:0]  io_enq_uops_3_ldst,
  input         io_enq_uops_3_ldst_val,
  input  [1:0]  io_enq_uops_3_dst_rtype,
  input         io_enq_uops_3_fp_val,
                io_enq_partial_stall,
  input  [39:0] io_xcpt_fetch_pc,
  input  [19:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input  [6:0]  io_brupdate_b2_uop_rob_idx,
  input         io_brupdate_b2_mispredict,
                io_wb_resps_0_valid,
  input  [6:0]  io_wb_resps_0_bits_uop_rob_idx,
                io_wb_resps_0_bits_uop_pdst,
  input         io_wb_resps_0_bits_predicated,
                io_wb_resps_1_valid,
  input  [6:0]  io_wb_resps_1_bits_uop_rob_idx,
                io_wb_resps_1_bits_uop_pdst,
  input         io_wb_resps_2_valid,
  input  [6:0]  io_wb_resps_2_bits_uop_rob_idx,
                io_wb_resps_2_bits_uop_pdst,
  input         io_wb_resps_3_valid,
  input  [6:0]  io_wb_resps_3_bits_uop_rob_idx,
                io_wb_resps_3_bits_uop_pdst,
  input         io_wb_resps_4_valid,
  input  [6:0]  io_wb_resps_4_bits_uop_rob_idx,
                io_wb_resps_4_bits_uop_pdst,
  input         io_wb_resps_5_valid,
  input  [6:0]  io_wb_resps_5_bits_uop_rob_idx,
                io_wb_resps_5_bits_uop_pdst,
  input         io_wb_resps_6_valid,
  input  [6:0]  io_wb_resps_6_bits_uop_rob_idx,
                io_wb_resps_6_bits_uop_pdst,
  input         io_wb_resps_6_bits_predicated,
                io_wb_resps_7_valid,
  input  [6:0]  io_wb_resps_7_bits_uop_rob_idx,
                io_wb_resps_7_bits_uop_pdst,
  input         io_wb_resps_8_valid,
  input  [6:0]  io_wb_resps_8_bits_uop_rob_idx,
                io_wb_resps_8_bits_uop_pdst,
  input         io_wb_resps_9_valid,
  input  [6:0]  io_wb_resps_9_bits_uop_rob_idx,
                io_wb_resps_9_bits_uop_pdst,
  input         io_lsu_clr_bsy_0_valid,
  input  [6:0]  io_lsu_clr_bsy_0_bits,
  input         io_lsu_clr_bsy_1_valid,
  input  [6:0]  io_lsu_clr_bsy_1_bits,
  input         io_lsu_clr_bsy_2_valid,
  input  [6:0]  io_lsu_clr_bsy_2_bits,
  input         io_fflags_0_valid,
  input  [6:0]  io_fflags_0_bits_uop_rob_idx,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_2_valid,
  input  [6:0]  io_fflags_2_bits_uop_rob_idx,
  input  [4:0]  io_fflags_2_bits_flags,
  input         io_fflags_3_valid,
  input  [6:0]  io_fflags_3_bits_uop_rob_idx,
  input  [4:0]  io_fflags_3_bits_flags,
  input         io_lxcpt_valid,
  input  [19:0] io_lxcpt_bits_uop_br_mask,
  input  [6:0]  io_lxcpt_bits_uop_rob_idx,
  input  [4:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  input         io_csr_stall,
  output [6:0]  io_rob_tail_idx,
                io_rob_head_idx,
  output        io_commit_valids_0,
                io_commit_valids_1,
                io_commit_valids_2,
                io_commit_valids_3,
                io_commit_arch_valids_0,
                io_commit_arch_valids_1,
                io_commit_arch_valids_2,
                io_commit_arch_valids_3,
  output [5:0]  io_commit_uops_0_ftq_idx,
  output [6:0]  io_commit_uops_0_pdst,
                io_commit_uops_0_stale_pdst,
  output        io_commit_uops_0_is_fencei,
                io_commit_uops_0_uses_ldq,
                io_commit_uops_0_uses_stq,
  output [5:0]  io_commit_uops_0_ldst,
  output        io_commit_uops_0_ldst_val,
  output [1:0]  io_commit_uops_0_dst_rtype,
  output [5:0]  io_commit_uops_1_ftq_idx,
  output [6:0]  io_commit_uops_1_pdst,
                io_commit_uops_1_stale_pdst,
  output        io_commit_uops_1_is_fencei,
                io_commit_uops_1_uses_ldq,
                io_commit_uops_1_uses_stq,
  output [5:0]  io_commit_uops_1_ldst,
  output        io_commit_uops_1_ldst_val,
  output [1:0]  io_commit_uops_1_dst_rtype,
  output [5:0]  io_commit_uops_2_ftq_idx,
  output [6:0]  io_commit_uops_2_pdst,
                io_commit_uops_2_stale_pdst,
  output        io_commit_uops_2_is_fencei,
                io_commit_uops_2_uses_ldq,
                io_commit_uops_2_uses_stq,
  output [5:0]  io_commit_uops_2_ldst,
  output        io_commit_uops_2_ldst_val,
  output [1:0]  io_commit_uops_2_dst_rtype,
  output [5:0]  io_commit_uops_3_ftq_idx,
  output [6:0]  io_commit_uops_3_pdst,
                io_commit_uops_3_stale_pdst,
  output        io_commit_uops_3_is_fencei,
                io_commit_uops_3_uses_ldq,
                io_commit_uops_3_uses_stq,
  output [5:0]  io_commit_uops_3_ldst,
  output        io_commit_uops_3_ldst_val,
  output [1:0]  io_commit_uops_3_dst_rtype,
  output        io_commit_fflags_valid,
  output [4:0]  io_commit_fflags_bits,
  output        io_commit_rbk_valids_0,
                io_commit_rbk_valids_1,
                io_commit_rbk_valids_2,
                io_commit_rbk_valids_3,
                io_commit_rollback,
                io_com_load_is_at_rob_head,
                io_com_xcpt_valid,
  output [5:0]  io_com_xcpt_bits_ftq_idx,
  output        io_com_xcpt_bits_edge_inst,
  output [5:0]  io_com_xcpt_bits_pc_lob,
  output [63:0] io_com_xcpt_bits_cause,
                io_com_xcpt_bits_badvaddr,
  output        io_flush_valid,
  output [5:0]  io_flush_bits_ftq_idx,
  output        io_flush_bits_edge_inst,
                io_flush_bits_is_rvc,
  output [5:0]  io_flush_bits_pc_lob,
  output [2:0]  io_flush_bits_flush_typ,
  output        io_empty,
                io_ready,
                io_flush_frontend
);

  wire             empty;	// rob.scala:788:41
  wire             full;	// rob.scala:787:39
  wire             will_commit_3;	// rob.scala:547:70
  wire             will_commit_2;	// rob.scala:547:70
  wire             will_commit_1;	// rob.scala:547:70
  wire             will_commit_0;	// rob.scala:547:70
  wire [4:0]       _rob_fflags_3_ext_R0_data;	// rob.scala:313:28
  wire [4:0]       _rob_fflags_2_ext_R0_data;	// rob.scala:313:28
  wire [4:0]       _rob_fflags_1_ext_R0_data;	// rob.scala:313:28
  wire [4:0]       _rob_fflags_ext_R0_data;	// rob.scala:313:28
  reg  [1:0]       rob_state;	// rob.scala:221:26
  reg  [4:0]       rob_head;	// rob.scala:224:29
  reg  [1:0]       rob_head_lsb;	// rob.scala:225:29
  wire [6:0]       rob_head_idx = {rob_head, rob_head_lsb};	// Cat.scala:30:58, rob.scala:224:29, :225:29
  reg  [4:0]       rob_tail;	// rob.scala:228:29
  reg  [1:0]       rob_tail_lsb;	// rob.scala:229:29
  wire [6:0]       rob_tail_idx = {rob_tail, rob_tail_lsb};	// Cat.scala:30:58, rob.scala:228:29, :229:29
  reg  [4:0]       rob_pnr;	// rob.scala:232:29
  reg  [1:0]       rob_pnr_lsb;	// rob.scala:233:29
  wire             _io_commit_rollback_T_3 = rob_state == 2'h2;	// rob.scala:221:26, :236:31
  wire [4:0]       com_idx = _io_commit_rollback_T_3 ? rob_tail : rob_head;	// rob.scala:224:29, :228:29, :236:{20,31}
  reg              maybe_full;	// rob.scala:239:29
  reg              r_xcpt_val;	// rob.scala:258:33
  reg  [19:0]      r_xcpt_uop_br_mask;	// rob.scala:259:29
  reg  [6:0]       r_xcpt_uop_rob_idx;	// rob.scala:259:29
  reg  [63:0]      r_xcpt_uop_exc_cause;	// rob.scala:259:29
  reg  [39:0]      r_xcpt_badvaddr;	// rob.scala:260:29
  reg              rob_val_0;	// rob.scala:307:32
  reg              rob_val_1;	// rob.scala:307:32
  reg              rob_val_2;	// rob.scala:307:32
  reg              rob_val_3;	// rob.scala:307:32
  reg              rob_val_4;	// rob.scala:307:32
  reg              rob_val_5;	// rob.scala:307:32
  reg              rob_val_6;	// rob.scala:307:32
  reg              rob_val_7;	// rob.scala:307:32
  reg              rob_val_8;	// rob.scala:307:32
  reg              rob_val_9;	// rob.scala:307:32
  reg              rob_val_10;	// rob.scala:307:32
  reg              rob_val_11;	// rob.scala:307:32
  reg              rob_val_12;	// rob.scala:307:32
  reg              rob_val_13;	// rob.scala:307:32
  reg              rob_val_14;	// rob.scala:307:32
  reg              rob_val_15;	// rob.scala:307:32
  reg              rob_val_16;	// rob.scala:307:32
  reg              rob_val_17;	// rob.scala:307:32
  reg              rob_val_18;	// rob.scala:307:32
  reg              rob_val_19;	// rob.scala:307:32
  reg              rob_val_20;	// rob.scala:307:32
  reg              rob_val_21;	// rob.scala:307:32
  reg              rob_val_22;	// rob.scala:307:32
  reg              rob_val_23;	// rob.scala:307:32
  reg              rob_val_24;	// rob.scala:307:32
  reg              rob_val_25;	// rob.scala:307:32
  reg              rob_val_26;	// rob.scala:307:32
  reg              rob_val_27;	// rob.scala:307:32
  reg              rob_val_28;	// rob.scala:307:32
  reg              rob_val_29;	// rob.scala:307:32
  reg              rob_val_30;	// rob.scala:307:32
  reg              rob_val_31;	// rob.scala:307:32
  reg              rob_bsy_0;	// rob.scala:308:28
  reg              rob_bsy_1;	// rob.scala:308:28
  reg              rob_bsy_2;	// rob.scala:308:28
  reg              rob_bsy_3;	// rob.scala:308:28
  reg              rob_bsy_4;	// rob.scala:308:28
  reg              rob_bsy_5;	// rob.scala:308:28
  reg              rob_bsy_6;	// rob.scala:308:28
  reg              rob_bsy_7;	// rob.scala:308:28
  reg              rob_bsy_8;	// rob.scala:308:28
  reg              rob_bsy_9;	// rob.scala:308:28
  reg              rob_bsy_10;	// rob.scala:308:28
  reg              rob_bsy_11;	// rob.scala:308:28
  reg              rob_bsy_12;	// rob.scala:308:28
  reg              rob_bsy_13;	// rob.scala:308:28
  reg              rob_bsy_14;	// rob.scala:308:28
  reg              rob_bsy_15;	// rob.scala:308:28
  reg              rob_bsy_16;	// rob.scala:308:28
  reg              rob_bsy_17;	// rob.scala:308:28
  reg              rob_bsy_18;	// rob.scala:308:28
  reg              rob_bsy_19;	// rob.scala:308:28
  reg              rob_bsy_20;	// rob.scala:308:28
  reg              rob_bsy_21;	// rob.scala:308:28
  reg              rob_bsy_22;	// rob.scala:308:28
  reg              rob_bsy_23;	// rob.scala:308:28
  reg              rob_bsy_24;	// rob.scala:308:28
  reg              rob_bsy_25;	// rob.scala:308:28
  reg              rob_bsy_26;	// rob.scala:308:28
  reg              rob_bsy_27;	// rob.scala:308:28
  reg              rob_bsy_28;	// rob.scala:308:28
  reg              rob_bsy_29;	// rob.scala:308:28
  reg              rob_bsy_30;	// rob.scala:308:28
  reg              rob_bsy_31;	// rob.scala:308:28
  reg              rob_unsafe_0;	// rob.scala:309:28
  reg              rob_unsafe_1;	// rob.scala:309:28
  reg              rob_unsafe_2;	// rob.scala:309:28
  reg              rob_unsafe_3;	// rob.scala:309:28
  reg              rob_unsafe_4;	// rob.scala:309:28
  reg              rob_unsafe_5;	// rob.scala:309:28
  reg              rob_unsafe_6;	// rob.scala:309:28
  reg              rob_unsafe_7;	// rob.scala:309:28
  reg              rob_unsafe_8;	// rob.scala:309:28
  reg              rob_unsafe_9;	// rob.scala:309:28
  reg              rob_unsafe_10;	// rob.scala:309:28
  reg              rob_unsafe_11;	// rob.scala:309:28
  reg              rob_unsafe_12;	// rob.scala:309:28
  reg              rob_unsafe_13;	// rob.scala:309:28
  reg              rob_unsafe_14;	// rob.scala:309:28
  reg              rob_unsafe_15;	// rob.scala:309:28
  reg              rob_unsafe_16;	// rob.scala:309:28
  reg              rob_unsafe_17;	// rob.scala:309:28
  reg              rob_unsafe_18;	// rob.scala:309:28
  reg              rob_unsafe_19;	// rob.scala:309:28
  reg              rob_unsafe_20;	// rob.scala:309:28
  reg              rob_unsafe_21;	// rob.scala:309:28
  reg              rob_unsafe_22;	// rob.scala:309:28
  reg              rob_unsafe_23;	// rob.scala:309:28
  reg              rob_unsafe_24;	// rob.scala:309:28
  reg              rob_unsafe_25;	// rob.scala:309:28
  reg              rob_unsafe_26;	// rob.scala:309:28
  reg              rob_unsafe_27;	// rob.scala:309:28
  reg              rob_unsafe_28;	// rob.scala:309:28
  reg              rob_unsafe_29;	// rob.scala:309:28
  reg              rob_unsafe_30;	// rob.scala:309:28
  reg              rob_unsafe_31;	// rob.scala:309:28
  reg  [6:0]       rob_uop_0_uopc;	// rob.scala:310:28
  reg              rob_uop_0_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_0_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_0_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_0_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_0_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_0_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_0_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_0_is_fencei;	// rob.scala:310:28
  reg              rob_uop_0_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_0_uses_stq;	// rob.scala:310:28
  reg              rob_uop_0_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_0_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_0_ldst;	// rob.scala:310:28
  reg              rob_uop_0_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_0_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_0_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_uopc;	// rob.scala:310:28
  reg              rob_uop_1_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_ldst;	// rob.scala:310:28
  reg              rob_uop_1_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_uopc;	// rob.scala:310:28
  reg              rob_uop_2_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_ldst;	// rob.scala:310:28
  reg              rob_uop_2_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_uopc;	// rob.scala:310:28
  reg              rob_uop_3_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_ldst;	// rob.scala:310:28
  reg              rob_uop_3_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_4_uopc;	// rob.scala:310:28
  reg              rob_uop_4_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_4_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_4_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_4_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_4_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_4_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_4_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_4_is_fencei;	// rob.scala:310:28
  reg              rob_uop_4_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_4_uses_stq;	// rob.scala:310:28
  reg              rob_uop_4_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_4_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_4_ldst;	// rob.scala:310:28
  reg              rob_uop_4_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_4_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_4_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_5_uopc;	// rob.scala:310:28
  reg              rob_uop_5_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_5_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_5_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_5_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_5_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_5_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_5_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_5_is_fencei;	// rob.scala:310:28
  reg              rob_uop_5_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_5_uses_stq;	// rob.scala:310:28
  reg              rob_uop_5_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_5_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_5_ldst;	// rob.scala:310:28
  reg              rob_uop_5_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_5_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_5_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_6_uopc;	// rob.scala:310:28
  reg              rob_uop_6_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_6_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_6_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_6_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_6_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_6_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_6_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_6_is_fencei;	// rob.scala:310:28
  reg              rob_uop_6_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_6_uses_stq;	// rob.scala:310:28
  reg              rob_uop_6_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_6_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_6_ldst;	// rob.scala:310:28
  reg              rob_uop_6_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_6_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_6_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_7_uopc;	// rob.scala:310:28
  reg              rob_uop_7_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_7_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_7_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_7_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_7_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_7_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_7_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_7_is_fencei;	// rob.scala:310:28
  reg              rob_uop_7_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_7_uses_stq;	// rob.scala:310:28
  reg              rob_uop_7_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_7_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_7_ldst;	// rob.scala:310:28
  reg              rob_uop_7_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_7_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_7_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_8_uopc;	// rob.scala:310:28
  reg              rob_uop_8_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_8_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_8_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_8_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_8_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_8_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_8_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_8_is_fencei;	// rob.scala:310:28
  reg              rob_uop_8_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_8_uses_stq;	// rob.scala:310:28
  reg              rob_uop_8_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_8_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_8_ldst;	// rob.scala:310:28
  reg              rob_uop_8_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_8_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_8_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_9_uopc;	// rob.scala:310:28
  reg              rob_uop_9_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_9_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_9_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_9_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_9_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_9_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_9_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_9_is_fencei;	// rob.scala:310:28
  reg              rob_uop_9_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_9_uses_stq;	// rob.scala:310:28
  reg              rob_uop_9_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_9_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_9_ldst;	// rob.scala:310:28
  reg              rob_uop_9_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_9_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_9_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_10_uopc;	// rob.scala:310:28
  reg              rob_uop_10_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_10_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_10_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_10_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_10_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_10_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_10_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_10_is_fencei;	// rob.scala:310:28
  reg              rob_uop_10_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_10_uses_stq;	// rob.scala:310:28
  reg              rob_uop_10_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_10_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_10_ldst;	// rob.scala:310:28
  reg              rob_uop_10_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_10_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_10_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_11_uopc;	// rob.scala:310:28
  reg              rob_uop_11_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_11_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_11_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_11_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_11_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_11_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_11_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_11_is_fencei;	// rob.scala:310:28
  reg              rob_uop_11_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_11_uses_stq;	// rob.scala:310:28
  reg              rob_uop_11_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_11_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_11_ldst;	// rob.scala:310:28
  reg              rob_uop_11_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_11_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_11_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_12_uopc;	// rob.scala:310:28
  reg              rob_uop_12_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_12_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_12_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_12_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_12_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_12_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_12_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_12_is_fencei;	// rob.scala:310:28
  reg              rob_uop_12_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_12_uses_stq;	// rob.scala:310:28
  reg              rob_uop_12_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_12_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_12_ldst;	// rob.scala:310:28
  reg              rob_uop_12_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_12_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_12_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_13_uopc;	// rob.scala:310:28
  reg              rob_uop_13_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_13_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_13_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_13_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_13_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_13_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_13_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_13_is_fencei;	// rob.scala:310:28
  reg              rob_uop_13_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_13_uses_stq;	// rob.scala:310:28
  reg              rob_uop_13_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_13_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_13_ldst;	// rob.scala:310:28
  reg              rob_uop_13_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_13_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_13_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_14_uopc;	// rob.scala:310:28
  reg              rob_uop_14_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_14_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_14_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_14_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_14_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_14_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_14_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_14_is_fencei;	// rob.scala:310:28
  reg              rob_uop_14_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_14_uses_stq;	// rob.scala:310:28
  reg              rob_uop_14_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_14_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_14_ldst;	// rob.scala:310:28
  reg              rob_uop_14_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_14_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_14_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_15_uopc;	// rob.scala:310:28
  reg              rob_uop_15_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_15_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_15_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_15_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_15_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_15_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_15_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_15_is_fencei;	// rob.scala:310:28
  reg              rob_uop_15_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_15_uses_stq;	// rob.scala:310:28
  reg              rob_uop_15_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_15_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_15_ldst;	// rob.scala:310:28
  reg              rob_uop_15_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_15_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_15_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_16_uopc;	// rob.scala:310:28
  reg              rob_uop_16_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_16_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_16_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_16_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_16_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_16_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_16_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_16_is_fencei;	// rob.scala:310:28
  reg              rob_uop_16_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_16_uses_stq;	// rob.scala:310:28
  reg              rob_uop_16_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_16_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_16_ldst;	// rob.scala:310:28
  reg              rob_uop_16_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_16_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_16_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_17_uopc;	// rob.scala:310:28
  reg              rob_uop_17_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_17_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_17_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_17_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_17_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_17_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_17_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_17_is_fencei;	// rob.scala:310:28
  reg              rob_uop_17_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_17_uses_stq;	// rob.scala:310:28
  reg              rob_uop_17_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_17_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_17_ldst;	// rob.scala:310:28
  reg              rob_uop_17_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_17_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_17_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_18_uopc;	// rob.scala:310:28
  reg              rob_uop_18_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_18_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_18_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_18_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_18_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_18_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_18_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_18_is_fencei;	// rob.scala:310:28
  reg              rob_uop_18_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_18_uses_stq;	// rob.scala:310:28
  reg              rob_uop_18_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_18_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_18_ldst;	// rob.scala:310:28
  reg              rob_uop_18_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_18_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_18_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_19_uopc;	// rob.scala:310:28
  reg              rob_uop_19_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_19_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_19_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_19_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_19_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_19_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_19_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_19_is_fencei;	// rob.scala:310:28
  reg              rob_uop_19_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_19_uses_stq;	// rob.scala:310:28
  reg              rob_uop_19_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_19_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_19_ldst;	// rob.scala:310:28
  reg              rob_uop_19_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_19_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_19_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_20_uopc;	// rob.scala:310:28
  reg              rob_uop_20_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_20_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_20_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_20_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_20_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_20_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_20_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_20_is_fencei;	// rob.scala:310:28
  reg              rob_uop_20_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_20_uses_stq;	// rob.scala:310:28
  reg              rob_uop_20_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_20_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_20_ldst;	// rob.scala:310:28
  reg              rob_uop_20_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_20_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_20_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_21_uopc;	// rob.scala:310:28
  reg              rob_uop_21_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_21_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_21_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_21_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_21_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_21_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_21_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_21_is_fencei;	// rob.scala:310:28
  reg              rob_uop_21_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_21_uses_stq;	// rob.scala:310:28
  reg              rob_uop_21_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_21_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_21_ldst;	// rob.scala:310:28
  reg              rob_uop_21_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_21_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_21_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_22_uopc;	// rob.scala:310:28
  reg              rob_uop_22_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_22_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_22_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_22_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_22_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_22_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_22_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_22_is_fencei;	// rob.scala:310:28
  reg              rob_uop_22_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_22_uses_stq;	// rob.scala:310:28
  reg              rob_uop_22_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_22_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_22_ldst;	// rob.scala:310:28
  reg              rob_uop_22_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_22_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_22_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_23_uopc;	// rob.scala:310:28
  reg              rob_uop_23_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_23_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_23_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_23_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_23_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_23_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_23_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_23_is_fencei;	// rob.scala:310:28
  reg              rob_uop_23_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_23_uses_stq;	// rob.scala:310:28
  reg              rob_uop_23_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_23_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_23_ldst;	// rob.scala:310:28
  reg              rob_uop_23_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_23_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_23_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_24_uopc;	// rob.scala:310:28
  reg              rob_uop_24_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_24_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_24_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_24_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_24_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_24_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_24_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_24_is_fencei;	// rob.scala:310:28
  reg              rob_uop_24_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_24_uses_stq;	// rob.scala:310:28
  reg              rob_uop_24_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_24_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_24_ldst;	// rob.scala:310:28
  reg              rob_uop_24_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_24_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_24_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_25_uopc;	// rob.scala:310:28
  reg              rob_uop_25_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_25_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_25_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_25_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_25_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_25_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_25_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_25_is_fencei;	// rob.scala:310:28
  reg              rob_uop_25_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_25_uses_stq;	// rob.scala:310:28
  reg              rob_uop_25_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_25_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_25_ldst;	// rob.scala:310:28
  reg              rob_uop_25_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_25_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_25_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_26_uopc;	// rob.scala:310:28
  reg              rob_uop_26_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_26_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_26_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_26_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_26_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_26_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_26_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_26_is_fencei;	// rob.scala:310:28
  reg              rob_uop_26_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_26_uses_stq;	// rob.scala:310:28
  reg              rob_uop_26_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_26_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_26_ldst;	// rob.scala:310:28
  reg              rob_uop_26_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_26_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_26_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_27_uopc;	// rob.scala:310:28
  reg              rob_uop_27_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_27_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_27_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_27_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_27_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_27_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_27_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_27_is_fencei;	// rob.scala:310:28
  reg              rob_uop_27_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_27_uses_stq;	// rob.scala:310:28
  reg              rob_uop_27_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_27_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_27_ldst;	// rob.scala:310:28
  reg              rob_uop_27_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_27_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_27_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_28_uopc;	// rob.scala:310:28
  reg              rob_uop_28_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_28_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_28_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_28_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_28_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_28_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_28_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_28_is_fencei;	// rob.scala:310:28
  reg              rob_uop_28_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_28_uses_stq;	// rob.scala:310:28
  reg              rob_uop_28_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_28_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_28_ldst;	// rob.scala:310:28
  reg              rob_uop_28_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_28_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_28_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_29_uopc;	// rob.scala:310:28
  reg              rob_uop_29_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_29_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_29_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_29_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_29_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_29_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_29_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_29_is_fencei;	// rob.scala:310:28
  reg              rob_uop_29_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_29_uses_stq;	// rob.scala:310:28
  reg              rob_uop_29_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_29_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_29_ldst;	// rob.scala:310:28
  reg              rob_uop_29_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_29_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_29_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_30_uopc;	// rob.scala:310:28
  reg              rob_uop_30_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_30_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_30_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_30_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_30_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_30_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_30_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_30_is_fencei;	// rob.scala:310:28
  reg              rob_uop_30_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_30_uses_stq;	// rob.scala:310:28
  reg              rob_uop_30_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_30_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_30_ldst;	// rob.scala:310:28
  reg              rob_uop_30_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_30_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_30_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_31_uopc;	// rob.scala:310:28
  reg              rob_uop_31_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_31_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_31_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_31_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_31_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_31_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_31_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_31_is_fencei;	// rob.scala:310:28
  reg              rob_uop_31_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_31_uses_stq;	// rob.scala:310:28
  reg              rob_uop_31_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_31_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_31_ldst;	// rob.scala:310:28
  reg              rob_uop_31_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_31_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_31_fp_val;	// rob.scala:310:28
  reg              rob_exception_0;	// rob.scala:311:28
  reg              rob_exception_1;	// rob.scala:311:28
  reg              rob_exception_2;	// rob.scala:311:28
  reg              rob_exception_3;	// rob.scala:311:28
  reg              rob_exception_4;	// rob.scala:311:28
  reg              rob_exception_5;	// rob.scala:311:28
  reg              rob_exception_6;	// rob.scala:311:28
  reg              rob_exception_7;	// rob.scala:311:28
  reg              rob_exception_8;	// rob.scala:311:28
  reg              rob_exception_9;	// rob.scala:311:28
  reg              rob_exception_10;	// rob.scala:311:28
  reg              rob_exception_11;	// rob.scala:311:28
  reg              rob_exception_12;	// rob.scala:311:28
  reg              rob_exception_13;	// rob.scala:311:28
  reg              rob_exception_14;	// rob.scala:311:28
  reg              rob_exception_15;	// rob.scala:311:28
  reg              rob_exception_16;	// rob.scala:311:28
  reg              rob_exception_17;	// rob.scala:311:28
  reg              rob_exception_18;	// rob.scala:311:28
  reg              rob_exception_19;	// rob.scala:311:28
  reg              rob_exception_20;	// rob.scala:311:28
  reg              rob_exception_21;	// rob.scala:311:28
  reg              rob_exception_22;	// rob.scala:311:28
  reg              rob_exception_23;	// rob.scala:311:28
  reg              rob_exception_24;	// rob.scala:311:28
  reg              rob_exception_25;	// rob.scala:311:28
  reg              rob_exception_26;	// rob.scala:311:28
  reg              rob_exception_27;	// rob.scala:311:28
  reg              rob_exception_28;	// rob.scala:311:28
  reg              rob_exception_29;	// rob.scala:311:28
  reg              rob_exception_30;	// rob.scala:311:28
  reg              rob_exception_31;	// rob.scala:311:28
  reg              rob_predicated_0;	// rob.scala:312:29
  reg              rob_predicated_1;	// rob.scala:312:29
  reg              rob_predicated_2;	// rob.scala:312:29
  reg              rob_predicated_3;	// rob.scala:312:29
  reg              rob_predicated_4;	// rob.scala:312:29
  reg              rob_predicated_5;	// rob.scala:312:29
  reg              rob_predicated_6;	// rob.scala:312:29
  reg              rob_predicated_7;	// rob.scala:312:29
  reg              rob_predicated_8;	// rob.scala:312:29
  reg              rob_predicated_9;	// rob.scala:312:29
  reg              rob_predicated_10;	// rob.scala:312:29
  reg              rob_predicated_11;	// rob.scala:312:29
  reg              rob_predicated_12;	// rob.scala:312:29
  reg              rob_predicated_13;	// rob.scala:312:29
  reg              rob_predicated_14;	// rob.scala:312:29
  reg              rob_predicated_15;	// rob.scala:312:29
  reg              rob_predicated_16;	// rob.scala:312:29
  reg              rob_predicated_17;	// rob.scala:312:29
  reg              rob_predicated_18;	// rob.scala:312:29
  reg              rob_predicated_19;	// rob.scala:312:29
  reg              rob_predicated_20;	// rob.scala:312:29
  reg              rob_predicated_21;	// rob.scala:312:29
  reg              rob_predicated_22;	// rob.scala:312:29
  reg              rob_predicated_23;	// rob.scala:312:29
  reg              rob_predicated_24;	// rob.scala:312:29
  reg              rob_predicated_25;	// rob.scala:312:29
  reg              rob_predicated_26;	// rob.scala:312:29
  reg              rob_predicated_27;	// rob.scala:312:29
  reg              rob_predicated_28;	// rob.scala:312:29
  reg              rob_predicated_29;	// rob.scala:312:29
  reg              rob_predicated_30;	// rob.scala:312:29
  reg              rob_predicated_31;	// rob.scala:312:29
  wire [31:0]      _GEN =
    {{rob_val_31},
     {rob_val_30},
     {rob_val_29},
     {rob_val_28},
     {rob_val_27},
     {rob_val_26},
     {rob_val_25},
     {rob_val_24},
     {rob_val_23},
     {rob_val_22},
     {rob_val_21},
     {rob_val_20},
     {rob_val_19},
     {rob_val_18},
     {rob_val_17},
     {rob_val_16},
     {rob_val_15},
     {rob_val_14},
     {rob_val_13},
     {rob_val_12},
     {rob_val_11},
     {rob_val_10},
     {rob_val_9},
     {rob_val_8},
     {rob_val_7},
     {rob_val_6},
     {rob_val_5},
     {rob_val_4},
     {rob_val_3},
     {rob_val_2},
     {rob_val_1},
     {rob_val_0}};	// rob.scala:307:32, :324:31
  wire             rob_tail_vals_0 = _GEN[rob_tail];	// rob.scala:228:29, :324:31
  wire             _GEN_0 =
    io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_1 =
    io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_2 =
    io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_3 =
    io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_4 =
    io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_5 =
    io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_6 =
    io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_7 =
    io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_8 =
    io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_9 =
    io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_10 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :361:31
  wire [31:0]      _GEN_11 =
    {{rob_bsy_31},
     {rob_bsy_30},
     {rob_bsy_29},
     {rob_bsy_28},
     {rob_bsy_27},
     {rob_bsy_26},
     {rob_bsy_25},
     {rob_bsy_24},
     {rob_bsy_23},
     {rob_bsy_22},
     {rob_bsy_21},
     {rob_bsy_20},
     {rob_bsy_19},
     {rob_bsy_18},
     {rob_bsy_17},
     {rob_bsy_16},
     {rob_bsy_15},
     {rob_bsy_14},
     {rob_bsy_13},
     {rob_bsy_12},
     {rob_bsy_11},
     {rob_bsy_10},
     {rob_bsy_9},
     {rob_bsy_8},
     {rob_bsy_7},
     {rob_bsy_6},
     {rob_bsy_5},
     {rob_bsy_4},
     {rob_bsy_3},
     {rob_bsy_2},
     {rob_bsy_1},
     {rob_bsy_0}};	// rob.scala:308:28, :366:31
  wire             _GEN_12 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :361:31
  wire             _GEN_13 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :361:31
  wire             _GEN_14 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :390:26
  wire [31:0]      _GEN_15 =
    {{rob_unsafe_31},
     {rob_unsafe_30},
     {rob_unsafe_29},
     {rob_unsafe_28},
     {rob_unsafe_27},
     {rob_unsafe_26},
     {rob_unsafe_25},
     {rob_unsafe_24},
     {rob_unsafe_23},
     {rob_unsafe_22},
     {rob_unsafe_21},
     {rob_unsafe_20},
     {rob_unsafe_19},
     {rob_unsafe_18},
     {rob_unsafe_17},
     {rob_unsafe_16},
     {rob_unsafe_15},
     {rob_unsafe_14},
     {rob_unsafe_13},
     {rob_unsafe_12},
     {rob_unsafe_11},
     {rob_unsafe_10},
     {rob_unsafe_9},
     {rob_unsafe_8},
     {rob_unsafe_7},
     {rob_unsafe_6},
     {rob_unsafe_5},
     {rob_unsafe_4},
     {rob_unsafe_3},
     {rob_unsafe_2},
     {rob_unsafe_1},
     {rob_unsafe_0}};	// rob.scala:309:28, :394:15
  wire             rob_head_vals_0 = _GEN[rob_head];	// rob.scala:224:29, :324:31, :398:49
  wire [31:0]      _GEN_16 =
    {{rob_exception_31},
     {rob_exception_30},
     {rob_exception_29},
     {rob_exception_28},
     {rob_exception_27},
     {rob_exception_26},
     {rob_exception_25},
     {rob_exception_24},
     {rob_exception_23},
     {rob_exception_22},
     {rob_exception_21},
     {rob_exception_20},
     {rob_exception_19},
     {rob_exception_18},
     {rob_exception_17},
     {rob_exception_16},
     {rob_exception_15},
     {rob_exception_14},
     {rob_exception_13},
     {rob_exception_12},
     {rob_exception_11},
     {rob_exception_10},
     {rob_exception_9},
     {rob_exception_8},
     {rob_exception_7},
     {rob_exception_6},
     {rob_exception_5},
     {rob_exception_4},
     {rob_exception_3},
     {rob_exception_2},
     {rob_exception_1},
     {rob_exception_0}};	// rob.scala:311:28, :398:49
  wire             can_throw_exception_0 = rob_head_vals_0 & _GEN_16[rob_head];	// rob.scala:224:29, :398:49
  wire             can_commit_0 = rob_head_vals_0 & ~_GEN_11[rob_head] & ~io_csr_stall;	// rob.scala:224:29, :366:31, :398:49, :404:{43,64,67}
  wire [31:0]      _GEN_17 =
    {{rob_predicated_31},
     {rob_predicated_30},
     {rob_predicated_29},
     {rob_predicated_28},
     {rob_predicated_27},
     {rob_predicated_26},
     {rob_predicated_25},
     {rob_predicated_24},
     {rob_predicated_23},
     {rob_predicated_22},
     {rob_predicated_21},
     {rob_predicated_20},
     {rob_predicated_19},
     {rob_predicated_18},
     {rob_predicated_17},
     {rob_predicated_16},
     {rob_predicated_15},
     {rob_predicated_14},
     {rob_predicated_13},
     {rob_predicated_12},
     {rob_predicated_11},
     {rob_predicated_10},
     {rob_predicated_9},
     {rob_predicated_8},
     {rob_predicated_7},
     {rob_predicated_6},
     {rob_predicated_5},
     {rob_predicated_4},
     {rob_predicated_3},
     {rob_predicated_2},
     {rob_predicated_1},
     {rob_predicated_0}};	// rob.scala:312:29, :410:51
  wire [31:0][6:0] _GEN_18 =
    {{rob_uop_31_uopc},
     {rob_uop_30_uopc},
     {rob_uop_29_uopc},
     {rob_uop_28_uopc},
     {rob_uop_27_uopc},
     {rob_uop_26_uopc},
     {rob_uop_25_uopc},
     {rob_uop_24_uopc},
     {rob_uop_23_uopc},
     {rob_uop_22_uopc},
     {rob_uop_21_uopc},
     {rob_uop_20_uopc},
     {rob_uop_19_uopc},
     {rob_uop_18_uopc},
     {rob_uop_17_uopc},
     {rob_uop_16_uopc},
     {rob_uop_15_uopc},
     {rob_uop_14_uopc},
     {rob_uop_13_uopc},
     {rob_uop_12_uopc},
     {rob_uop_11_uopc},
     {rob_uop_10_uopc},
     {rob_uop_9_uopc},
     {rob_uop_8_uopc},
     {rob_uop_7_uopc},
     {rob_uop_6_uopc},
     {rob_uop_5_uopc},
     {rob_uop_4_uopc},
     {rob_uop_3_uopc},
     {rob_uop_2_uopc},
     {rob_uop_1_uopc},
     {rob_uop_0_uopc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_19 =
    {{rob_uop_31_is_rvc},
     {rob_uop_30_is_rvc},
     {rob_uop_29_is_rvc},
     {rob_uop_28_is_rvc},
     {rob_uop_27_is_rvc},
     {rob_uop_26_is_rvc},
     {rob_uop_25_is_rvc},
     {rob_uop_24_is_rvc},
     {rob_uop_23_is_rvc},
     {rob_uop_22_is_rvc},
     {rob_uop_21_is_rvc},
     {rob_uop_20_is_rvc},
     {rob_uop_19_is_rvc},
     {rob_uop_18_is_rvc},
     {rob_uop_17_is_rvc},
     {rob_uop_16_is_rvc},
     {rob_uop_15_is_rvc},
     {rob_uop_14_is_rvc},
     {rob_uop_13_is_rvc},
     {rob_uop_12_is_rvc},
     {rob_uop_11_is_rvc},
     {rob_uop_10_is_rvc},
     {rob_uop_9_is_rvc},
     {rob_uop_8_is_rvc},
     {rob_uop_7_is_rvc},
     {rob_uop_6_is_rvc},
     {rob_uop_5_is_rvc},
     {rob_uop_4_is_rvc},
     {rob_uop_3_is_rvc},
     {rob_uop_2_is_rvc},
     {rob_uop_1_is_rvc},
     {rob_uop_0_is_rvc}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_20 =
    {{rob_uop_31_ftq_idx},
     {rob_uop_30_ftq_idx},
     {rob_uop_29_ftq_idx},
     {rob_uop_28_ftq_idx},
     {rob_uop_27_ftq_idx},
     {rob_uop_26_ftq_idx},
     {rob_uop_25_ftq_idx},
     {rob_uop_24_ftq_idx},
     {rob_uop_23_ftq_idx},
     {rob_uop_22_ftq_idx},
     {rob_uop_21_ftq_idx},
     {rob_uop_20_ftq_idx},
     {rob_uop_19_ftq_idx},
     {rob_uop_18_ftq_idx},
     {rob_uop_17_ftq_idx},
     {rob_uop_16_ftq_idx},
     {rob_uop_15_ftq_idx},
     {rob_uop_14_ftq_idx},
     {rob_uop_13_ftq_idx},
     {rob_uop_12_ftq_idx},
     {rob_uop_11_ftq_idx},
     {rob_uop_10_ftq_idx},
     {rob_uop_9_ftq_idx},
     {rob_uop_8_ftq_idx},
     {rob_uop_7_ftq_idx},
     {rob_uop_6_ftq_idx},
     {rob_uop_5_ftq_idx},
     {rob_uop_4_ftq_idx},
     {rob_uop_3_ftq_idx},
     {rob_uop_2_ftq_idx},
     {rob_uop_1_ftq_idx},
     {rob_uop_0_ftq_idx}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_21 =
    {{rob_uop_31_edge_inst},
     {rob_uop_30_edge_inst},
     {rob_uop_29_edge_inst},
     {rob_uop_28_edge_inst},
     {rob_uop_27_edge_inst},
     {rob_uop_26_edge_inst},
     {rob_uop_25_edge_inst},
     {rob_uop_24_edge_inst},
     {rob_uop_23_edge_inst},
     {rob_uop_22_edge_inst},
     {rob_uop_21_edge_inst},
     {rob_uop_20_edge_inst},
     {rob_uop_19_edge_inst},
     {rob_uop_18_edge_inst},
     {rob_uop_17_edge_inst},
     {rob_uop_16_edge_inst},
     {rob_uop_15_edge_inst},
     {rob_uop_14_edge_inst},
     {rob_uop_13_edge_inst},
     {rob_uop_12_edge_inst},
     {rob_uop_11_edge_inst},
     {rob_uop_10_edge_inst},
     {rob_uop_9_edge_inst},
     {rob_uop_8_edge_inst},
     {rob_uop_7_edge_inst},
     {rob_uop_6_edge_inst},
     {rob_uop_5_edge_inst},
     {rob_uop_4_edge_inst},
     {rob_uop_3_edge_inst},
     {rob_uop_2_edge_inst},
     {rob_uop_1_edge_inst},
     {rob_uop_0_edge_inst}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_22 =
    {{rob_uop_31_pc_lob},
     {rob_uop_30_pc_lob},
     {rob_uop_29_pc_lob},
     {rob_uop_28_pc_lob},
     {rob_uop_27_pc_lob},
     {rob_uop_26_pc_lob},
     {rob_uop_25_pc_lob},
     {rob_uop_24_pc_lob},
     {rob_uop_23_pc_lob},
     {rob_uop_22_pc_lob},
     {rob_uop_21_pc_lob},
     {rob_uop_20_pc_lob},
     {rob_uop_19_pc_lob},
     {rob_uop_18_pc_lob},
     {rob_uop_17_pc_lob},
     {rob_uop_16_pc_lob},
     {rob_uop_15_pc_lob},
     {rob_uop_14_pc_lob},
     {rob_uop_13_pc_lob},
     {rob_uop_12_pc_lob},
     {rob_uop_11_pc_lob},
     {rob_uop_10_pc_lob},
     {rob_uop_9_pc_lob},
     {rob_uop_8_pc_lob},
     {rob_uop_7_pc_lob},
     {rob_uop_6_pc_lob},
     {rob_uop_5_pc_lob},
     {rob_uop_4_pc_lob},
     {rob_uop_3_pc_lob},
     {rob_uop_2_pc_lob},
     {rob_uop_1_pc_lob},
     {rob_uop_0_pc_lob}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_23 =
    {{rob_uop_31_pdst},
     {rob_uop_30_pdst},
     {rob_uop_29_pdst},
     {rob_uop_28_pdst},
     {rob_uop_27_pdst},
     {rob_uop_26_pdst},
     {rob_uop_25_pdst},
     {rob_uop_24_pdst},
     {rob_uop_23_pdst},
     {rob_uop_22_pdst},
     {rob_uop_21_pdst},
     {rob_uop_20_pdst},
     {rob_uop_19_pdst},
     {rob_uop_18_pdst},
     {rob_uop_17_pdst},
     {rob_uop_16_pdst},
     {rob_uop_15_pdst},
     {rob_uop_14_pdst},
     {rob_uop_13_pdst},
     {rob_uop_12_pdst},
     {rob_uop_11_pdst},
     {rob_uop_10_pdst},
     {rob_uop_9_pdst},
     {rob_uop_8_pdst},
     {rob_uop_7_pdst},
     {rob_uop_6_pdst},
     {rob_uop_5_pdst},
     {rob_uop_4_pdst},
     {rob_uop_3_pdst},
     {rob_uop_2_pdst},
     {rob_uop_1_pdst},
     {rob_uop_0_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_24 =
    {{rob_uop_31_stale_pdst},
     {rob_uop_30_stale_pdst},
     {rob_uop_29_stale_pdst},
     {rob_uop_28_stale_pdst},
     {rob_uop_27_stale_pdst},
     {rob_uop_26_stale_pdst},
     {rob_uop_25_stale_pdst},
     {rob_uop_24_stale_pdst},
     {rob_uop_23_stale_pdst},
     {rob_uop_22_stale_pdst},
     {rob_uop_21_stale_pdst},
     {rob_uop_20_stale_pdst},
     {rob_uop_19_stale_pdst},
     {rob_uop_18_stale_pdst},
     {rob_uop_17_stale_pdst},
     {rob_uop_16_stale_pdst},
     {rob_uop_15_stale_pdst},
     {rob_uop_14_stale_pdst},
     {rob_uop_13_stale_pdst},
     {rob_uop_12_stale_pdst},
     {rob_uop_11_stale_pdst},
     {rob_uop_10_stale_pdst},
     {rob_uop_9_stale_pdst},
     {rob_uop_8_stale_pdst},
     {rob_uop_7_stale_pdst},
     {rob_uop_6_stale_pdst},
     {rob_uop_5_stale_pdst},
     {rob_uop_4_stale_pdst},
     {rob_uop_3_stale_pdst},
     {rob_uop_2_stale_pdst},
     {rob_uop_1_stale_pdst},
     {rob_uop_0_stale_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_25 =
    {{rob_uop_31_is_fencei},
     {rob_uop_30_is_fencei},
     {rob_uop_29_is_fencei},
     {rob_uop_28_is_fencei},
     {rob_uop_27_is_fencei},
     {rob_uop_26_is_fencei},
     {rob_uop_25_is_fencei},
     {rob_uop_24_is_fencei},
     {rob_uop_23_is_fencei},
     {rob_uop_22_is_fencei},
     {rob_uop_21_is_fencei},
     {rob_uop_20_is_fencei},
     {rob_uop_19_is_fencei},
     {rob_uop_18_is_fencei},
     {rob_uop_17_is_fencei},
     {rob_uop_16_is_fencei},
     {rob_uop_15_is_fencei},
     {rob_uop_14_is_fencei},
     {rob_uop_13_is_fencei},
     {rob_uop_12_is_fencei},
     {rob_uop_11_is_fencei},
     {rob_uop_10_is_fencei},
     {rob_uop_9_is_fencei},
     {rob_uop_8_is_fencei},
     {rob_uop_7_is_fencei},
     {rob_uop_6_is_fencei},
     {rob_uop_5_is_fencei},
     {rob_uop_4_is_fencei},
     {rob_uop_3_is_fencei},
     {rob_uop_2_is_fencei},
     {rob_uop_1_is_fencei},
     {rob_uop_0_is_fencei}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_26 =
    {{rob_uop_31_uses_ldq},
     {rob_uop_30_uses_ldq},
     {rob_uop_29_uses_ldq},
     {rob_uop_28_uses_ldq},
     {rob_uop_27_uses_ldq},
     {rob_uop_26_uses_ldq},
     {rob_uop_25_uses_ldq},
     {rob_uop_24_uses_ldq},
     {rob_uop_23_uses_ldq},
     {rob_uop_22_uses_ldq},
     {rob_uop_21_uses_ldq},
     {rob_uop_20_uses_ldq},
     {rob_uop_19_uses_ldq},
     {rob_uop_18_uses_ldq},
     {rob_uop_17_uses_ldq},
     {rob_uop_16_uses_ldq},
     {rob_uop_15_uses_ldq},
     {rob_uop_14_uses_ldq},
     {rob_uop_13_uses_ldq},
     {rob_uop_12_uses_ldq},
     {rob_uop_11_uses_ldq},
     {rob_uop_10_uses_ldq},
     {rob_uop_9_uses_ldq},
     {rob_uop_8_uses_ldq},
     {rob_uop_7_uses_ldq},
     {rob_uop_6_uses_ldq},
     {rob_uop_5_uses_ldq},
     {rob_uop_4_uses_ldq},
     {rob_uop_3_uses_ldq},
     {rob_uop_2_uses_ldq},
     {rob_uop_1_uses_ldq},
     {rob_uop_0_uses_ldq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_27 =
    {{rob_uop_31_uses_stq},
     {rob_uop_30_uses_stq},
     {rob_uop_29_uses_stq},
     {rob_uop_28_uses_stq},
     {rob_uop_27_uses_stq},
     {rob_uop_26_uses_stq},
     {rob_uop_25_uses_stq},
     {rob_uop_24_uses_stq},
     {rob_uop_23_uses_stq},
     {rob_uop_22_uses_stq},
     {rob_uop_21_uses_stq},
     {rob_uop_20_uses_stq},
     {rob_uop_19_uses_stq},
     {rob_uop_18_uses_stq},
     {rob_uop_17_uses_stq},
     {rob_uop_16_uses_stq},
     {rob_uop_15_uses_stq},
     {rob_uop_14_uses_stq},
     {rob_uop_13_uses_stq},
     {rob_uop_12_uses_stq},
     {rob_uop_11_uses_stq},
     {rob_uop_10_uses_stq},
     {rob_uop_9_uses_stq},
     {rob_uop_8_uses_stq},
     {rob_uop_7_uses_stq},
     {rob_uop_6_uses_stq},
     {rob_uop_5_uses_stq},
     {rob_uop_4_uses_stq},
     {rob_uop_3_uses_stq},
     {rob_uop_2_uses_stq},
     {rob_uop_1_uses_stq},
     {rob_uop_0_uses_stq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_28 =
    {{rob_uop_31_is_sys_pc2epc},
     {rob_uop_30_is_sys_pc2epc},
     {rob_uop_29_is_sys_pc2epc},
     {rob_uop_28_is_sys_pc2epc},
     {rob_uop_27_is_sys_pc2epc},
     {rob_uop_26_is_sys_pc2epc},
     {rob_uop_25_is_sys_pc2epc},
     {rob_uop_24_is_sys_pc2epc},
     {rob_uop_23_is_sys_pc2epc},
     {rob_uop_22_is_sys_pc2epc},
     {rob_uop_21_is_sys_pc2epc},
     {rob_uop_20_is_sys_pc2epc},
     {rob_uop_19_is_sys_pc2epc},
     {rob_uop_18_is_sys_pc2epc},
     {rob_uop_17_is_sys_pc2epc},
     {rob_uop_16_is_sys_pc2epc},
     {rob_uop_15_is_sys_pc2epc},
     {rob_uop_14_is_sys_pc2epc},
     {rob_uop_13_is_sys_pc2epc},
     {rob_uop_12_is_sys_pc2epc},
     {rob_uop_11_is_sys_pc2epc},
     {rob_uop_10_is_sys_pc2epc},
     {rob_uop_9_is_sys_pc2epc},
     {rob_uop_8_is_sys_pc2epc},
     {rob_uop_7_is_sys_pc2epc},
     {rob_uop_6_is_sys_pc2epc},
     {rob_uop_5_is_sys_pc2epc},
     {rob_uop_4_is_sys_pc2epc},
     {rob_uop_3_is_sys_pc2epc},
     {rob_uop_2_is_sys_pc2epc},
     {rob_uop_1_is_sys_pc2epc},
     {rob_uop_0_is_sys_pc2epc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_29 =
    {{rob_uop_31_flush_on_commit},
     {rob_uop_30_flush_on_commit},
     {rob_uop_29_flush_on_commit},
     {rob_uop_28_flush_on_commit},
     {rob_uop_27_flush_on_commit},
     {rob_uop_26_flush_on_commit},
     {rob_uop_25_flush_on_commit},
     {rob_uop_24_flush_on_commit},
     {rob_uop_23_flush_on_commit},
     {rob_uop_22_flush_on_commit},
     {rob_uop_21_flush_on_commit},
     {rob_uop_20_flush_on_commit},
     {rob_uop_19_flush_on_commit},
     {rob_uop_18_flush_on_commit},
     {rob_uop_17_flush_on_commit},
     {rob_uop_16_flush_on_commit},
     {rob_uop_15_flush_on_commit},
     {rob_uop_14_flush_on_commit},
     {rob_uop_13_flush_on_commit},
     {rob_uop_12_flush_on_commit},
     {rob_uop_11_flush_on_commit},
     {rob_uop_10_flush_on_commit},
     {rob_uop_9_flush_on_commit},
     {rob_uop_8_flush_on_commit},
     {rob_uop_7_flush_on_commit},
     {rob_uop_6_flush_on_commit},
     {rob_uop_5_flush_on_commit},
     {rob_uop_4_flush_on_commit},
     {rob_uop_3_flush_on_commit},
     {rob_uop_2_flush_on_commit},
     {rob_uop_1_flush_on_commit},
     {rob_uop_0_flush_on_commit}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_30 =
    {{rob_uop_31_ldst},
     {rob_uop_30_ldst},
     {rob_uop_29_ldst},
     {rob_uop_28_ldst},
     {rob_uop_27_ldst},
     {rob_uop_26_ldst},
     {rob_uop_25_ldst},
     {rob_uop_24_ldst},
     {rob_uop_23_ldst},
     {rob_uop_22_ldst},
     {rob_uop_21_ldst},
     {rob_uop_20_ldst},
     {rob_uop_19_ldst},
     {rob_uop_18_ldst},
     {rob_uop_17_ldst},
     {rob_uop_16_ldst},
     {rob_uop_15_ldst},
     {rob_uop_14_ldst},
     {rob_uop_13_ldst},
     {rob_uop_12_ldst},
     {rob_uop_11_ldst},
     {rob_uop_10_ldst},
     {rob_uop_9_ldst},
     {rob_uop_8_ldst},
     {rob_uop_7_ldst},
     {rob_uop_6_ldst},
     {rob_uop_5_ldst},
     {rob_uop_4_ldst},
     {rob_uop_3_ldst},
     {rob_uop_2_ldst},
     {rob_uop_1_ldst},
     {rob_uop_0_ldst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_31 =
    {{rob_uop_31_ldst_val},
     {rob_uop_30_ldst_val},
     {rob_uop_29_ldst_val},
     {rob_uop_28_ldst_val},
     {rob_uop_27_ldst_val},
     {rob_uop_26_ldst_val},
     {rob_uop_25_ldst_val},
     {rob_uop_24_ldst_val},
     {rob_uop_23_ldst_val},
     {rob_uop_22_ldst_val},
     {rob_uop_21_ldst_val},
     {rob_uop_20_ldst_val},
     {rob_uop_19_ldst_val},
     {rob_uop_18_ldst_val},
     {rob_uop_17_ldst_val},
     {rob_uop_16_ldst_val},
     {rob_uop_15_ldst_val},
     {rob_uop_14_ldst_val},
     {rob_uop_13_ldst_val},
     {rob_uop_12_ldst_val},
     {rob_uop_11_ldst_val},
     {rob_uop_10_ldst_val},
     {rob_uop_9_ldst_val},
     {rob_uop_8_ldst_val},
     {rob_uop_7_ldst_val},
     {rob_uop_6_ldst_val},
     {rob_uop_5_ldst_val},
     {rob_uop_4_ldst_val},
     {rob_uop_3_ldst_val},
     {rob_uop_2_ldst_val},
     {rob_uop_1_ldst_val},
     {rob_uop_0_ldst_val}};	// rob.scala:310:28, :411:25
  wire [31:0][1:0] _GEN_32 =
    {{rob_uop_31_dst_rtype},
     {rob_uop_30_dst_rtype},
     {rob_uop_29_dst_rtype},
     {rob_uop_28_dst_rtype},
     {rob_uop_27_dst_rtype},
     {rob_uop_26_dst_rtype},
     {rob_uop_25_dst_rtype},
     {rob_uop_24_dst_rtype},
     {rob_uop_23_dst_rtype},
     {rob_uop_22_dst_rtype},
     {rob_uop_21_dst_rtype},
     {rob_uop_20_dst_rtype},
     {rob_uop_19_dst_rtype},
     {rob_uop_18_dst_rtype},
     {rob_uop_17_dst_rtype},
     {rob_uop_16_dst_rtype},
     {rob_uop_15_dst_rtype},
     {rob_uop_14_dst_rtype},
     {rob_uop_13_dst_rtype},
     {rob_uop_12_dst_rtype},
     {rob_uop_11_dst_rtype},
     {rob_uop_10_dst_rtype},
     {rob_uop_9_dst_rtype},
     {rob_uop_8_dst_rtype},
     {rob_uop_7_dst_rtype},
     {rob_uop_6_dst_rtype},
     {rob_uop_5_dst_rtype},
     {rob_uop_4_dst_rtype},
     {rob_uop_3_dst_rtype},
     {rob_uop_2_dst_rtype},
     {rob_uop_1_dst_rtype},
     {rob_uop_0_dst_rtype}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_33 =
    {{rob_uop_31_fp_val},
     {rob_uop_30_fp_val},
     {rob_uop_29_fp_val},
     {rob_uop_28_fp_val},
     {rob_uop_27_fp_val},
     {rob_uop_26_fp_val},
     {rob_uop_25_fp_val},
     {rob_uop_24_fp_val},
     {rob_uop_23_fp_val},
     {rob_uop_22_fp_val},
     {rob_uop_21_fp_val},
     {rob_uop_20_fp_val},
     {rob_uop_19_fp_val},
     {rob_uop_18_fp_val},
     {rob_uop_17_fp_val},
     {rob_uop_16_fp_val},
     {rob_uop_15_fp_val},
     {rob_uop_14_fp_val},
     {rob_uop_13_fp_val},
     {rob_uop_12_fp_val},
     {rob_uop_11_fp_val},
     {rob_uop_10_fp_val},
     {rob_uop_9_fp_val},
     {rob_uop_8_fp_val},
     {rob_uop_7_fp_val},
     {rob_uop_6_fp_val},
     {rob_uop_5_fp_val},
     {rob_uop_4_fp_val},
     {rob_uop_3_fp_val},
     {rob_uop_2_fp_val},
     {rob_uop_1_fp_val},
     {rob_uop_0_fp_val}};	// rob.scala:310:28, :411:25
  wire             rbk_row = _io_commit_rollback_T_3 & ~full;	// rob.scala:236:31, :425:{44,47}, :787:39
  wire             _io_commit_rbk_valids_0_output = rbk_row & _GEN[com_idx];	// rob.scala:236:20, :324:31, :425:44, :427:40
  reg              rob_val_1_0;	// rob.scala:307:32
  reg              rob_val_1_1;	// rob.scala:307:32
  reg              rob_val_1_2;	// rob.scala:307:32
  reg              rob_val_1_3;	// rob.scala:307:32
  reg              rob_val_1_4;	// rob.scala:307:32
  reg              rob_val_1_5;	// rob.scala:307:32
  reg              rob_val_1_6;	// rob.scala:307:32
  reg              rob_val_1_7;	// rob.scala:307:32
  reg              rob_val_1_8;	// rob.scala:307:32
  reg              rob_val_1_9;	// rob.scala:307:32
  reg              rob_val_1_10;	// rob.scala:307:32
  reg              rob_val_1_11;	// rob.scala:307:32
  reg              rob_val_1_12;	// rob.scala:307:32
  reg              rob_val_1_13;	// rob.scala:307:32
  reg              rob_val_1_14;	// rob.scala:307:32
  reg              rob_val_1_15;	// rob.scala:307:32
  reg              rob_val_1_16;	// rob.scala:307:32
  reg              rob_val_1_17;	// rob.scala:307:32
  reg              rob_val_1_18;	// rob.scala:307:32
  reg              rob_val_1_19;	// rob.scala:307:32
  reg              rob_val_1_20;	// rob.scala:307:32
  reg              rob_val_1_21;	// rob.scala:307:32
  reg              rob_val_1_22;	// rob.scala:307:32
  reg              rob_val_1_23;	// rob.scala:307:32
  reg              rob_val_1_24;	// rob.scala:307:32
  reg              rob_val_1_25;	// rob.scala:307:32
  reg              rob_val_1_26;	// rob.scala:307:32
  reg              rob_val_1_27;	// rob.scala:307:32
  reg              rob_val_1_28;	// rob.scala:307:32
  reg              rob_val_1_29;	// rob.scala:307:32
  reg              rob_val_1_30;	// rob.scala:307:32
  reg              rob_val_1_31;	// rob.scala:307:32
  reg              rob_bsy_1_0;	// rob.scala:308:28
  reg              rob_bsy_1_1;	// rob.scala:308:28
  reg              rob_bsy_1_2;	// rob.scala:308:28
  reg              rob_bsy_1_3;	// rob.scala:308:28
  reg              rob_bsy_1_4;	// rob.scala:308:28
  reg              rob_bsy_1_5;	// rob.scala:308:28
  reg              rob_bsy_1_6;	// rob.scala:308:28
  reg              rob_bsy_1_7;	// rob.scala:308:28
  reg              rob_bsy_1_8;	// rob.scala:308:28
  reg              rob_bsy_1_9;	// rob.scala:308:28
  reg              rob_bsy_1_10;	// rob.scala:308:28
  reg              rob_bsy_1_11;	// rob.scala:308:28
  reg              rob_bsy_1_12;	// rob.scala:308:28
  reg              rob_bsy_1_13;	// rob.scala:308:28
  reg              rob_bsy_1_14;	// rob.scala:308:28
  reg              rob_bsy_1_15;	// rob.scala:308:28
  reg              rob_bsy_1_16;	// rob.scala:308:28
  reg              rob_bsy_1_17;	// rob.scala:308:28
  reg              rob_bsy_1_18;	// rob.scala:308:28
  reg              rob_bsy_1_19;	// rob.scala:308:28
  reg              rob_bsy_1_20;	// rob.scala:308:28
  reg              rob_bsy_1_21;	// rob.scala:308:28
  reg              rob_bsy_1_22;	// rob.scala:308:28
  reg              rob_bsy_1_23;	// rob.scala:308:28
  reg              rob_bsy_1_24;	// rob.scala:308:28
  reg              rob_bsy_1_25;	// rob.scala:308:28
  reg              rob_bsy_1_26;	// rob.scala:308:28
  reg              rob_bsy_1_27;	// rob.scala:308:28
  reg              rob_bsy_1_28;	// rob.scala:308:28
  reg              rob_bsy_1_29;	// rob.scala:308:28
  reg              rob_bsy_1_30;	// rob.scala:308:28
  reg              rob_bsy_1_31;	// rob.scala:308:28
  reg              rob_unsafe_1_0;	// rob.scala:309:28
  reg              rob_unsafe_1_1;	// rob.scala:309:28
  reg              rob_unsafe_1_2;	// rob.scala:309:28
  reg              rob_unsafe_1_3;	// rob.scala:309:28
  reg              rob_unsafe_1_4;	// rob.scala:309:28
  reg              rob_unsafe_1_5;	// rob.scala:309:28
  reg              rob_unsafe_1_6;	// rob.scala:309:28
  reg              rob_unsafe_1_7;	// rob.scala:309:28
  reg              rob_unsafe_1_8;	// rob.scala:309:28
  reg              rob_unsafe_1_9;	// rob.scala:309:28
  reg              rob_unsafe_1_10;	// rob.scala:309:28
  reg              rob_unsafe_1_11;	// rob.scala:309:28
  reg              rob_unsafe_1_12;	// rob.scala:309:28
  reg              rob_unsafe_1_13;	// rob.scala:309:28
  reg              rob_unsafe_1_14;	// rob.scala:309:28
  reg              rob_unsafe_1_15;	// rob.scala:309:28
  reg              rob_unsafe_1_16;	// rob.scala:309:28
  reg              rob_unsafe_1_17;	// rob.scala:309:28
  reg              rob_unsafe_1_18;	// rob.scala:309:28
  reg              rob_unsafe_1_19;	// rob.scala:309:28
  reg              rob_unsafe_1_20;	// rob.scala:309:28
  reg              rob_unsafe_1_21;	// rob.scala:309:28
  reg              rob_unsafe_1_22;	// rob.scala:309:28
  reg              rob_unsafe_1_23;	// rob.scala:309:28
  reg              rob_unsafe_1_24;	// rob.scala:309:28
  reg              rob_unsafe_1_25;	// rob.scala:309:28
  reg              rob_unsafe_1_26;	// rob.scala:309:28
  reg              rob_unsafe_1_27;	// rob.scala:309:28
  reg              rob_unsafe_1_28;	// rob.scala:309:28
  reg              rob_unsafe_1_29;	// rob.scala:309:28
  reg              rob_unsafe_1_30;	// rob.scala:309:28
  reg              rob_unsafe_1_31;	// rob.scala:309:28
  reg  [6:0]       rob_uop_1_0_uopc;	// rob.scala:310:28
  reg              rob_uop_1_0_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_0_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_0_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_0_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_0_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_0_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_0_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_0_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_0_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_0_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_0_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_0_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_0_ldst;	// rob.scala:310:28
  reg              rob_uop_1_0_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_0_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_0_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_1_uopc;	// rob.scala:310:28
  reg              rob_uop_1_1_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_1_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_1_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_1_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_1_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_1_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_1_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_1_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_1_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_1_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_1_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_1_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_1_ldst;	// rob.scala:310:28
  reg              rob_uop_1_1_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_1_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_1_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_2_uopc;	// rob.scala:310:28
  reg              rob_uop_1_2_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_2_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_2_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_2_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_2_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_2_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_2_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_2_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_2_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_2_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_2_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_2_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_2_ldst;	// rob.scala:310:28
  reg              rob_uop_1_2_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_2_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_2_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_3_uopc;	// rob.scala:310:28
  reg              rob_uop_1_3_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_3_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_3_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_3_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_3_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_3_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_3_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_3_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_3_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_3_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_3_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_3_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_3_ldst;	// rob.scala:310:28
  reg              rob_uop_1_3_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_3_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_3_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_4_uopc;	// rob.scala:310:28
  reg              rob_uop_1_4_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_4_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_4_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_4_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_4_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_4_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_4_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_4_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_4_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_4_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_4_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_4_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_4_ldst;	// rob.scala:310:28
  reg              rob_uop_1_4_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_4_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_4_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_5_uopc;	// rob.scala:310:28
  reg              rob_uop_1_5_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_5_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_5_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_5_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_5_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_5_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_5_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_5_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_5_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_5_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_5_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_5_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_5_ldst;	// rob.scala:310:28
  reg              rob_uop_1_5_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_5_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_5_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_6_uopc;	// rob.scala:310:28
  reg              rob_uop_1_6_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_6_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_6_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_6_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_6_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_6_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_6_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_6_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_6_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_6_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_6_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_6_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_6_ldst;	// rob.scala:310:28
  reg              rob_uop_1_6_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_6_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_6_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_7_uopc;	// rob.scala:310:28
  reg              rob_uop_1_7_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_7_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_7_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_7_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_7_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_7_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_7_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_7_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_7_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_7_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_7_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_7_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_7_ldst;	// rob.scala:310:28
  reg              rob_uop_1_7_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_7_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_7_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_8_uopc;	// rob.scala:310:28
  reg              rob_uop_1_8_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_8_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_8_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_8_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_8_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_8_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_8_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_8_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_8_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_8_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_8_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_8_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_8_ldst;	// rob.scala:310:28
  reg              rob_uop_1_8_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_8_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_8_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_9_uopc;	// rob.scala:310:28
  reg              rob_uop_1_9_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_9_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_9_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_9_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_9_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_9_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_9_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_9_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_9_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_9_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_9_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_9_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_9_ldst;	// rob.scala:310:28
  reg              rob_uop_1_9_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_9_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_9_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_10_uopc;	// rob.scala:310:28
  reg              rob_uop_1_10_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_10_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_10_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_10_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_10_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_10_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_10_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_10_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_10_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_10_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_10_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_10_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_10_ldst;	// rob.scala:310:28
  reg              rob_uop_1_10_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_10_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_10_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_11_uopc;	// rob.scala:310:28
  reg              rob_uop_1_11_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_11_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_11_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_11_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_11_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_11_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_11_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_11_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_11_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_11_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_11_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_11_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_11_ldst;	// rob.scala:310:28
  reg              rob_uop_1_11_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_11_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_11_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_12_uopc;	// rob.scala:310:28
  reg              rob_uop_1_12_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_12_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_12_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_12_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_12_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_12_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_12_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_12_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_12_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_12_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_12_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_12_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_12_ldst;	// rob.scala:310:28
  reg              rob_uop_1_12_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_12_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_12_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_13_uopc;	// rob.scala:310:28
  reg              rob_uop_1_13_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_13_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_13_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_13_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_13_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_13_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_13_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_13_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_13_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_13_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_13_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_13_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_13_ldst;	// rob.scala:310:28
  reg              rob_uop_1_13_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_13_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_13_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_14_uopc;	// rob.scala:310:28
  reg              rob_uop_1_14_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_14_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_14_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_14_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_14_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_14_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_14_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_14_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_14_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_14_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_14_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_14_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_14_ldst;	// rob.scala:310:28
  reg              rob_uop_1_14_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_14_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_14_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_15_uopc;	// rob.scala:310:28
  reg              rob_uop_1_15_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_15_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_15_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_15_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_15_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_15_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_15_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_15_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_15_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_15_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_15_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_15_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_15_ldst;	// rob.scala:310:28
  reg              rob_uop_1_15_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_15_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_15_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_16_uopc;	// rob.scala:310:28
  reg              rob_uop_1_16_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_16_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_16_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_16_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_16_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_16_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_16_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_16_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_16_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_16_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_16_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_16_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_16_ldst;	// rob.scala:310:28
  reg              rob_uop_1_16_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_16_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_16_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_17_uopc;	// rob.scala:310:28
  reg              rob_uop_1_17_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_17_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_17_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_17_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_17_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_17_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_17_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_17_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_17_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_17_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_17_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_17_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_17_ldst;	// rob.scala:310:28
  reg              rob_uop_1_17_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_17_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_17_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_18_uopc;	// rob.scala:310:28
  reg              rob_uop_1_18_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_18_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_18_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_18_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_18_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_18_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_18_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_18_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_18_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_18_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_18_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_18_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_18_ldst;	// rob.scala:310:28
  reg              rob_uop_1_18_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_18_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_18_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_19_uopc;	// rob.scala:310:28
  reg              rob_uop_1_19_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_19_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_19_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_19_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_19_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_19_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_19_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_19_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_19_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_19_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_19_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_19_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_19_ldst;	// rob.scala:310:28
  reg              rob_uop_1_19_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_19_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_19_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_20_uopc;	// rob.scala:310:28
  reg              rob_uop_1_20_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_20_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_20_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_20_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_20_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_20_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_20_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_20_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_20_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_20_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_20_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_20_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_20_ldst;	// rob.scala:310:28
  reg              rob_uop_1_20_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_20_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_20_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_21_uopc;	// rob.scala:310:28
  reg              rob_uop_1_21_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_21_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_21_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_21_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_21_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_21_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_21_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_21_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_21_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_21_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_21_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_21_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_21_ldst;	// rob.scala:310:28
  reg              rob_uop_1_21_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_21_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_21_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_22_uopc;	// rob.scala:310:28
  reg              rob_uop_1_22_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_22_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_22_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_22_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_22_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_22_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_22_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_22_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_22_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_22_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_22_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_22_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_22_ldst;	// rob.scala:310:28
  reg              rob_uop_1_22_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_22_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_22_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_23_uopc;	// rob.scala:310:28
  reg              rob_uop_1_23_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_23_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_23_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_23_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_23_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_23_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_23_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_23_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_23_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_23_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_23_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_23_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_23_ldst;	// rob.scala:310:28
  reg              rob_uop_1_23_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_23_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_23_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_24_uopc;	// rob.scala:310:28
  reg              rob_uop_1_24_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_24_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_24_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_24_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_24_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_24_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_24_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_24_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_24_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_24_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_24_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_24_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_24_ldst;	// rob.scala:310:28
  reg              rob_uop_1_24_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_24_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_24_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_25_uopc;	// rob.scala:310:28
  reg              rob_uop_1_25_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_25_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_25_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_25_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_25_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_25_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_25_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_25_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_25_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_25_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_25_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_25_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_25_ldst;	// rob.scala:310:28
  reg              rob_uop_1_25_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_25_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_25_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_26_uopc;	// rob.scala:310:28
  reg              rob_uop_1_26_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_26_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_26_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_26_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_26_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_26_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_26_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_26_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_26_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_26_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_26_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_26_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_26_ldst;	// rob.scala:310:28
  reg              rob_uop_1_26_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_26_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_26_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_27_uopc;	// rob.scala:310:28
  reg              rob_uop_1_27_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_27_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_27_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_27_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_27_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_27_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_27_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_27_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_27_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_27_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_27_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_27_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_27_ldst;	// rob.scala:310:28
  reg              rob_uop_1_27_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_27_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_27_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_28_uopc;	// rob.scala:310:28
  reg              rob_uop_1_28_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_28_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_28_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_28_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_28_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_28_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_28_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_28_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_28_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_28_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_28_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_28_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_28_ldst;	// rob.scala:310:28
  reg              rob_uop_1_28_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_28_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_28_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_29_uopc;	// rob.scala:310:28
  reg              rob_uop_1_29_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_29_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_29_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_29_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_29_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_29_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_29_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_29_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_29_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_29_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_29_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_29_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_29_ldst;	// rob.scala:310:28
  reg              rob_uop_1_29_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_29_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_29_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_30_uopc;	// rob.scala:310:28
  reg              rob_uop_1_30_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_30_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_30_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_30_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_30_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_30_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_30_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_30_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_30_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_30_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_30_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_30_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_30_ldst;	// rob.scala:310:28
  reg              rob_uop_1_30_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_30_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_30_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_31_uopc;	// rob.scala:310:28
  reg              rob_uop_1_31_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_1_31_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_31_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_31_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_31_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_31_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_31_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_31_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_31_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_31_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_31_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_31_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_31_ldst;	// rob.scala:310:28
  reg              rob_uop_1_31_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_31_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_31_fp_val;	// rob.scala:310:28
  reg              rob_exception_1_0;	// rob.scala:311:28
  reg              rob_exception_1_1;	// rob.scala:311:28
  reg              rob_exception_1_2;	// rob.scala:311:28
  reg              rob_exception_1_3;	// rob.scala:311:28
  reg              rob_exception_1_4;	// rob.scala:311:28
  reg              rob_exception_1_5;	// rob.scala:311:28
  reg              rob_exception_1_6;	// rob.scala:311:28
  reg              rob_exception_1_7;	// rob.scala:311:28
  reg              rob_exception_1_8;	// rob.scala:311:28
  reg              rob_exception_1_9;	// rob.scala:311:28
  reg              rob_exception_1_10;	// rob.scala:311:28
  reg              rob_exception_1_11;	// rob.scala:311:28
  reg              rob_exception_1_12;	// rob.scala:311:28
  reg              rob_exception_1_13;	// rob.scala:311:28
  reg              rob_exception_1_14;	// rob.scala:311:28
  reg              rob_exception_1_15;	// rob.scala:311:28
  reg              rob_exception_1_16;	// rob.scala:311:28
  reg              rob_exception_1_17;	// rob.scala:311:28
  reg              rob_exception_1_18;	// rob.scala:311:28
  reg              rob_exception_1_19;	// rob.scala:311:28
  reg              rob_exception_1_20;	// rob.scala:311:28
  reg              rob_exception_1_21;	// rob.scala:311:28
  reg              rob_exception_1_22;	// rob.scala:311:28
  reg              rob_exception_1_23;	// rob.scala:311:28
  reg              rob_exception_1_24;	// rob.scala:311:28
  reg              rob_exception_1_25;	// rob.scala:311:28
  reg              rob_exception_1_26;	// rob.scala:311:28
  reg              rob_exception_1_27;	// rob.scala:311:28
  reg              rob_exception_1_28;	// rob.scala:311:28
  reg              rob_exception_1_29;	// rob.scala:311:28
  reg              rob_exception_1_30;	// rob.scala:311:28
  reg              rob_exception_1_31;	// rob.scala:311:28
  reg              rob_predicated_1_0;	// rob.scala:312:29
  reg              rob_predicated_1_1;	// rob.scala:312:29
  reg              rob_predicated_1_2;	// rob.scala:312:29
  reg              rob_predicated_1_3;	// rob.scala:312:29
  reg              rob_predicated_1_4;	// rob.scala:312:29
  reg              rob_predicated_1_5;	// rob.scala:312:29
  reg              rob_predicated_1_6;	// rob.scala:312:29
  reg              rob_predicated_1_7;	// rob.scala:312:29
  reg              rob_predicated_1_8;	// rob.scala:312:29
  reg              rob_predicated_1_9;	// rob.scala:312:29
  reg              rob_predicated_1_10;	// rob.scala:312:29
  reg              rob_predicated_1_11;	// rob.scala:312:29
  reg              rob_predicated_1_12;	// rob.scala:312:29
  reg              rob_predicated_1_13;	// rob.scala:312:29
  reg              rob_predicated_1_14;	// rob.scala:312:29
  reg              rob_predicated_1_15;	// rob.scala:312:29
  reg              rob_predicated_1_16;	// rob.scala:312:29
  reg              rob_predicated_1_17;	// rob.scala:312:29
  reg              rob_predicated_1_18;	// rob.scala:312:29
  reg              rob_predicated_1_19;	// rob.scala:312:29
  reg              rob_predicated_1_20;	// rob.scala:312:29
  reg              rob_predicated_1_21;	// rob.scala:312:29
  reg              rob_predicated_1_22;	// rob.scala:312:29
  reg              rob_predicated_1_23;	// rob.scala:312:29
  reg              rob_predicated_1_24;	// rob.scala:312:29
  reg              rob_predicated_1_25;	// rob.scala:312:29
  reg              rob_predicated_1_26;	// rob.scala:312:29
  reg              rob_predicated_1_27;	// rob.scala:312:29
  reg              rob_predicated_1_28;	// rob.scala:312:29
  reg              rob_predicated_1_29;	// rob.scala:312:29
  reg              rob_predicated_1_30;	// rob.scala:312:29
  reg              rob_predicated_1_31;	// rob.scala:312:29
  wire [31:0]      _GEN_34 =
    {{rob_val_1_31},
     {rob_val_1_30},
     {rob_val_1_29},
     {rob_val_1_28},
     {rob_val_1_27},
     {rob_val_1_26},
     {rob_val_1_25},
     {rob_val_1_24},
     {rob_val_1_23},
     {rob_val_1_22},
     {rob_val_1_21},
     {rob_val_1_20},
     {rob_val_1_19},
     {rob_val_1_18},
     {rob_val_1_17},
     {rob_val_1_16},
     {rob_val_1_15},
     {rob_val_1_14},
     {rob_val_1_13},
     {rob_val_1_12},
     {rob_val_1_11},
     {rob_val_1_10},
     {rob_val_1_9},
     {rob_val_1_8},
     {rob_val_1_7},
     {rob_val_1_6},
     {rob_val_1_5},
     {rob_val_1_4},
     {rob_val_1_3},
     {rob_val_1_2},
     {rob_val_1_1},
     {rob_val_1_0}};	// rob.scala:307:32, :324:31
  wire             rob_tail_vals_1 = _GEN_34[rob_tail];	// rob.scala:228:29, :324:31
  wire             _GEN_35 =
    io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_36 =
    io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_37 =
    io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_38 =
    io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_39 =
    io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_40 =
    io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_41 =
    io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_42 =
    io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_43 =
    io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_44 =
    io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_45 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :361:31, :540:33
  wire [31:0]      _GEN_46 =
    {{rob_bsy_1_31},
     {rob_bsy_1_30},
     {rob_bsy_1_29},
     {rob_bsy_1_28},
     {rob_bsy_1_27},
     {rob_bsy_1_26},
     {rob_bsy_1_25},
     {rob_bsy_1_24},
     {rob_bsy_1_23},
     {rob_bsy_1_22},
     {rob_bsy_1_21},
     {rob_bsy_1_20},
     {rob_bsy_1_19},
     {rob_bsy_1_18},
     {rob_bsy_1_17},
     {rob_bsy_1_16},
     {rob_bsy_1_15},
     {rob_bsy_1_14},
     {rob_bsy_1_13},
     {rob_bsy_1_12},
     {rob_bsy_1_11},
     {rob_bsy_1_10},
     {rob_bsy_1_9},
     {rob_bsy_1_8},
     {rob_bsy_1_7},
     {rob_bsy_1_6},
     {rob_bsy_1_5},
     {rob_bsy_1_4},
     {rob_bsy_1_3},
     {rob_bsy_1_2},
     {rob_bsy_1_1},
     {rob_bsy_1_0}};	// rob.scala:308:28, :366:31
  wire             _GEN_47 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :361:31, :540:33
  wire             _GEN_48 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :361:31, :540:33
  wire             _GEN_49 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :390:26, :540:33
  wire [31:0]      _GEN_50 =
    {{rob_unsafe_1_31},
     {rob_unsafe_1_30},
     {rob_unsafe_1_29},
     {rob_unsafe_1_28},
     {rob_unsafe_1_27},
     {rob_unsafe_1_26},
     {rob_unsafe_1_25},
     {rob_unsafe_1_24},
     {rob_unsafe_1_23},
     {rob_unsafe_1_22},
     {rob_unsafe_1_21},
     {rob_unsafe_1_20},
     {rob_unsafe_1_19},
     {rob_unsafe_1_18},
     {rob_unsafe_1_17},
     {rob_unsafe_1_16},
     {rob_unsafe_1_15},
     {rob_unsafe_1_14},
     {rob_unsafe_1_13},
     {rob_unsafe_1_12},
     {rob_unsafe_1_11},
     {rob_unsafe_1_10},
     {rob_unsafe_1_9},
     {rob_unsafe_1_8},
     {rob_unsafe_1_7},
     {rob_unsafe_1_6},
     {rob_unsafe_1_5},
     {rob_unsafe_1_4},
     {rob_unsafe_1_3},
     {rob_unsafe_1_2},
     {rob_unsafe_1_1},
     {rob_unsafe_1_0}};	// rob.scala:309:28, :394:15
  wire             rob_head_vals_1 = _GEN_34[rob_head];	// rob.scala:224:29, :324:31, :398:49
  wire [31:0]      _GEN_51 =
    {{rob_exception_1_31},
     {rob_exception_1_30},
     {rob_exception_1_29},
     {rob_exception_1_28},
     {rob_exception_1_27},
     {rob_exception_1_26},
     {rob_exception_1_25},
     {rob_exception_1_24},
     {rob_exception_1_23},
     {rob_exception_1_22},
     {rob_exception_1_21},
     {rob_exception_1_20},
     {rob_exception_1_19},
     {rob_exception_1_18},
     {rob_exception_1_17},
     {rob_exception_1_16},
     {rob_exception_1_15},
     {rob_exception_1_14},
     {rob_exception_1_13},
     {rob_exception_1_12},
     {rob_exception_1_11},
     {rob_exception_1_10},
     {rob_exception_1_9},
     {rob_exception_1_8},
     {rob_exception_1_7},
     {rob_exception_1_6},
     {rob_exception_1_5},
     {rob_exception_1_4},
     {rob_exception_1_3},
     {rob_exception_1_2},
     {rob_exception_1_1},
     {rob_exception_1_0}};	// rob.scala:311:28, :398:49
  wire             can_throw_exception_1 = rob_head_vals_1 & _GEN_51[rob_head];	// rob.scala:224:29, :398:49
  wire             can_commit_1 = rob_head_vals_1 & ~_GEN_46[rob_head] & ~io_csr_stall;	// rob.scala:224:29, :366:31, :398:49, :404:{43,64,67}
  wire [31:0]      _GEN_52 =
    {{rob_predicated_1_31},
     {rob_predicated_1_30},
     {rob_predicated_1_29},
     {rob_predicated_1_28},
     {rob_predicated_1_27},
     {rob_predicated_1_26},
     {rob_predicated_1_25},
     {rob_predicated_1_24},
     {rob_predicated_1_23},
     {rob_predicated_1_22},
     {rob_predicated_1_21},
     {rob_predicated_1_20},
     {rob_predicated_1_19},
     {rob_predicated_1_18},
     {rob_predicated_1_17},
     {rob_predicated_1_16},
     {rob_predicated_1_15},
     {rob_predicated_1_14},
     {rob_predicated_1_13},
     {rob_predicated_1_12},
     {rob_predicated_1_11},
     {rob_predicated_1_10},
     {rob_predicated_1_9},
     {rob_predicated_1_8},
     {rob_predicated_1_7},
     {rob_predicated_1_6},
     {rob_predicated_1_5},
     {rob_predicated_1_4},
     {rob_predicated_1_3},
     {rob_predicated_1_2},
     {rob_predicated_1_1},
     {rob_predicated_1_0}};	// rob.scala:312:29, :410:51
  wire [31:0][6:0] _GEN_53 =
    {{rob_uop_1_31_uopc},
     {rob_uop_1_30_uopc},
     {rob_uop_1_29_uopc},
     {rob_uop_1_28_uopc},
     {rob_uop_1_27_uopc},
     {rob_uop_1_26_uopc},
     {rob_uop_1_25_uopc},
     {rob_uop_1_24_uopc},
     {rob_uop_1_23_uopc},
     {rob_uop_1_22_uopc},
     {rob_uop_1_21_uopc},
     {rob_uop_1_20_uopc},
     {rob_uop_1_19_uopc},
     {rob_uop_1_18_uopc},
     {rob_uop_1_17_uopc},
     {rob_uop_1_16_uopc},
     {rob_uop_1_15_uopc},
     {rob_uop_1_14_uopc},
     {rob_uop_1_13_uopc},
     {rob_uop_1_12_uopc},
     {rob_uop_1_11_uopc},
     {rob_uop_1_10_uopc},
     {rob_uop_1_9_uopc},
     {rob_uop_1_8_uopc},
     {rob_uop_1_7_uopc},
     {rob_uop_1_6_uopc},
     {rob_uop_1_5_uopc},
     {rob_uop_1_4_uopc},
     {rob_uop_1_3_uopc},
     {rob_uop_1_2_uopc},
     {rob_uop_1_1_uopc},
     {rob_uop_1_0_uopc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_54 =
    {{rob_uop_1_31_is_rvc},
     {rob_uop_1_30_is_rvc},
     {rob_uop_1_29_is_rvc},
     {rob_uop_1_28_is_rvc},
     {rob_uop_1_27_is_rvc},
     {rob_uop_1_26_is_rvc},
     {rob_uop_1_25_is_rvc},
     {rob_uop_1_24_is_rvc},
     {rob_uop_1_23_is_rvc},
     {rob_uop_1_22_is_rvc},
     {rob_uop_1_21_is_rvc},
     {rob_uop_1_20_is_rvc},
     {rob_uop_1_19_is_rvc},
     {rob_uop_1_18_is_rvc},
     {rob_uop_1_17_is_rvc},
     {rob_uop_1_16_is_rvc},
     {rob_uop_1_15_is_rvc},
     {rob_uop_1_14_is_rvc},
     {rob_uop_1_13_is_rvc},
     {rob_uop_1_12_is_rvc},
     {rob_uop_1_11_is_rvc},
     {rob_uop_1_10_is_rvc},
     {rob_uop_1_9_is_rvc},
     {rob_uop_1_8_is_rvc},
     {rob_uop_1_7_is_rvc},
     {rob_uop_1_6_is_rvc},
     {rob_uop_1_5_is_rvc},
     {rob_uop_1_4_is_rvc},
     {rob_uop_1_3_is_rvc},
     {rob_uop_1_2_is_rvc},
     {rob_uop_1_1_is_rvc},
     {rob_uop_1_0_is_rvc}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_55 =
    {{rob_uop_1_31_ftq_idx},
     {rob_uop_1_30_ftq_idx},
     {rob_uop_1_29_ftq_idx},
     {rob_uop_1_28_ftq_idx},
     {rob_uop_1_27_ftq_idx},
     {rob_uop_1_26_ftq_idx},
     {rob_uop_1_25_ftq_idx},
     {rob_uop_1_24_ftq_idx},
     {rob_uop_1_23_ftq_idx},
     {rob_uop_1_22_ftq_idx},
     {rob_uop_1_21_ftq_idx},
     {rob_uop_1_20_ftq_idx},
     {rob_uop_1_19_ftq_idx},
     {rob_uop_1_18_ftq_idx},
     {rob_uop_1_17_ftq_idx},
     {rob_uop_1_16_ftq_idx},
     {rob_uop_1_15_ftq_idx},
     {rob_uop_1_14_ftq_idx},
     {rob_uop_1_13_ftq_idx},
     {rob_uop_1_12_ftq_idx},
     {rob_uop_1_11_ftq_idx},
     {rob_uop_1_10_ftq_idx},
     {rob_uop_1_9_ftq_idx},
     {rob_uop_1_8_ftq_idx},
     {rob_uop_1_7_ftq_idx},
     {rob_uop_1_6_ftq_idx},
     {rob_uop_1_5_ftq_idx},
     {rob_uop_1_4_ftq_idx},
     {rob_uop_1_3_ftq_idx},
     {rob_uop_1_2_ftq_idx},
     {rob_uop_1_1_ftq_idx},
     {rob_uop_1_0_ftq_idx}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_56 =
    {{rob_uop_1_31_edge_inst},
     {rob_uop_1_30_edge_inst},
     {rob_uop_1_29_edge_inst},
     {rob_uop_1_28_edge_inst},
     {rob_uop_1_27_edge_inst},
     {rob_uop_1_26_edge_inst},
     {rob_uop_1_25_edge_inst},
     {rob_uop_1_24_edge_inst},
     {rob_uop_1_23_edge_inst},
     {rob_uop_1_22_edge_inst},
     {rob_uop_1_21_edge_inst},
     {rob_uop_1_20_edge_inst},
     {rob_uop_1_19_edge_inst},
     {rob_uop_1_18_edge_inst},
     {rob_uop_1_17_edge_inst},
     {rob_uop_1_16_edge_inst},
     {rob_uop_1_15_edge_inst},
     {rob_uop_1_14_edge_inst},
     {rob_uop_1_13_edge_inst},
     {rob_uop_1_12_edge_inst},
     {rob_uop_1_11_edge_inst},
     {rob_uop_1_10_edge_inst},
     {rob_uop_1_9_edge_inst},
     {rob_uop_1_8_edge_inst},
     {rob_uop_1_7_edge_inst},
     {rob_uop_1_6_edge_inst},
     {rob_uop_1_5_edge_inst},
     {rob_uop_1_4_edge_inst},
     {rob_uop_1_3_edge_inst},
     {rob_uop_1_2_edge_inst},
     {rob_uop_1_1_edge_inst},
     {rob_uop_1_0_edge_inst}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_57 =
    {{rob_uop_1_31_pc_lob},
     {rob_uop_1_30_pc_lob},
     {rob_uop_1_29_pc_lob},
     {rob_uop_1_28_pc_lob},
     {rob_uop_1_27_pc_lob},
     {rob_uop_1_26_pc_lob},
     {rob_uop_1_25_pc_lob},
     {rob_uop_1_24_pc_lob},
     {rob_uop_1_23_pc_lob},
     {rob_uop_1_22_pc_lob},
     {rob_uop_1_21_pc_lob},
     {rob_uop_1_20_pc_lob},
     {rob_uop_1_19_pc_lob},
     {rob_uop_1_18_pc_lob},
     {rob_uop_1_17_pc_lob},
     {rob_uop_1_16_pc_lob},
     {rob_uop_1_15_pc_lob},
     {rob_uop_1_14_pc_lob},
     {rob_uop_1_13_pc_lob},
     {rob_uop_1_12_pc_lob},
     {rob_uop_1_11_pc_lob},
     {rob_uop_1_10_pc_lob},
     {rob_uop_1_9_pc_lob},
     {rob_uop_1_8_pc_lob},
     {rob_uop_1_7_pc_lob},
     {rob_uop_1_6_pc_lob},
     {rob_uop_1_5_pc_lob},
     {rob_uop_1_4_pc_lob},
     {rob_uop_1_3_pc_lob},
     {rob_uop_1_2_pc_lob},
     {rob_uop_1_1_pc_lob},
     {rob_uop_1_0_pc_lob}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_58 =
    {{rob_uop_1_31_pdst},
     {rob_uop_1_30_pdst},
     {rob_uop_1_29_pdst},
     {rob_uop_1_28_pdst},
     {rob_uop_1_27_pdst},
     {rob_uop_1_26_pdst},
     {rob_uop_1_25_pdst},
     {rob_uop_1_24_pdst},
     {rob_uop_1_23_pdst},
     {rob_uop_1_22_pdst},
     {rob_uop_1_21_pdst},
     {rob_uop_1_20_pdst},
     {rob_uop_1_19_pdst},
     {rob_uop_1_18_pdst},
     {rob_uop_1_17_pdst},
     {rob_uop_1_16_pdst},
     {rob_uop_1_15_pdst},
     {rob_uop_1_14_pdst},
     {rob_uop_1_13_pdst},
     {rob_uop_1_12_pdst},
     {rob_uop_1_11_pdst},
     {rob_uop_1_10_pdst},
     {rob_uop_1_9_pdst},
     {rob_uop_1_8_pdst},
     {rob_uop_1_7_pdst},
     {rob_uop_1_6_pdst},
     {rob_uop_1_5_pdst},
     {rob_uop_1_4_pdst},
     {rob_uop_1_3_pdst},
     {rob_uop_1_2_pdst},
     {rob_uop_1_1_pdst},
     {rob_uop_1_0_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_59 =
    {{rob_uop_1_31_stale_pdst},
     {rob_uop_1_30_stale_pdst},
     {rob_uop_1_29_stale_pdst},
     {rob_uop_1_28_stale_pdst},
     {rob_uop_1_27_stale_pdst},
     {rob_uop_1_26_stale_pdst},
     {rob_uop_1_25_stale_pdst},
     {rob_uop_1_24_stale_pdst},
     {rob_uop_1_23_stale_pdst},
     {rob_uop_1_22_stale_pdst},
     {rob_uop_1_21_stale_pdst},
     {rob_uop_1_20_stale_pdst},
     {rob_uop_1_19_stale_pdst},
     {rob_uop_1_18_stale_pdst},
     {rob_uop_1_17_stale_pdst},
     {rob_uop_1_16_stale_pdst},
     {rob_uop_1_15_stale_pdst},
     {rob_uop_1_14_stale_pdst},
     {rob_uop_1_13_stale_pdst},
     {rob_uop_1_12_stale_pdst},
     {rob_uop_1_11_stale_pdst},
     {rob_uop_1_10_stale_pdst},
     {rob_uop_1_9_stale_pdst},
     {rob_uop_1_8_stale_pdst},
     {rob_uop_1_7_stale_pdst},
     {rob_uop_1_6_stale_pdst},
     {rob_uop_1_5_stale_pdst},
     {rob_uop_1_4_stale_pdst},
     {rob_uop_1_3_stale_pdst},
     {rob_uop_1_2_stale_pdst},
     {rob_uop_1_1_stale_pdst},
     {rob_uop_1_0_stale_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_60 =
    {{rob_uop_1_31_is_fencei},
     {rob_uop_1_30_is_fencei},
     {rob_uop_1_29_is_fencei},
     {rob_uop_1_28_is_fencei},
     {rob_uop_1_27_is_fencei},
     {rob_uop_1_26_is_fencei},
     {rob_uop_1_25_is_fencei},
     {rob_uop_1_24_is_fencei},
     {rob_uop_1_23_is_fencei},
     {rob_uop_1_22_is_fencei},
     {rob_uop_1_21_is_fencei},
     {rob_uop_1_20_is_fencei},
     {rob_uop_1_19_is_fencei},
     {rob_uop_1_18_is_fencei},
     {rob_uop_1_17_is_fencei},
     {rob_uop_1_16_is_fencei},
     {rob_uop_1_15_is_fencei},
     {rob_uop_1_14_is_fencei},
     {rob_uop_1_13_is_fencei},
     {rob_uop_1_12_is_fencei},
     {rob_uop_1_11_is_fencei},
     {rob_uop_1_10_is_fencei},
     {rob_uop_1_9_is_fencei},
     {rob_uop_1_8_is_fencei},
     {rob_uop_1_7_is_fencei},
     {rob_uop_1_6_is_fencei},
     {rob_uop_1_5_is_fencei},
     {rob_uop_1_4_is_fencei},
     {rob_uop_1_3_is_fencei},
     {rob_uop_1_2_is_fencei},
     {rob_uop_1_1_is_fencei},
     {rob_uop_1_0_is_fencei}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_61 =
    {{rob_uop_1_31_uses_ldq},
     {rob_uop_1_30_uses_ldq},
     {rob_uop_1_29_uses_ldq},
     {rob_uop_1_28_uses_ldq},
     {rob_uop_1_27_uses_ldq},
     {rob_uop_1_26_uses_ldq},
     {rob_uop_1_25_uses_ldq},
     {rob_uop_1_24_uses_ldq},
     {rob_uop_1_23_uses_ldq},
     {rob_uop_1_22_uses_ldq},
     {rob_uop_1_21_uses_ldq},
     {rob_uop_1_20_uses_ldq},
     {rob_uop_1_19_uses_ldq},
     {rob_uop_1_18_uses_ldq},
     {rob_uop_1_17_uses_ldq},
     {rob_uop_1_16_uses_ldq},
     {rob_uop_1_15_uses_ldq},
     {rob_uop_1_14_uses_ldq},
     {rob_uop_1_13_uses_ldq},
     {rob_uop_1_12_uses_ldq},
     {rob_uop_1_11_uses_ldq},
     {rob_uop_1_10_uses_ldq},
     {rob_uop_1_9_uses_ldq},
     {rob_uop_1_8_uses_ldq},
     {rob_uop_1_7_uses_ldq},
     {rob_uop_1_6_uses_ldq},
     {rob_uop_1_5_uses_ldq},
     {rob_uop_1_4_uses_ldq},
     {rob_uop_1_3_uses_ldq},
     {rob_uop_1_2_uses_ldq},
     {rob_uop_1_1_uses_ldq},
     {rob_uop_1_0_uses_ldq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_62 =
    {{rob_uop_1_31_uses_stq},
     {rob_uop_1_30_uses_stq},
     {rob_uop_1_29_uses_stq},
     {rob_uop_1_28_uses_stq},
     {rob_uop_1_27_uses_stq},
     {rob_uop_1_26_uses_stq},
     {rob_uop_1_25_uses_stq},
     {rob_uop_1_24_uses_stq},
     {rob_uop_1_23_uses_stq},
     {rob_uop_1_22_uses_stq},
     {rob_uop_1_21_uses_stq},
     {rob_uop_1_20_uses_stq},
     {rob_uop_1_19_uses_stq},
     {rob_uop_1_18_uses_stq},
     {rob_uop_1_17_uses_stq},
     {rob_uop_1_16_uses_stq},
     {rob_uop_1_15_uses_stq},
     {rob_uop_1_14_uses_stq},
     {rob_uop_1_13_uses_stq},
     {rob_uop_1_12_uses_stq},
     {rob_uop_1_11_uses_stq},
     {rob_uop_1_10_uses_stq},
     {rob_uop_1_9_uses_stq},
     {rob_uop_1_8_uses_stq},
     {rob_uop_1_7_uses_stq},
     {rob_uop_1_6_uses_stq},
     {rob_uop_1_5_uses_stq},
     {rob_uop_1_4_uses_stq},
     {rob_uop_1_3_uses_stq},
     {rob_uop_1_2_uses_stq},
     {rob_uop_1_1_uses_stq},
     {rob_uop_1_0_uses_stq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_63 =
    {{rob_uop_1_31_is_sys_pc2epc},
     {rob_uop_1_30_is_sys_pc2epc},
     {rob_uop_1_29_is_sys_pc2epc},
     {rob_uop_1_28_is_sys_pc2epc},
     {rob_uop_1_27_is_sys_pc2epc},
     {rob_uop_1_26_is_sys_pc2epc},
     {rob_uop_1_25_is_sys_pc2epc},
     {rob_uop_1_24_is_sys_pc2epc},
     {rob_uop_1_23_is_sys_pc2epc},
     {rob_uop_1_22_is_sys_pc2epc},
     {rob_uop_1_21_is_sys_pc2epc},
     {rob_uop_1_20_is_sys_pc2epc},
     {rob_uop_1_19_is_sys_pc2epc},
     {rob_uop_1_18_is_sys_pc2epc},
     {rob_uop_1_17_is_sys_pc2epc},
     {rob_uop_1_16_is_sys_pc2epc},
     {rob_uop_1_15_is_sys_pc2epc},
     {rob_uop_1_14_is_sys_pc2epc},
     {rob_uop_1_13_is_sys_pc2epc},
     {rob_uop_1_12_is_sys_pc2epc},
     {rob_uop_1_11_is_sys_pc2epc},
     {rob_uop_1_10_is_sys_pc2epc},
     {rob_uop_1_9_is_sys_pc2epc},
     {rob_uop_1_8_is_sys_pc2epc},
     {rob_uop_1_7_is_sys_pc2epc},
     {rob_uop_1_6_is_sys_pc2epc},
     {rob_uop_1_5_is_sys_pc2epc},
     {rob_uop_1_4_is_sys_pc2epc},
     {rob_uop_1_3_is_sys_pc2epc},
     {rob_uop_1_2_is_sys_pc2epc},
     {rob_uop_1_1_is_sys_pc2epc},
     {rob_uop_1_0_is_sys_pc2epc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_64 =
    {{rob_uop_1_31_flush_on_commit},
     {rob_uop_1_30_flush_on_commit},
     {rob_uop_1_29_flush_on_commit},
     {rob_uop_1_28_flush_on_commit},
     {rob_uop_1_27_flush_on_commit},
     {rob_uop_1_26_flush_on_commit},
     {rob_uop_1_25_flush_on_commit},
     {rob_uop_1_24_flush_on_commit},
     {rob_uop_1_23_flush_on_commit},
     {rob_uop_1_22_flush_on_commit},
     {rob_uop_1_21_flush_on_commit},
     {rob_uop_1_20_flush_on_commit},
     {rob_uop_1_19_flush_on_commit},
     {rob_uop_1_18_flush_on_commit},
     {rob_uop_1_17_flush_on_commit},
     {rob_uop_1_16_flush_on_commit},
     {rob_uop_1_15_flush_on_commit},
     {rob_uop_1_14_flush_on_commit},
     {rob_uop_1_13_flush_on_commit},
     {rob_uop_1_12_flush_on_commit},
     {rob_uop_1_11_flush_on_commit},
     {rob_uop_1_10_flush_on_commit},
     {rob_uop_1_9_flush_on_commit},
     {rob_uop_1_8_flush_on_commit},
     {rob_uop_1_7_flush_on_commit},
     {rob_uop_1_6_flush_on_commit},
     {rob_uop_1_5_flush_on_commit},
     {rob_uop_1_4_flush_on_commit},
     {rob_uop_1_3_flush_on_commit},
     {rob_uop_1_2_flush_on_commit},
     {rob_uop_1_1_flush_on_commit},
     {rob_uop_1_0_flush_on_commit}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_65 =
    {{rob_uop_1_31_ldst},
     {rob_uop_1_30_ldst},
     {rob_uop_1_29_ldst},
     {rob_uop_1_28_ldst},
     {rob_uop_1_27_ldst},
     {rob_uop_1_26_ldst},
     {rob_uop_1_25_ldst},
     {rob_uop_1_24_ldst},
     {rob_uop_1_23_ldst},
     {rob_uop_1_22_ldst},
     {rob_uop_1_21_ldst},
     {rob_uop_1_20_ldst},
     {rob_uop_1_19_ldst},
     {rob_uop_1_18_ldst},
     {rob_uop_1_17_ldst},
     {rob_uop_1_16_ldst},
     {rob_uop_1_15_ldst},
     {rob_uop_1_14_ldst},
     {rob_uop_1_13_ldst},
     {rob_uop_1_12_ldst},
     {rob_uop_1_11_ldst},
     {rob_uop_1_10_ldst},
     {rob_uop_1_9_ldst},
     {rob_uop_1_8_ldst},
     {rob_uop_1_7_ldst},
     {rob_uop_1_6_ldst},
     {rob_uop_1_5_ldst},
     {rob_uop_1_4_ldst},
     {rob_uop_1_3_ldst},
     {rob_uop_1_2_ldst},
     {rob_uop_1_1_ldst},
     {rob_uop_1_0_ldst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_66 =
    {{rob_uop_1_31_ldst_val},
     {rob_uop_1_30_ldst_val},
     {rob_uop_1_29_ldst_val},
     {rob_uop_1_28_ldst_val},
     {rob_uop_1_27_ldst_val},
     {rob_uop_1_26_ldst_val},
     {rob_uop_1_25_ldst_val},
     {rob_uop_1_24_ldst_val},
     {rob_uop_1_23_ldst_val},
     {rob_uop_1_22_ldst_val},
     {rob_uop_1_21_ldst_val},
     {rob_uop_1_20_ldst_val},
     {rob_uop_1_19_ldst_val},
     {rob_uop_1_18_ldst_val},
     {rob_uop_1_17_ldst_val},
     {rob_uop_1_16_ldst_val},
     {rob_uop_1_15_ldst_val},
     {rob_uop_1_14_ldst_val},
     {rob_uop_1_13_ldst_val},
     {rob_uop_1_12_ldst_val},
     {rob_uop_1_11_ldst_val},
     {rob_uop_1_10_ldst_val},
     {rob_uop_1_9_ldst_val},
     {rob_uop_1_8_ldst_val},
     {rob_uop_1_7_ldst_val},
     {rob_uop_1_6_ldst_val},
     {rob_uop_1_5_ldst_val},
     {rob_uop_1_4_ldst_val},
     {rob_uop_1_3_ldst_val},
     {rob_uop_1_2_ldst_val},
     {rob_uop_1_1_ldst_val},
     {rob_uop_1_0_ldst_val}};	// rob.scala:310:28, :411:25
  wire [31:0][1:0] _GEN_67 =
    {{rob_uop_1_31_dst_rtype},
     {rob_uop_1_30_dst_rtype},
     {rob_uop_1_29_dst_rtype},
     {rob_uop_1_28_dst_rtype},
     {rob_uop_1_27_dst_rtype},
     {rob_uop_1_26_dst_rtype},
     {rob_uop_1_25_dst_rtype},
     {rob_uop_1_24_dst_rtype},
     {rob_uop_1_23_dst_rtype},
     {rob_uop_1_22_dst_rtype},
     {rob_uop_1_21_dst_rtype},
     {rob_uop_1_20_dst_rtype},
     {rob_uop_1_19_dst_rtype},
     {rob_uop_1_18_dst_rtype},
     {rob_uop_1_17_dst_rtype},
     {rob_uop_1_16_dst_rtype},
     {rob_uop_1_15_dst_rtype},
     {rob_uop_1_14_dst_rtype},
     {rob_uop_1_13_dst_rtype},
     {rob_uop_1_12_dst_rtype},
     {rob_uop_1_11_dst_rtype},
     {rob_uop_1_10_dst_rtype},
     {rob_uop_1_9_dst_rtype},
     {rob_uop_1_8_dst_rtype},
     {rob_uop_1_7_dst_rtype},
     {rob_uop_1_6_dst_rtype},
     {rob_uop_1_5_dst_rtype},
     {rob_uop_1_4_dst_rtype},
     {rob_uop_1_3_dst_rtype},
     {rob_uop_1_2_dst_rtype},
     {rob_uop_1_1_dst_rtype},
     {rob_uop_1_0_dst_rtype}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_68 =
    {{rob_uop_1_31_fp_val},
     {rob_uop_1_30_fp_val},
     {rob_uop_1_29_fp_val},
     {rob_uop_1_28_fp_val},
     {rob_uop_1_27_fp_val},
     {rob_uop_1_26_fp_val},
     {rob_uop_1_25_fp_val},
     {rob_uop_1_24_fp_val},
     {rob_uop_1_23_fp_val},
     {rob_uop_1_22_fp_val},
     {rob_uop_1_21_fp_val},
     {rob_uop_1_20_fp_val},
     {rob_uop_1_19_fp_val},
     {rob_uop_1_18_fp_val},
     {rob_uop_1_17_fp_val},
     {rob_uop_1_16_fp_val},
     {rob_uop_1_15_fp_val},
     {rob_uop_1_14_fp_val},
     {rob_uop_1_13_fp_val},
     {rob_uop_1_12_fp_val},
     {rob_uop_1_11_fp_val},
     {rob_uop_1_10_fp_val},
     {rob_uop_1_9_fp_val},
     {rob_uop_1_8_fp_val},
     {rob_uop_1_7_fp_val},
     {rob_uop_1_6_fp_val},
     {rob_uop_1_5_fp_val},
     {rob_uop_1_4_fp_val},
     {rob_uop_1_3_fp_val},
     {rob_uop_1_2_fp_val},
     {rob_uop_1_1_fp_val},
     {rob_uop_1_0_fp_val}};	// rob.scala:310:28, :411:25
  wire             rbk_row_1 = _io_commit_rollback_T_3 & ~full;	// rob.scala:236:31, :425:{44,47}, :787:39
  wire             _io_commit_rbk_valids_1_output = rbk_row_1 & _GEN_34[com_idx];	// rob.scala:236:20, :324:31, :425:44, :427:40
  reg              rob_val_2_0;	// rob.scala:307:32
  reg              rob_val_2_1;	// rob.scala:307:32
  reg              rob_val_2_2;	// rob.scala:307:32
  reg              rob_val_2_3;	// rob.scala:307:32
  reg              rob_val_2_4;	// rob.scala:307:32
  reg              rob_val_2_5;	// rob.scala:307:32
  reg              rob_val_2_6;	// rob.scala:307:32
  reg              rob_val_2_7;	// rob.scala:307:32
  reg              rob_val_2_8;	// rob.scala:307:32
  reg              rob_val_2_9;	// rob.scala:307:32
  reg              rob_val_2_10;	// rob.scala:307:32
  reg              rob_val_2_11;	// rob.scala:307:32
  reg              rob_val_2_12;	// rob.scala:307:32
  reg              rob_val_2_13;	// rob.scala:307:32
  reg              rob_val_2_14;	// rob.scala:307:32
  reg              rob_val_2_15;	// rob.scala:307:32
  reg              rob_val_2_16;	// rob.scala:307:32
  reg              rob_val_2_17;	// rob.scala:307:32
  reg              rob_val_2_18;	// rob.scala:307:32
  reg              rob_val_2_19;	// rob.scala:307:32
  reg              rob_val_2_20;	// rob.scala:307:32
  reg              rob_val_2_21;	// rob.scala:307:32
  reg              rob_val_2_22;	// rob.scala:307:32
  reg              rob_val_2_23;	// rob.scala:307:32
  reg              rob_val_2_24;	// rob.scala:307:32
  reg              rob_val_2_25;	// rob.scala:307:32
  reg              rob_val_2_26;	// rob.scala:307:32
  reg              rob_val_2_27;	// rob.scala:307:32
  reg              rob_val_2_28;	// rob.scala:307:32
  reg              rob_val_2_29;	// rob.scala:307:32
  reg              rob_val_2_30;	// rob.scala:307:32
  reg              rob_val_2_31;	// rob.scala:307:32
  reg              rob_bsy_2_0;	// rob.scala:308:28
  reg              rob_bsy_2_1;	// rob.scala:308:28
  reg              rob_bsy_2_2;	// rob.scala:308:28
  reg              rob_bsy_2_3;	// rob.scala:308:28
  reg              rob_bsy_2_4;	// rob.scala:308:28
  reg              rob_bsy_2_5;	// rob.scala:308:28
  reg              rob_bsy_2_6;	// rob.scala:308:28
  reg              rob_bsy_2_7;	// rob.scala:308:28
  reg              rob_bsy_2_8;	// rob.scala:308:28
  reg              rob_bsy_2_9;	// rob.scala:308:28
  reg              rob_bsy_2_10;	// rob.scala:308:28
  reg              rob_bsy_2_11;	// rob.scala:308:28
  reg              rob_bsy_2_12;	// rob.scala:308:28
  reg              rob_bsy_2_13;	// rob.scala:308:28
  reg              rob_bsy_2_14;	// rob.scala:308:28
  reg              rob_bsy_2_15;	// rob.scala:308:28
  reg              rob_bsy_2_16;	// rob.scala:308:28
  reg              rob_bsy_2_17;	// rob.scala:308:28
  reg              rob_bsy_2_18;	// rob.scala:308:28
  reg              rob_bsy_2_19;	// rob.scala:308:28
  reg              rob_bsy_2_20;	// rob.scala:308:28
  reg              rob_bsy_2_21;	// rob.scala:308:28
  reg              rob_bsy_2_22;	// rob.scala:308:28
  reg              rob_bsy_2_23;	// rob.scala:308:28
  reg              rob_bsy_2_24;	// rob.scala:308:28
  reg              rob_bsy_2_25;	// rob.scala:308:28
  reg              rob_bsy_2_26;	// rob.scala:308:28
  reg              rob_bsy_2_27;	// rob.scala:308:28
  reg              rob_bsy_2_28;	// rob.scala:308:28
  reg              rob_bsy_2_29;	// rob.scala:308:28
  reg              rob_bsy_2_30;	// rob.scala:308:28
  reg              rob_bsy_2_31;	// rob.scala:308:28
  reg              rob_unsafe_2_0;	// rob.scala:309:28
  reg              rob_unsafe_2_1;	// rob.scala:309:28
  reg              rob_unsafe_2_2;	// rob.scala:309:28
  reg              rob_unsafe_2_3;	// rob.scala:309:28
  reg              rob_unsafe_2_4;	// rob.scala:309:28
  reg              rob_unsafe_2_5;	// rob.scala:309:28
  reg              rob_unsafe_2_6;	// rob.scala:309:28
  reg              rob_unsafe_2_7;	// rob.scala:309:28
  reg              rob_unsafe_2_8;	// rob.scala:309:28
  reg              rob_unsafe_2_9;	// rob.scala:309:28
  reg              rob_unsafe_2_10;	// rob.scala:309:28
  reg              rob_unsafe_2_11;	// rob.scala:309:28
  reg              rob_unsafe_2_12;	// rob.scala:309:28
  reg              rob_unsafe_2_13;	// rob.scala:309:28
  reg              rob_unsafe_2_14;	// rob.scala:309:28
  reg              rob_unsafe_2_15;	// rob.scala:309:28
  reg              rob_unsafe_2_16;	// rob.scala:309:28
  reg              rob_unsafe_2_17;	// rob.scala:309:28
  reg              rob_unsafe_2_18;	// rob.scala:309:28
  reg              rob_unsafe_2_19;	// rob.scala:309:28
  reg              rob_unsafe_2_20;	// rob.scala:309:28
  reg              rob_unsafe_2_21;	// rob.scala:309:28
  reg              rob_unsafe_2_22;	// rob.scala:309:28
  reg              rob_unsafe_2_23;	// rob.scala:309:28
  reg              rob_unsafe_2_24;	// rob.scala:309:28
  reg              rob_unsafe_2_25;	// rob.scala:309:28
  reg              rob_unsafe_2_26;	// rob.scala:309:28
  reg              rob_unsafe_2_27;	// rob.scala:309:28
  reg              rob_unsafe_2_28;	// rob.scala:309:28
  reg              rob_unsafe_2_29;	// rob.scala:309:28
  reg              rob_unsafe_2_30;	// rob.scala:309:28
  reg              rob_unsafe_2_31;	// rob.scala:309:28
  reg  [6:0]       rob_uop_2_0_uopc;	// rob.scala:310:28
  reg              rob_uop_2_0_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_0_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_0_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_0_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_0_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_0_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_0_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_0_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_0_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_0_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_0_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_0_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_0_ldst;	// rob.scala:310:28
  reg              rob_uop_2_0_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_0_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_0_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_1_uopc;	// rob.scala:310:28
  reg              rob_uop_2_1_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_1_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_1_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_1_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_1_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_1_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_1_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_1_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_1_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_1_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_1_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_1_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_1_ldst;	// rob.scala:310:28
  reg              rob_uop_2_1_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_1_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_1_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_2_uopc;	// rob.scala:310:28
  reg              rob_uop_2_2_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_2_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_2_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_2_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_2_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_2_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_2_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_2_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_2_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_2_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_2_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_2_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_2_ldst;	// rob.scala:310:28
  reg              rob_uop_2_2_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_2_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_2_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_3_uopc;	// rob.scala:310:28
  reg              rob_uop_2_3_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_3_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_3_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_3_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_3_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_3_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_3_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_3_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_3_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_3_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_3_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_3_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_3_ldst;	// rob.scala:310:28
  reg              rob_uop_2_3_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_3_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_3_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_4_uopc;	// rob.scala:310:28
  reg              rob_uop_2_4_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_4_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_4_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_4_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_4_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_4_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_4_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_4_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_4_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_4_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_4_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_4_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_4_ldst;	// rob.scala:310:28
  reg              rob_uop_2_4_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_4_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_4_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_5_uopc;	// rob.scala:310:28
  reg              rob_uop_2_5_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_5_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_5_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_5_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_5_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_5_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_5_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_5_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_5_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_5_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_5_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_5_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_5_ldst;	// rob.scala:310:28
  reg              rob_uop_2_5_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_5_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_5_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_6_uopc;	// rob.scala:310:28
  reg              rob_uop_2_6_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_6_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_6_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_6_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_6_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_6_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_6_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_6_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_6_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_6_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_6_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_6_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_6_ldst;	// rob.scala:310:28
  reg              rob_uop_2_6_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_6_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_6_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_7_uopc;	// rob.scala:310:28
  reg              rob_uop_2_7_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_7_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_7_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_7_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_7_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_7_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_7_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_7_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_7_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_7_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_7_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_7_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_7_ldst;	// rob.scala:310:28
  reg              rob_uop_2_7_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_7_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_7_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_8_uopc;	// rob.scala:310:28
  reg              rob_uop_2_8_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_8_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_8_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_8_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_8_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_8_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_8_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_8_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_8_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_8_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_8_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_8_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_8_ldst;	// rob.scala:310:28
  reg              rob_uop_2_8_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_8_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_8_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_9_uopc;	// rob.scala:310:28
  reg              rob_uop_2_9_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_9_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_9_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_9_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_9_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_9_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_9_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_9_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_9_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_9_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_9_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_9_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_9_ldst;	// rob.scala:310:28
  reg              rob_uop_2_9_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_9_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_9_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_10_uopc;	// rob.scala:310:28
  reg              rob_uop_2_10_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_10_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_10_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_10_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_10_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_10_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_10_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_10_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_10_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_10_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_10_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_10_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_10_ldst;	// rob.scala:310:28
  reg              rob_uop_2_10_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_10_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_10_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_11_uopc;	// rob.scala:310:28
  reg              rob_uop_2_11_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_11_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_11_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_11_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_11_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_11_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_11_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_11_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_11_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_11_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_11_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_11_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_11_ldst;	// rob.scala:310:28
  reg              rob_uop_2_11_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_11_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_11_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_12_uopc;	// rob.scala:310:28
  reg              rob_uop_2_12_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_12_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_12_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_12_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_12_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_12_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_12_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_12_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_12_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_12_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_12_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_12_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_12_ldst;	// rob.scala:310:28
  reg              rob_uop_2_12_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_12_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_12_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_13_uopc;	// rob.scala:310:28
  reg              rob_uop_2_13_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_13_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_13_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_13_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_13_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_13_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_13_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_13_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_13_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_13_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_13_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_13_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_13_ldst;	// rob.scala:310:28
  reg              rob_uop_2_13_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_13_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_13_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_14_uopc;	// rob.scala:310:28
  reg              rob_uop_2_14_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_14_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_14_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_14_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_14_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_14_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_14_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_14_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_14_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_14_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_14_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_14_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_14_ldst;	// rob.scala:310:28
  reg              rob_uop_2_14_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_14_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_14_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_15_uopc;	// rob.scala:310:28
  reg              rob_uop_2_15_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_15_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_15_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_15_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_15_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_15_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_15_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_15_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_15_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_15_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_15_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_15_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_15_ldst;	// rob.scala:310:28
  reg              rob_uop_2_15_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_15_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_15_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_16_uopc;	// rob.scala:310:28
  reg              rob_uop_2_16_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_16_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_16_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_16_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_16_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_16_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_16_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_16_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_16_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_16_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_16_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_16_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_16_ldst;	// rob.scala:310:28
  reg              rob_uop_2_16_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_16_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_16_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_17_uopc;	// rob.scala:310:28
  reg              rob_uop_2_17_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_17_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_17_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_17_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_17_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_17_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_17_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_17_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_17_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_17_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_17_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_17_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_17_ldst;	// rob.scala:310:28
  reg              rob_uop_2_17_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_17_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_17_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_18_uopc;	// rob.scala:310:28
  reg              rob_uop_2_18_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_18_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_18_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_18_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_18_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_18_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_18_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_18_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_18_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_18_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_18_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_18_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_18_ldst;	// rob.scala:310:28
  reg              rob_uop_2_18_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_18_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_18_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_19_uopc;	// rob.scala:310:28
  reg              rob_uop_2_19_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_19_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_19_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_19_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_19_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_19_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_19_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_19_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_19_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_19_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_19_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_19_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_19_ldst;	// rob.scala:310:28
  reg              rob_uop_2_19_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_19_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_19_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_20_uopc;	// rob.scala:310:28
  reg              rob_uop_2_20_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_20_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_20_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_20_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_20_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_20_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_20_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_20_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_20_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_20_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_20_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_20_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_20_ldst;	// rob.scala:310:28
  reg              rob_uop_2_20_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_20_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_20_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_21_uopc;	// rob.scala:310:28
  reg              rob_uop_2_21_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_21_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_21_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_21_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_21_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_21_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_21_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_21_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_21_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_21_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_21_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_21_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_21_ldst;	// rob.scala:310:28
  reg              rob_uop_2_21_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_21_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_21_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_22_uopc;	// rob.scala:310:28
  reg              rob_uop_2_22_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_22_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_22_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_22_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_22_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_22_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_22_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_22_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_22_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_22_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_22_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_22_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_22_ldst;	// rob.scala:310:28
  reg              rob_uop_2_22_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_22_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_22_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_23_uopc;	// rob.scala:310:28
  reg              rob_uop_2_23_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_23_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_23_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_23_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_23_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_23_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_23_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_23_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_23_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_23_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_23_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_23_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_23_ldst;	// rob.scala:310:28
  reg              rob_uop_2_23_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_23_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_23_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_24_uopc;	// rob.scala:310:28
  reg              rob_uop_2_24_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_24_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_24_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_24_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_24_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_24_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_24_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_24_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_24_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_24_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_24_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_24_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_24_ldst;	// rob.scala:310:28
  reg              rob_uop_2_24_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_24_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_24_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_25_uopc;	// rob.scala:310:28
  reg              rob_uop_2_25_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_25_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_25_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_25_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_25_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_25_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_25_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_25_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_25_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_25_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_25_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_25_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_25_ldst;	// rob.scala:310:28
  reg              rob_uop_2_25_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_25_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_25_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_26_uopc;	// rob.scala:310:28
  reg              rob_uop_2_26_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_26_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_26_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_26_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_26_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_26_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_26_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_26_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_26_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_26_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_26_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_26_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_26_ldst;	// rob.scala:310:28
  reg              rob_uop_2_26_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_26_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_26_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_27_uopc;	// rob.scala:310:28
  reg              rob_uop_2_27_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_27_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_27_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_27_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_27_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_27_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_27_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_27_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_27_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_27_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_27_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_27_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_27_ldst;	// rob.scala:310:28
  reg              rob_uop_2_27_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_27_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_27_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_28_uopc;	// rob.scala:310:28
  reg              rob_uop_2_28_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_28_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_28_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_28_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_28_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_28_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_28_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_28_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_28_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_28_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_28_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_28_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_28_ldst;	// rob.scala:310:28
  reg              rob_uop_2_28_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_28_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_28_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_29_uopc;	// rob.scala:310:28
  reg              rob_uop_2_29_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_29_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_29_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_29_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_29_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_29_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_29_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_29_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_29_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_29_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_29_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_29_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_29_ldst;	// rob.scala:310:28
  reg              rob_uop_2_29_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_29_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_29_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_30_uopc;	// rob.scala:310:28
  reg              rob_uop_2_30_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_30_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_30_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_30_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_30_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_30_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_30_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_30_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_30_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_30_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_30_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_30_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_30_ldst;	// rob.scala:310:28
  reg              rob_uop_2_30_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_30_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_30_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_31_uopc;	// rob.scala:310:28
  reg              rob_uop_2_31_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_2_31_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_31_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_31_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_31_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_31_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_31_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_31_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_31_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_31_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_31_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_31_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_31_ldst;	// rob.scala:310:28
  reg              rob_uop_2_31_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_31_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_31_fp_val;	// rob.scala:310:28
  reg              rob_exception_2_0;	// rob.scala:311:28
  reg              rob_exception_2_1;	// rob.scala:311:28
  reg              rob_exception_2_2;	// rob.scala:311:28
  reg              rob_exception_2_3;	// rob.scala:311:28
  reg              rob_exception_2_4;	// rob.scala:311:28
  reg              rob_exception_2_5;	// rob.scala:311:28
  reg              rob_exception_2_6;	// rob.scala:311:28
  reg              rob_exception_2_7;	// rob.scala:311:28
  reg              rob_exception_2_8;	// rob.scala:311:28
  reg              rob_exception_2_9;	// rob.scala:311:28
  reg              rob_exception_2_10;	// rob.scala:311:28
  reg              rob_exception_2_11;	// rob.scala:311:28
  reg              rob_exception_2_12;	// rob.scala:311:28
  reg              rob_exception_2_13;	// rob.scala:311:28
  reg              rob_exception_2_14;	// rob.scala:311:28
  reg              rob_exception_2_15;	// rob.scala:311:28
  reg              rob_exception_2_16;	// rob.scala:311:28
  reg              rob_exception_2_17;	// rob.scala:311:28
  reg              rob_exception_2_18;	// rob.scala:311:28
  reg              rob_exception_2_19;	// rob.scala:311:28
  reg              rob_exception_2_20;	// rob.scala:311:28
  reg              rob_exception_2_21;	// rob.scala:311:28
  reg              rob_exception_2_22;	// rob.scala:311:28
  reg              rob_exception_2_23;	// rob.scala:311:28
  reg              rob_exception_2_24;	// rob.scala:311:28
  reg              rob_exception_2_25;	// rob.scala:311:28
  reg              rob_exception_2_26;	// rob.scala:311:28
  reg              rob_exception_2_27;	// rob.scala:311:28
  reg              rob_exception_2_28;	// rob.scala:311:28
  reg              rob_exception_2_29;	// rob.scala:311:28
  reg              rob_exception_2_30;	// rob.scala:311:28
  reg              rob_exception_2_31;	// rob.scala:311:28
  reg              rob_predicated_2_0;	// rob.scala:312:29
  reg              rob_predicated_2_1;	// rob.scala:312:29
  reg              rob_predicated_2_2;	// rob.scala:312:29
  reg              rob_predicated_2_3;	// rob.scala:312:29
  reg              rob_predicated_2_4;	// rob.scala:312:29
  reg              rob_predicated_2_5;	// rob.scala:312:29
  reg              rob_predicated_2_6;	// rob.scala:312:29
  reg              rob_predicated_2_7;	// rob.scala:312:29
  reg              rob_predicated_2_8;	// rob.scala:312:29
  reg              rob_predicated_2_9;	// rob.scala:312:29
  reg              rob_predicated_2_10;	// rob.scala:312:29
  reg              rob_predicated_2_11;	// rob.scala:312:29
  reg              rob_predicated_2_12;	// rob.scala:312:29
  reg              rob_predicated_2_13;	// rob.scala:312:29
  reg              rob_predicated_2_14;	// rob.scala:312:29
  reg              rob_predicated_2_15;	// rob.scala:312:29
  reg              rob_predicated_2_16;	// rob.scala:312:29
  reg              rob_predicated_2_17;	// rob.scala:312:29
  reg              rob_predicated_2_18;	// rob.scala:312:29
  reg              rob_predicated_2_19;	// rob.scala:312:29
  reg              rob_predicated_2_20;	// rob.scala:312:29
  reg              rob_predicated_2_21;	// rob.scala:312:29
  reg              rob_predicated_2_22;	// rob.scala:312:29
  reg              rob_predicated_2_23;	// rob.scala:312:29
  reg              rob_predicated_2_24;	// rob.scala:312:29
  reg              rob_predicated_2_25;	// rob.scala:312:29
  reg              rob_predicated_2_26;	// rob.scala:312:29
  reg              rob_predicated_2_27;	// rob.scala:312:29
  reg              rob_predicated_2_28;	// rob.scala:312:29
  reg              rob_predicated_2_29;	// rob.scala:312:29
  reg              rob_predicated_2_30;	// rob.scala:312:29
  reg              rob_predicated_2_31;	// rob.scala:312:29
  wire [31:0]      _GEN_69 =
    {{rob_val_2_31},
     {rob_val_2_30},
     {rob_val_2_29},
     {rob_val_2_28},
     {rob_val_2_27},
     {rob_val_2_26},
     {rob_val_2_25},
     {rob_val_2_24},
     {rob_val_2_23},
     {rob_val_2_22},
     {rob_val_2_21},
     {rob_val_2_20},
     {rob_val_2_19},
     {rob_val_2_18},
     {rob_val_2_17},
     {rob_val_2_16},
     {rob_val_2_15},
     {rob_val_2_14},
     {rob_val_2_13},
     {rob_val_2_12},
     {rob_val_2_11},
     {rob_val_2_10},
     {rob_val_2_9},
     {rob_val_2_8},
     {rob_val_2_7},
     {rob_val_2_6},
     {rob_val_2_5},
     {rob_val_2_4},
     {rob_val_2_3},
     {rob_val_2_2},
     {rob_val_2_1},
     {rob_val_2_0}};	// rob.scala:307:32, :324:31
  wire             rob_tail_vals_2 = _GEN_69[rob_tail];	// rob.scala:228:29, :324:31
  wire             _GEN_70 =
    io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_71 =
    io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_72 =
    io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_73 =
    io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_74 =
    io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_75 =
    io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_76 =
    io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_77 =
    io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_78 =
    io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_79 =
    io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_80 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :361:31
  wire [31:0]      _GEN_81 =
    {{rob_bsy_2_31},
     {rob_bsy_2_30},
     {rob_bsy_2_29},
     {rob_bsy_2_28},
     {rob_bsy_2_27},
     {rob_bsy_2_26},
     {rob_bsy_2_25},
     {rob_bsy_2_24},
     {rob_bsy_2_23},
     {rob_bsy_2_22},
     {rob_bsy_2_21},
     {rob_bsy_2_20},
     {rob_bsy_2_19},
     {rob_bsy_2_18},
     {rob_bsy_2_17},
     {rob_bsy_2_16},
     {rob_bsy_2_15},
     {rob_bsy_2_14},
     {rob_bsy_2_13},
     {rob_bsy_2_12},
     {rob_bsy_2_11},
     {rob_bsy_2_10},
     {rob_bsy_2_9},
     {rob_bsy_2_8},
     {rob_bsy_2_7},
     {rob_bsy_2_6},
     {rob_bsy_2_5},
     {rob_bsy_2_4},
     {rob_bsy_2_3},
     {rob_bsy_2_2},
     {rob_bsy_2_1},
     {rob_bsy_2_0}};	// rob.scala:308:28, :366:31
  wire             _GEN_82 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :361:31
  wire             _GEN_83 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :361:31
  wire             _GEN_84 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :390:26
  wire [31:0]      _GEN_85 =
    {{rob_unsafe_2_31},
     {rob_unsafe_2_30},
     {rob_unsafe_2_29},
     {rob_unsafe_2_28},
     {rob_unsafe_2_27},
     {rob_unsafe_2_26},
     {rob_unsafe_2_25},
     {rob_unsafe_2_24},
     {rob_unsafe_2_23},
     {rob_unsafe_2_22},
     {rob_unsafe_2_21},
     {rob_unsafe_2_20},
     {rob_unsafe_2_19},
     {rob_unsafe_2_18},
     {rob_unsafe_2_17},
     {rob_unsafe_2_16},
     {rob_unsafe_2_15},
     {rob_unsafe_2_14},
     {rob_unsafe_2_13},
     {rob_unsafe_2_12},
     {rob_unsafe_2_11},
     {rob_unsafe_2_10},
     {rob_unsafe_2_9},
     {rob_unsafe_2_8},
     {rob_unsafe_2_7},
     {rob_unsafe_2_6},
     {rob_unsafe_2_5},
     {rob_unsafe_2_4},
     {rob_unsafe_2_3},
     {rob_unsafe_2_2},
     {rob_unsafe_2_1},
     {rob_unsafe_2_0}};	// rob.scala:309:28, :394:15
  wire             rob_head_vals_2 = _GEN_69[rob_head];	// rob.scala:224:29, :324:31, :398:49
  wire [31:0]      _GEN_86 =
    {{rob_exception_2_31},
     {rob_exception_2_30},
     {rob_exception_2_29},
     {rob_exception_2_28},
     {rob_exception_2_27},
     {rob_exception_2_26},
     {rob_exception_2_25},
     {rob_exception_2_24},
     {rob_exception_2_23},
     {rob_exception_2_22},
     {rob_exception_2_21},
     {rob_exception_2_20},
     {rob_exception_2_19},
     {rob_exception_2_18},
     {rob_exception_2_17},
     {rob_exception_2_16},
     {rob_exception_2_15},
     {rob_exception_2_14},
     {rob_exception_2_13},
     {rob_exception_2_12},
     {rob_exception_2_11},
     {rob_exception_2_10},
     {rob_exception_2_9},
     {rob_exception_2_8},
     {rob_exception_2_7},
     {rob_exception_2_6},
     {rob_exception_2_5},
     {rob_exception_2_4},
     {rob_exception_2_3},
     {rob_exception_2_2},
     {rob_exception_2_1},
     {rob_exception_2_0}};	// rob.scala:311:28, :398:49
  wire             can_throw_exception_2 = rob_head_vals_2 & _GEN_86[rob_head];	// rob.scala:224:29, :398:49
  wire             can_commit_2 = rob_head_vals_2 & ~_GEN_81[rob_head] & ~io_csr_stall;	// rob.scala:224:29, :366:31, :398:49, :404:{43,64,67}
  wire [31:0]      _GEN_87 =
    {{rob_predicated_2_31},
     {rob_predicated_2_30},
     {rob_predicated_2_29},
     {rob_predicated_2_28},
     {rob_predicated_2_27},
     {rob_predicated_2_26},
     {rob_predicated_2_25},
     {rob_predicated_2_24},
     {rob_predicated_2_23},
     {rob_predicated_2_22},
     {rob_predicated_2_21},
     {rob_predicated_2_20},
     {rob_predicated_2_19},
     {rob_predicated_2_18},
     {rob_predicated_2_17},
     {rob_predicated_2_16},
     {rob_predicated_2_15},
     {rob_predicated_2_14},
     {rob_predicated_2_13},
     {rob_predicated_2_12},
     {rob_predicated_2_11},
     {rob_predicated_2_10},
     {rob_predicated_2_9},
     {rob_predicated_2_8},
     {rob_predicated_2_7},
     {rob_predicated_2_6},
     {rob_predicated_2_5},
     {rob_predicated_2_4},
     {rob_predicated_2_3},
     {rob_predicated_2_2},
     {rob_predicated_2_1},
     {rob_predicated_2_0}};	// rob.scala:312:29, :410:51
  wire [31:0][6:0] _GEN_88 =
    {{rob_uop_2_31_uopc},
     {rob_uop_2_30_uopc},
     {rob_uop_2_29_uopc},
     {rob_uop_2_28_uopc},
     {rob_uop_2_27_uopc},
     {rob_uop_2_26_uopc},
     {rob_uop_2_25_uopc},
     {rob_uop_2_24_uopc},
     {rob_uop_2_23_uopc},
     {rob_uop_2_22_uopc},
     {rob_uop_2_21_uopc},
     {rob_uop_2_20_uopc},
     {rob_uop_2_19_uopc},
     {rob_uop_2_18_uopc},
     {rob_uop_2_17_uopc},
     {rob_uop_2_16_uopc},
     {rob_uop_2_15_uopc},
     {rob_uop_2_14_uopc},
     {rob_uop_2_13_uopc},
     {rob_uop_2_12_uopc},
     {rob_uop_2_11_uopc},
     {rob_uop_2_10_uopc},
     {rob_uop_2_9_uopc},
     {rob_uop_2_8_uopc},
     {rob_uop_2_7_uopc},
     {rob_uop_2_6_uopc},
     {rob_uop_2_5_uopc},
     {rob_uop_2_4_uopc},
     {rob_uop_2_3_uopc},
     {rob_uop_2_2_uopc},
     {rob_uop_2_1_uopc},
     {rob_uop_2_0_uopc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_89 =
    {{rob_uop_2_31_is_rvc},
     {rob_uop_2_30_is_rvc},
     {rob_uop_2_29_is_rvc},
     {rob_uop_2_28_is_rvc},
     {rob_uop_2_27_is_rvc},
     {rob_uop_2_26_is_rvc},
     {rob_uop_2_25_is_rvc},
     {rob_uop_2_24_is_rvc},
     {rob_uop_2_23_is_rvc},
     {rob_uop_2_22_is_rvc},
     {rob_uop_2_21_is_rvc},
     {rob_uop_2_20_is_rvc},
     {rob_uop_2_19_is_rvc},
     {rob_uop_2_18_is_rvc},
     {rob_uop_2_17_is_rvc},
     {rob_uop_2_16_is_rvc},
     {rob_uop_2_15_is_rvc},
     {rob_uop_2_14_is_rvc},
     {rob_uop_2_13_is_rvc},
     {rob_uop_2_12_is_rvc},
     {rob_uop_2_11_is_rvc},
     {rob_uop_2_10_is_rvc},
     {rob_uop_2_9_is_rvc},
     {rob_uop_2_8_is_rvc},
     {rob_uop_2_7_is_rvc},
     {rob_uop_2_6_is_rvc},
     {rob_uop_2_5_is_rvc},
     {rob_uop_2_4_is_rvc},
     {rob_uop_2_3_is_rvc},
     {rob_uop_2_2_is_rvc},
     {rob_uop_2_1_is_rvc},
     {rob_uop_2_0_is_rvc}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_90 =
    {{rob_uop_2_31_ftq_idx},
     {rob_uop_2_30_ftq_idx},
     {rob_uop_2_29_ftq_idx},
     {rob_uop_2_28_ftq_idx},
     {rob_uop_2_27_ftq_idx},
     {rob_uop_2_26_ftq_idx},
     {rob_uop_2_25_ftq_idx},
     {rob_uop_2_24_ftq_idx},
     {rob_uop_2_23_ftq_idx},
     {rob_uop_2_22_ftq_idx},
     {rob_uop_2_21_ftq_idx},
     {rob_uop_2_20_ftq_idx},
     {rob_uop_2_19_ftq_idx},
     {rob_uop_2_18_ftq_idx},
     {rob_uop_2_17_ftq_idx},
     {rob_uop_2_16_ftq_idx},
     {rob_uop_2_15_ftq_idx},
     {rob_uop_2_14_ftq_idx},
     {rob_uop_2_13_ftq_idx},
     {rob_uop_2_12_ftq_idx},
     {rob_uop_2_11_ftq_idx},
     {rob_uop_2_10_ftq_idx},
     {rob_uop_2_9_ftq_idx},
     {rob_uop_2_8_ftq_idx},
     {rob_uop_2_7_ftq_idx},
     {rob_uop_2_6_ftq_idx},
     {rob_uop_2_5_ftq_idx},
     {rob_uop_2_4_ftq_idx},
     {rob_uop_2_3_ftq_idx},
     {rob_uop_2_2_ftq_idx},
     {rob_uop_2_1_ftq_idx},
     {rob_uop_2_0_ftq_idx}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_91 =
    {{rob_uop_2_31_edge_inst},
     {rob_uop_2_30_edge_inst},
     {rob_uop_2_29_edge_inst},
     {rob_uop_2_28_edge_inst},
     {rob_uop_2_27_edge_inst},
     {rob_uop_2_26_edge_inst},
     {rob_uop_2_25_edge_inst},
     {rob_uop_2_24_edge_inst},
     {rob_uop_2_23_edge_inst},
     {rob_uop_2_22_edge_inst},
     {rob_uop_2_21_edge_inst},
     {rob_uop_2_20_edge_inst},
     {rob_uop_2_19_edge_inst},
     {rob_uop_2_18_edge_inst},
     {rob_uop_2_17_edge_inst},
     {rob_uop_2_16_edge_inst},
     {rob_uop_2_15_edge_inst},
     {rob_uop_2_14_edge_inst},
     {rob_uop_2_13_edge_inst},
     {rob_uop_2_12_edge_inst},
     {rob_uop_2_11_edge_inst},
     {rob_uop_2_10_edge_inst},
     {rob_uop_2_9_edge_inst},
     {rob_uop_2_8_edge_inst},
     {rob_uop_2_7_edge_inst},
     {rob_uop_2_6_edge_inst},
     {rob_uop_2_5_edge_inst},
     {rob_uop_2_4_edge_inst},
     {rob_uop_2_3_edge_inst},
     {rob_uop_2_2_edge_inst},
     {rob_uop_2_1_edge_inst},
     {rob_uop_2_0_edge_inst}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_92 =
    {{rob_uop_2_31_pc_lob},
     {rob_uop_2_30_pc_lob},
     {rob_uop_2_29_pc_lob},
     {rob_uop_2_28_pc_lob},
     {rob_uop_2_27_pc_lob},
     {rob_uop_2_26_pc_lob},
     {rob_uop_2_25_pc_lob},
     {rob_uop_2_24_pc_lob},
     {rob_uop_2_23_pc_lob},
     {rob_uop_2_22_pc_lob},
     {rob_uop_2_21_pc_lob},
     {rob_uop_2_20_pc_lob},
     {rob_uop_2_19_pc_lob},
     {rob_uop_2_18_pc_lob},
     {rob_uop_2_17_pc_lob},
     {rob_uop_2_16_pc_lob},
     {rob_uop_2_15_pc_lob},
     {rob_uop_2_14_pc_lob},
     {rob_uop_2_13_pc_lob},
     {rob_uop_2_12_pc_lob},
     {rob_uop_2_11_pc_lob},
     {rob_uop_2_10_pc_lob},
     {rob_uop_2_9_pc_lob},
     {rob_uop_2_8_pc_lob},
     {rob_uop_2_7_pc_lob},
     {rob_uop_2_6_pc_lob},
     {rob_uop_2_5_pc_lob},
     {rob_uop_2_4_pc_lob},
     {rob_uop_2_3_pc_lob},
     {rob_uop_2_2_pc_lob},
     {rob_uop_2_1_pc_lob},
     {rob_uop_2_0_pc_lob}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_93 =
    {{rob_uop_2_31_pdst},
     {rob_uop_2_30_pdst},
     {rob_uop_2_29_pdst},
     {rob_uop_2_28_pdst},
     {rob_uop_2_27_pdst},
     {rob_uop_2_26_pdst},
     {rob_uop_2_25_pdst},
     {rob_uop_2_24_pdst},
     {rob_uop_2_23_pdst},
     {rob_uop_2_22_pdst},
     {rob_uop_2_21_pdst},
     {rob_uop_2_20_pdst},
     {rob_uop_2_19_pdst},
     {rob_uop_2_18_pdst},
     {rob_uop_2_17_pdst},
     {rob_uop_2_16_pdst},
     {rob_uop_2_15_pdst},
     {rob_uop_2_14_pdst},
     {rob_uop_2_13_pdst},
     {rob_uop_2_12_pdst},
     {rob_uop_2_11_pdst},
     {rob_uop_2_10_pdst},
     {rob_uop_2_9_pdst},
     {rob_uop_2_8_pdst},
     {rob_uop_2_7_pdst},
     {rob_uop_2_6_pdst},
     {rob_uop_2_5_pdst},
     {rob_uop_2_4_pdst},
     {rob_uop_2_3_pdst},
     {rob_uop_2_2_pdst},
     {rob_uop_2_1_pdst},
     {rob_uop_2_0_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_94 =
    {{rob_uop_2_31_stale_pdst},
     {rob_uop_2_30_stale_pdst},
     {rob_uop_2_29_stale_pdst},
     {rob_uop_2_28_stale_pdst},
     {rob_uop_2_27_stale_pdst},
     {rob_uop_2_26_stale_pdst},
     {rob_uop_2_25_stale_pdst},
     {rob_uop_2_24_stale_pdst},
     {rob_uop_2_23_stale_pdst},
     {rob_uop_2_22_stale_pdst},
     {rob_uop_2_21_stale_pdst},
     {rob_uop_2_20_stale_pdst},
     {rob_uop_2_19_stale_pdst},
     {rob_uop_2_18_stale_pdst},
     {rob_uop_2_17_stale_pdst},
     {rob_uop_2_16_stale_pdst},
     {rob_uop_2_15_stale_pdst},
     {rob_uop_2_14_stale_pdst},
     {rob_uop_2_13_stale_pdst},
     {rob_uop_2_12_stale_pdst},
     {rob_uop_2_11_stale_pdst},
     {rob_uop_2_10_stale_pdst},
     {rob_uop_2_9_stale_pdst},
     {rob_uop_2_8_stale_pdst},
     {rob_uop_2_7_stale_pdst},
     {rob_uop_2_6_stale_pdst},
     {rob_uop_2_5_stale_pdst},
     {rob_uop_2_4_stale_pdst},
     {rob_uop_2_3_stale_pdst},
     {rob_uop_2_2_stale_pdst},
     {rob_uop_2_1_stale_pdst},
     {rob_uop_2_0_stale_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_95 =
    {{rob_uop_2_31_is_fencei},
     {rob_uop_2_30_is_fencei},
     {rob_uop_2_29_is_fencei},
     {rob_uop_2_28_is_fencei},
     {rob_uop_2_27_is_fencei},
     {rob_uop_2_26_is_fencei},
     {rob_uop_2_25_is_fencei},
     {rob_uop_2_24_is_fencei},
     {rob_uop_2_23_is_fencei},
     {rob_uop_2_22_is_fencei},
     {rob_uop_2_21_is_fencei},
     {rob_uop_2_20_is_fencei},
     {rob_uop_2_19_is_fencei},
     {rob_uop_2_18_is_fencei},
     {rob_uop_2_17_is_fencei},
     {rob_uop_2_16_is_fencei},
     {rob_uop_2_15_is_fencei},
     {rob_uop_2_14_is_fencei},
     {rob_uop_2_13_is_fencei},
     {rob_uop_2_12_is_fencei},
     {rob_uop_2_11_is_fencei},
     {rob_uop_2_10_is_fencei},
     {rob_uop_2_9_is_fencei},
     {rob_uop_2_8_is_fencei},
     {rob_uop_2_7_is_fencei},
     {rob_uop_2_6_is_fencei},
     {rob_uop_2_5_is_fencei},
     {rob_uop_2_4_is_fencei},
     {rob_uop_2_3_is_fencei},
     {rob_uop_2_2_is_fencei},
     {rob_uop_2_1_is_fencei},
     {rob_uop_2_0_is_fencei}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_96 =
    {{rob_uop_2_31_uses_ldq},
     {rob_uop_2_30_uses_ldq},
     {rob_uop_2_29_uses_ldq},
     {rob_uop_2_28_uses_ldq},
     {rob_uop_2_27_uses_ldq},
     {rob_uop_2_26_uses_ldq},
     {rob_uop_2_25_uses_ldq},
     {rob_uop_2_24_uses_ldq},
     {rob_uop_2_23_uses_ldq},
     {rob_uop_2_22_uses_ldq},
     {rob_uop_2_21_uses_ldq},
     {rob_uop_2_20_uses_ldq},
     {rob_uop_2_19_uses_ldq},
     {rob_uop_2_18_uses_ldq},
     {rob_uop_2_17_uses_ldq},
     {rob_uop_2_16_uses_ldq},
     {rob_uop_2_15_uses_ldq},
     {rob_uop_2_14_uses_ldq},
     {rob_uop_2_13_uses_ldq},
     {rob_uop_2_12_uses_ldq},
     {rob_uop_2_11_uses_ldq},
     {rob_uop_2_10_uses_ldq},
     {rob_uop_2_9_uses_ldq},
     {rob_uop_2_8_uses_ldq},
     {rob_uop_2_7_uses_ldq},
     {rob_uop_2_6_uses_ldq},
     {rob_uop_2_5_uses_ldq},
     {rob_uop_2_4_uses_ldq},
     {rob_uop_2_3_uses_ldq},
     {rob_uop_2_2_uses_ldq},
     {rob_uop_2_1_uses_ldq},
     {rob_uop_2_0_uses_ldq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_97 =
    {{rob_uop_2_31_uses_stq},
     {rob_uop_2_30_uses_stq},
     {rob_uop_2_29_uses_stq},
     {rob_uop_2_28_uses_stq},
     {rob_uop_2_27_uses_stq},
     {rob_uop_2_26_uses_stq},
     {rob_uop_2_25_uses_stq},
     {rob_uop_2_24_uses_stq},
     {rob_uop_2_23_uses_stq},
     {rob_uop_2_22_uses_stq},
     {rob_uop_2_21_uses_stq},
     {rob_uop_2_20_uses_stq},
     {rob_uop_2_19_uses_stq},
     {rob_uop_2_18_uses_stq},
     {rob_uop_2_17_uses_stq},
     {rob_uop_2_16_uses_stq},
     {rob_uop_2_15_uses_stq},
     {rob_uop_2_14_uses_stq},
     {rob_uop_2_13_uses_stq},
     {rob_uop_2_12_uses_stq},
     {rob_uop_2_11_uses_stq},
     {rob_uop_2_10_uses_stq},
     {rob_uop_2_9_uses_stq},
     {rob_uop_2_8_uses_stq},
     {rob_uop_2_7_uses_stq},
     {rob_uop_2_6_uses_stq},
     {rob_uop_2_5_uses_stq},
     {rob_uop_2_4_uses_stq},
     {rob_uop_2_3_uses_stq},
     {rob_uop_2_2_uses_stq},
     {rob_uop_2_1_uses_stq},
     {rob_uop_2_0_uses_stq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_98 =
    {{rob_uop_2_31_is_sys_pc2epc},
     {rob_uop_2_30_is_sys_pc2epc},
     {rob_uop_2_29_is_sys_pc2epc},
     {rob_uop_2_28_is_sys_pc2epc},
     {rob_uop_2_27_is_sys_pc2epc},
     {rob_uop_2_26_is_sys_pc2epc},
     {rob_uop_2_25_is_sys_pc2epc},
     {rob_uop_2_24_is_sys_pc2epc},
     {rob_uop_2_23_is_sys_pc2epc},
     {rob_uop_2_22_is_sys_pc2epc},
     {rob_uop_2_21_is_sys_pc2epc},
     {rob_uop_2_20_is_sys_pc2epc},
     {rob_uop_2_19_is_sys_pc2epc},
     {rob_uop_2_18_is_sys_pc2epc},
     {rob_uop_2_17_is_sys_pc2epc},
     {rob_uop_2_16_is_sys_pc2epc},
     {rob_uop_2_15_is_sys_pc2epc},
     {rob_uop_2_14_is_sys_pc2epc},
     {rob_uop_2_13_is_sys_pc2epc},
     {rob_uop_2_12_is_sys_pc2epc},
     {rob_uop_2_11_is_sys_pc2epc},
     {rob_uop_2_10_is_sys_pc2epc},
     {rob_uop_2_9_is_sys_pc2epc},
     {rob_uop_2_8_is_sys_pc2epc},
     {rob_uop_2_7_is_sys_pc2epc},
     {rob_uop_2_6_is_sys_pc2epc},
     {rob_uop_2_5_is_sys_pc2epc},
     {rob_uop_2_4_is_sys_pc2epc},
     {rob_uop_2_3_is_sys_pc2epc},
     {rob_uop_2_2_is_sys_pc2epc},
     {rob_uop_2_1_is_sys_pc2epc},
     {rob_uop_2_0_is_sys_pc2epc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_99 =
    {{rob_uop_2_31_flush_on_commit},
     {rob_uop_2_30_flush_on_commit},
     {rob_uop_2_29_flush_on_commit},
     {rob_uop_2_28_flush_on_commit},
     {rob_uop_2_27_flush_on_commit},
     {rob_uop_2_26_flush_on_commit},
     {rob_uop_2_25_flush_on_commit},
     {rob_uop_2_24_flush_on_commit},
     {rob_uop_2_23_flush_on_commit},
     {rob_uop_2_22_flush_on_commit},
     {rob_uop_2_21_flush_on_commit},
     {rob_uop_2_20_flush_on_commit},
     {rob_uop_2_19_flush_on_commit},
     {rob_uop_2_18_flush_on_commit},
     {rob_uop_2_17_flush_on_commit},
     {rob_uop_2_16_flush_on_commit},
     {rob_uop_2_15_flush_on_commit},
     {rob_uop_2_14_flush_on_commit},
     {rob_uop_2_13_flush_on_commit},
     {rob_uop_2_12_flush_on_commit},
     {rob_uop_2_11_flush_on_commit},
     {rob_uop_2_10_flush_on_commit},
     {rob_uop_2_9_flush_on_commit},
     {rob_uop_2_8_flush_on_commit},
     {rob_uop_2_7_flush_on_commit},
     {rob_uop_2_6_flush_on_commit},
     {rob_uop_2_5_flush_on_commit},
     {rob_uop_2_4_flush_on_commit},
     {rob_uop_2_3_flush_on_commit},
     {rob_uop_2_2_flush_on_commit},
     {rob_uop_2_1_flush_on_commit},
     {rob_uop_2_0_flush_on_commit}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_100 =
    {{rob_uop_2_31_ldst},
     {rob_uop_2_30_ldst},
     {rob_uop_2_29_ldst},
     {rob_uop_2_28_ldst},
     {rob_uop_2_27_ldst},
     {rob_uop_2_26_ldst},
     {rob_uop_2_25_ldst},
     {rob_uop_2_24_ldst},
     {rob_uop_2_23_ldst},
     {rob_uop_2_22_ldst},
     {rob_uop_2_21_ldst},
     {rob_uop_2_20_ldst},
     {rob_uop_2_19_ldst},
     {rob_uop_2_18_ldst},
     {rob_uop_2_17_ldst},
     {rob_uop_2_16_ldst},
     {rob_uop_2_15_ldst},
     {rob_uop_2_14_ldst},
     {rob_uop_2_13_ldst},
     {rob_uop_2_12_ldst},
     {rob_uop_2_11_ldst},
     {rob_uop_2_10_ldst},
     {rob_uop_2_9_ldst},
     {rob_uop_2_8_ldst},
     {rob_uop_2_7_ldst},
     {rob_uop_2_6_ldst},
     {rob_uop_2_5_ldst},
     {rob_uop_2_4_ldst},
     {rob_uop_2_3_ldst},
     {rob_uop_2_2_ldst},
     {rob_uop_2_1_ldst},
     {rob_uop_2_0_ldst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_101 =
    {{rob_uop_2_31_ldst_val},
     {rob_uop_2_30_ldst_val},
     {rob_uop_2_29_ldst_val},
     {rob_uop_2_28_ldst_val},
     {rob_uop_2_27_ldst_val},
     {rob_uop_2_26_ldst_val},
     {rob_uop_2_25_ldst_val},
     {rob_uop_2_24_ldst_val},
     {rob_uop_2_23_ldst_val},
     {rob_uop_2_22_ldst_val},
     {rob_uop_2_21_ldst_val},
     {rob_uop_2_20_ldst_val},
     {rob_uop_2_19_ldst_val},
     {rob_uop_2_18_ldst_val},
     {rob_uop_2_17_ldst_val},
     {rob_uop_2_16_ldst_val},
     {rob_uop_2_15_ldst_val},
     {rob_uop_2_14_ldst_val},
     {rob_uop_2_13_ldst_val},
     {rob_uop_2_12_ldst_val},
     {rob_uop_2_11_ldst_val},
     {rob_uop_2_10_ldst_val},
     {rob_uop_2_9_ldst_val},
     {rob_uop_2_8_ldst_val},
     {rob_uop_2_7_ldst_val},
     {rob_uop_2_6_ldst_val},
     {rob_uop_2_5_ldst_val},
     {rob_uop_2_4_ldst_val},
     {rob_uop_2_3_ldst_val},
     {rob_uop_2_2_ldst_val},
     {rob_uop_2_1_ldst_val},
     {rob_uop_2_0_ldst_val}};	// rob.scala:310:28, :411:25
  wire [31:0][1:0] _GEN_102 =
    {{rob_uop_2_31_dst_rtype},
     {rob_uop_2_30_dst_rtype},
     {rob_uop_2_29_dst_rtype},
     {rob_uop_2_28_dst_rtype},
     {rob_uop_2_27_dst_rtype},
     {rob_uop_2_26_dst_rtype},
     {rob_uop_2_25_dst_rtype},
     {rob_uop_2_24_dst_rtype},
     {rob_uop_2_23_dst_rtype},
     {rob_uop_2_22_dst_rtype},
     {rob_uop_2_21_dst_rtype},
     {rob_uop_2_20_dst_rtype},
     {rob_uop_2_19_dst_rtype},
     {rob_uop_2_18_dst_rtype},
     {rob_uop_2_17_dst_rtype},
     {rob_uop_2_16_dst_rtype},
     {rob_uop_2_15_dst_rtype},
     {rob_uop_2_14_dst_rtype},
     {rob_uop_2_13_dst_rtype},
     {rob_uop_2_12_dst_rtype},
     {rob_uop_2_11_dst_rtype},
     {rob_uop_2_10_dst_rtype},
     {rob_uop_2_9_dst_rtype},
     {rob_uop_2_8_dst_rtype},
     {rob_uop_2_7_dst_rtype},
     {rob_uop_2_6_dst_rtype},
     {rob_uop_2_5_dst_rtype},
     {rob_uop_2_4_dst_rtype},
     {rob_uop_2_3_dst_rtype},
     {rob_uop_2_2_dst_rtype},
     {rob_uop_2_1_dst_rtype},
     {rob_uop_2_0_dst_rtype}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_103 =
    {{rob_uop_2_31_fp_val},
     {rob_uop_2_30_fp_val},
     {rob_uop_2_29_fp_val},
     {rob_uop_2_28_fp_val},
     {rob_uop_2_27_fp_val},
     {rob_uop_2_26_fp_val},
     {rob_uop_2_25_fp_val},
     {rob_uop_2_24_fp_val},
     {rob_uop_2_23_fp_val},
     {rob_uop_2_22_fp_val},
     {rob_uop_2_21_fp_val},
     {rob_uop_2_20_fp_val},
     {rob_uop_2_19_fp_val},
     {rob_uop_2_18_fp_val},
     {rob_uop_2_17_fp_val},
     {rob_uop_2_16_fp_val},
     {rob_uop_2_15_fp_val},
     {rob_uop_2_14_fp_val},
     {rob_uop_2_13_fp_val},
     {rob_uop_2_12_fp_val},
     {rob_uop_2_11_fp_val},
     {rob_uop_2_10_fp_val},
     {rob_uop_2_9_fp_val},
     {rob_uop_2_8_fp_val},
     {rob_uop_2_7_fp_val},
     {rob_uop_2_6_fp_val},
     {rob_uop_2_5_fp_val},
     {rob_uop_2_4_fp_val},
     {rob_uop_2_3_fp_val},
     {rob_uop_2_2_fp_val},
     {rob_uop_2_1_fp_val},
     {rob_uop_2_0_fp_val}};	// rob.scala:310:28, :411:25
  wire             rbk_row_2 = _io_commit_rollback_T_3 & ~full;	// rob.scala:236:31, :425:{44,47}, :787:39
  wire             _io_commit_rbk_valids_2_output = rbk_row_2 & _GEN_69[com_idx];	// rob.scala:236:20, :324:31, :425:44, :427:40
  reg              rob_val_3_0;	// rob.scala:307:32
  reg              rob_val_3_1;	// rob.scala:307:32
  reg              rob_val_3_2;	// rob.scala:307:32
  reg              rob_val_3_3;	// rob.scala:307:32
  reg              rob_val_3_4;	// rob.scala:307:32
  reg              rob_val_3_5;	// rob.scala:307:32
  reg              rob_val_3_6;	// rob.scala:307:32
  reg              rob_val_3_7;	// rob.scala:307:32
  reg              rob_val_3_8;	// rob.scala:307:32
  reg              rob_val_3_9;	// rob.scala:307:32
  reg              rob_val_3_10;	// rob.scala:307:32
  reg              rob_val_3_11;	// rob.scala:307:32
  reg              rob_val_3_12;	// rob.scala:307:32
  reg              rob_val_3_13;	// rob.scala:307:32
  reg              rob_val_3_14;	// rob.scala:307:32
  reg              rob_val_3_15;	// rob.scala:307:32
  reg              rob_val_3_16;	// rob.scala:307:32
  reg              rob_val_3_17;	// rob.scala:307:32
  reg              rob_val_3_18;	// rob.scala:307:32
  reg              rob_val_3_19;	// rob.scala:307:32
  reg              rob_val_3_20;	// rob.scala:307:32
  reg              rob_val_3_21;	// rob.scala:307:32
  reg              rob_val_3_22;	// rob.scala:307:32
  reg              rob_val_3_23;	// rob.scala:307:32
  reg              rob_val_3_24;	// rob.scala:307:32
  reg              rob_val_3_25;	// rob.scala:307:32
  reg              rob_val_3_26;	// rob.scala:307:32
  reg              rob_val_3_27;	// rob.scala:307:32
  reg              rob_val_3_28;	// rob.scala:307:32
  reg              rob_val_3_29;	// rob.scala:307:32
  reg              rob_val_3_30;	// rob.scala:307:32
  reg              rob_val_3_31;	// rob.scala:307:32
  reg              rob_bsy_3_0;	// rob.scala:308:28
  reg              rob_bsy_3_1;	// rob.scala:308:28
  reg              rob_bsy_3_2;	// rob.scala:308:28
  reg              rob_bsy_3_3;	// rob.scala:308:28
  reg              rob_bsy_3_4;	// rob.scala:308:28
  reg              rob_bsy_3_5;	// rob.scala:308:28
  reg              rob_bsy_3_6;	// rob.scala:308:28
  reg              rob_bsy_3_7;	// rob.scala:308:28
  reg              rob_bsy_3_8;	// rob.scala:308:28
  reg              rob_bsy_3_9;	// rob.scala:308:28
  reg              rob_bsy_3_10;	// rob.scala:308:28
  reg              rob_bsy_3_11;	// rob.scala:308:28
  reg              rob_bsy_3_12;	// rob.scala:308:28
  reg              rob_bsy_3_13;	// rob.scala:308:28
  reg              rob_bsy_3_14;	// rob.scala:308:28
  reg              rob_bsy_3_15;	// rob.scala:308:28
  reg              rob_bsy_3_16;	// rob.scala:308:28
  reg              rob_bsy_3_17;	// rob.scala:308:28
  reg              rob_bsy_3_18;	// rob.scala:308:28
  reg              rob_bsy_3_19;	// rob.scala:308:28
  reg              rob_bsy_3_20;	// rob.scala:308:28
  reg              rob_bsy_3_21;	// rob.scala:308:28
  reg              rob_bsy_3_22;	// rob.scala:308:28
  reg              rob_bsy_3_23;	// rob.scala:308:28
  reg              rob_bsy_3_24;	// rob.scala:308:28
  reg              rob_bsy_3_25;	// rob.scala:308:28
  reg              rob_bsy_3_26;	// rob.scala:308:28
  reg              rob_bsy_3_27;	// rob.scala:308:28
  reg              rob_bsy_3_28;	// rob.scala:308:28
  reg              rob_bsy_3_29;	// rob.scala:308:28
  reg              rob_bsy_3_30;	// rob.scala:308:28
  reg              rob_bsy_3_31;	// rob.scala:308:28
  reg              rob_unsafe_3_0;	// rob.scala:309:28
  reg              rob_unsafe_3_1;	// rob.scala:309:28
  reg              rob_unsafe_3_2;	// rob.scala:309:28
  reg              rob_unsafe_3_3;	// rob.scala:309:28
  reg              rob_unsafe_3_4;	// rob.scala:309:28
  reg              rob_unsafe_3_5;	// rob.scala:309:28
  reg              rob_unsafe_3_6;	// rob.scala:309:28
  reg              rob_unsafe_3_7;	// rob.scala:309:28
  reg              rob_unsafe_3_8;	// rob.scala:309:28
  reg              rob_unsafe_3_9;	// rob.scala:309:28
  reg              rob_unsafe_3_10;	// rob.scala:309:28
  reg              rob_unsafe_3_11;	// rob.scala:309:28
  reg              rob_unsafe_3_12;	// rob.scala:309:28
  reg              rob_unsafe_3_13;	// rob.scala:309:28
  reg              rob_unsafe_3_14;	// rob.scala:309:28
  reg              rob_unsafe_3_15;	// rob.scala:309:28
  reg              rob_unsafe_3_16;	// rob.scala:309:28
  reg              rob_unsafe_3_17;	// rob.scala:309:28
  reg              rob_unsafe_3_18;	// rob.scala:309:28
  reg              rob_unsafe_3_19;	// rob.scala:309:28
  reg              rob_unsafe_3_20;	// rob.scala:309:28
  reg              rob_unsafe_3_21;	// rob.scala:309:28
  reg              rob_unsafe_3_22;	// rob.scala:309:28
  reg              rob_unsafe_3_23;	// rob.scala:309:28
  reg              rob_unsafe_3_24;	// rob.scala:309:28
  reg              rob_unsafe_3_25;	// rob.scala:309:28
  reg              rob_unsafe_3_26;	// rob.scala:309:28
  reg              rob_unsafe_3_27;	// rob.scala:309:28
  reg              rob_unsafe_3_28;	// rob.scala:309:28
  reg              rob_unsafe_3_29;	// rob.scala:309:28
  reg              rob_unsafe_3_30;	// rob.scala:309:28
  reg              rob_unsafe_3_31;	// rob.scala:309:28
  reg  [6:0]       rob_uop_3_0_uopc;	// rob.scala:310:28
  reg              rob_uop_3_0_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_0_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_0_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_0_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_0_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_0_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_0_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_0_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_0_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_0_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_0_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_0_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_0_ldst;	// rob.scala:310:28
  reg              rob_uop_3_0_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_0_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_0_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_1_uopc;	// rob.scala:310:28
  reg              rob_uop_3_1_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_1_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_1_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_1_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_1_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_1_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_1_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_1_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_1_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_1_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_1_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_1_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_1_ldst;	// rob.scala:310:28
  reg              rob_uop_3_1_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_1_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_1_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_2_uopc;	// rob.scala:310:28
  reg              rob_uop_3_2_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_2_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_2_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_2_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_2_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_2_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_2_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_2_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_2_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_2_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_2_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_2_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_2_ldst;	// rob.scala:310:28
  reg              rob_uop_3_2_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_2_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_2_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_3_uopc;	// rob.scala:310:28
  reg              rob_uop_3_3_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_3_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_3_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_3_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_3_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_3_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_3_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_3_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_3_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_3_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_3_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_3_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_3_ldst;	// rob.scala:310:28
  reg              rob_uop_3_3_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_3_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_3_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_4_uopc;	// rob.scala:310:28
  reg              rob_uop_3_4_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_4_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_4_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_4_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_4_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_4_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_4_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_4_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_4_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_4_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_4_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_4_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_4_ldst;	// rob.scala:310:28
  reg              rob_uop_3_4_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_4_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_4_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_5_uopc;	// rob.scala:310:28
  reg              rob_uop_3_5_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_5_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_5_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_5_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_5_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_5_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_5_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_5_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_5_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_5_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_5_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_5_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_5_ldst;	// rob.scala:310:28
  reg              rob_uop_3_5_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_5_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_5_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_6_uopc;	// rob.scala:310:28
  reg              rob_uop_3_6_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_6_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_6_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_6_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_6_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_6_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_6_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_6_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_6_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_6_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_6_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_6_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_6_ldst;	// rob.scala:310:28
  reg              rob_uop_3_6_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_6_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_6_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_7_uopc;	// rob.scala:310:28
  reg              rob_uop_3_7_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_7_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_7_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_7_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_7_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_7_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_7_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_7_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_7_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_7_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_7_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_7_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_7_ldst;	// rob.scala:310:28
  reg              rob_uop_3_7_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_7_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_7_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_8_uopc;	// rob.scala:310:28
  reg              rob_uop_3_8_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_8_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_8_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_8_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_8_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_8_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_8_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_8_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_8_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_8_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_8_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_8_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_8_ldst;	// rob.scala:310:28
  reg              rob_uop_3_8_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_8_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_8_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_9_uopc;	// rob.scala:310:28
  reg              rob_uop_3_9_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_9_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_9_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_9_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_9_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_9_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_9_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_9_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_9_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_9_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_9_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_9_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_9_ldst;	// rob.scala:310:28
  reg              rob_uop_3_9_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_9_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_9_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_10_uopc;	// rob.scala:310:28
  reg              rob_uop_3_10_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_10_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_10_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_10_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_10_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_10_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_10_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_10_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_10_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_10_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_10_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_10_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_10_ldst;	// rob.scala:310:28
  reg              rob_uop_3_10_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_10_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_10_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_11_uopc;	// rob.scala:310:28
  reg              rob_uop_3_11_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_11_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_11_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_11_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_11_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_11_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_11_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_11_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_11_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_11_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_11_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_11_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_11_ldst;	// rob.scala:310:28
  reg              rob_uop_3_11_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_11_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_11_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_12_uopc;	// rob.scala:310:28
  reg              rob_uop_3_12_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_12_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_12_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_12_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_12_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_12_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_12_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_12_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_12_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_12_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_12_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_12_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_12_ldst;	// rob.scala:310:28
  reg              rob_uop_3_12_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_12_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_12_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_13_uopc;	// rob.scala:310:28
  reg              rob_uop_3_13_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_13_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_13_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_13_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_13_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_13_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_13_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_13_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_13_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_13_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_13_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_13_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_13_ldst;	// rob.scala:310:28
  reg              rob_uop_3_13_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_13_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_13_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_14_uopc;	// rob.scala:310:28
  reg              rob_uop_3_14_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_14_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_14_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_14_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_14_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_14_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_14_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_14_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_14_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_14_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_14_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_14_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_14_ldst;	// rob.scala:310:28
  reg              rob_uop_3_14_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_14_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_14_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_15_uopc;	// rob.scala:310:28
  reg              rob_uop_3_15_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_15_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_15_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_15_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_15_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_15_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_15_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_15_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_15_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_15_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_15_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_15_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_15_ldst;	// rob.scala:310:28
  reg              rob_uop_3_15_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_15_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_15_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_16_uopc;	// rob.scala:310:28
  reg              rob_uop_3_16_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_16_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_16_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_16_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_16_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_16_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_16_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_16_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_16_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_16_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_16_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_16_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_16_ldst;	// rob.scala:310:28
  reg              rob_uop_3_16_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_16_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_16_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_17_uopc;	// rob.scala:310:28
  reg              rob_uop_3_17_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_17_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_17_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_17_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_17_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_17_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_17_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_17_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_17_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_17_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_17_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_17_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_17_ldst;	// rob.scala:310:28
  reg              rob_uop_3_17_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_17_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_17_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_18_uopc;	// rob.scala:310:28
  reg              rob_uop_3_18_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_18_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_18_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_18_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_18_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_18_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_18_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_18_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_18_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_18_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_18_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_18_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_18_ldst;	// rob.scala:310:28
  reg              rob_uop_3_18_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_18_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_18_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_19_uopc;	// rob.scala:310:28
  reg              rob_uop_3_19_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_19_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_19_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_19_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_19_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_19_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_19_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_19_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_19_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_19_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_19_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_19_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_19_ldst;	// rob.scala:310:28
  reg              rob_uop_3_19_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_19_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_19_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_20_uopc;	// rob.scala:310:28
  reg              rob_uop_3_20_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_20_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_20_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_20_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_20_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_20_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_20_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_20_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_20_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_20_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_20_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_20_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_20_ldst;	// rob.scala:310:28
  reg              rob_uop_3_20_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_20_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_20_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_21_uopc;	// rob.scala:310:28
  reg              rob_uop_3_21_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_21_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_21_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_21_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_21_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_21_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_21_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_21_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_21_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_21_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_21_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_21_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_21_ldst;	// rob.scala:310:28
  reg              rob_uop_3_21_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_21_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_21_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_22_uopc;	// rob.scala:310:28
  reg              rob_uop_3_22_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_22_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_22_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_22_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_22_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_22_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_22_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_22_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_22_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_22_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_22_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_22_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_22_ldst;	// rob.scala:310:28
  reg              rob_uop_3_22_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_22_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_22_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_23_uopc;	// rob.scala:310:28
  reg              rob_uop_3_23_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_23_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_23_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_23_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_23_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_23_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_23_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_23_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_23_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_23_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_23_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_23_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_23_ldst;	// rob.scala:310:28
  reg              rob_uop_3_23_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_23_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_23_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_24_uopc;	// rob.scala:310:28
  reg              rob_uop_3_24_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_24_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_24_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_24_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_24_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_24_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_24_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_24_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_24_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_24_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_24_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_24_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_24_ldst;	// rob.scala:310:28
  reg              rob_uop_3_24_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_24_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_24_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_25_uopc;	// rob.scala:310:28
  reg              rob_uop_3_25_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_25_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_25_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_25_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_25_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_25_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_25_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_25_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_25_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_25_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_25_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_25_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_25_ldst;	// rob.scala:310:28
  reg              rob_uop_3_25_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_25_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_25_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_26_uopc;	// rob.scala:310:28
  reg              rob_uop_3_26_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_26_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_26_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_26_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_26_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_26_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_26_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_26_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_26_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_26_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_26_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_26_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_26_ldst;	// rob.scala:310:28
  reg              rob_uop_3_26_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_26_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_26_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_27_uopc;	// rob.scala:310:28
  reg              rob_uop_3_27_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_27_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_27_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_27_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_27_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_27_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_27_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_27_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_27_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_27_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_27_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_27_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_27_ldst;	// rob.scala:310:28
  reg              rob_uop_3_27_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_27_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_27_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_28_uopc;	// rob.scala:310:28
  reg              rob_uop_3_28_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_28_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_28_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_28_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_28_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_28_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_28_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_28_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_28_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_28_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_28_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_28_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_28_ldst;	// rob.scala:310:28
  reg              rob_uop_3_28_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_28_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_28_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_29_uopc;	// rob.scala:310:28
  reg              rob_uop_3_29_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_29_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_29_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_29_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_29_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_29_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_29_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_29_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_29_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_29_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_29_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_29_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_29_ldst;	// rob.scala:310:28
  reg              rob_uop_3_29_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_29_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_29_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_30_uopc;	// rob.scala:310:28
  reg              rob_uop_3_30_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_30_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_30_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_30_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_30_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_30_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_30_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_30_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_30_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_30_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_30_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_30_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_30_ldst;	// rob.scala:310:28
  reg              rob_uop_3_30_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_30_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_30_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_31_uopc;	// rob.scala:310:28
  reg              rob_uop_3_31_is_rvc;	// rob.scala:310:28
  reg  [19:0]      rob_uop_3_31_br_mask;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_31_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_31_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_31_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_31_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_31_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_31_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_31_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_31_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_31_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_31_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_31_ldst;	// rob.scala:310:28
  reg              rob_uop_3_31_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_31_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_31_fp_val;	// rob.scala:310:28
  reg              rob_exception_3_0;	// rob.scala:311:28
  reg              rob_exception_3_1;	// rob.scala:311:28
  reg              rob_exception_3_2;	// rob.scala:311:28
  reg              rob_exception_3_3;	// rob.scala:311:28
  reg              rob_exception_3_4;	// rob.scala:311:28
  reg              rob_exception_3_5;	// rob.scala:311:28
  reg              rob_exception_3_6;	// rob.scala:311:28
  reg              rob_exception_3_7;	// rob.scala:311:28
  reg              rob_exception_3_8;	// rob.scala:311:28
  reg              rob_exception_3_9;	// rob.scala:311:28
  reg              rob_exception_3_10;	// rob.scala:311:28
  reg              rob_exception_3_11;	// rob.scala:311:28
  reg              rob_exception_3_12;	// rob.scala:311:28
  reg              rob_exception_3_13;	// rob.scala:311:28
  reg              rob_exception_3_14;	// rob.scala:311:28
  reg              rob_exception_3_15;	// rob.scala:311:28
  reg              rob_exception_3_16;	// rob.scala:311:28
  reg              rob_exception_3_17;	// rob.scala:311:28
  reg              rob_exception_3_18;	// rob.scala:311:28
  reg              rob_exception_3_19;	// rob.scala:311:28
  reg              rob_exception_3_20;	// rob.scala:311:28
  reg              rob_exception_3_21;	// rob.scala:311:28
  reg              rob_exception_3_22;	// rob.scala:311:28
  reg              rob_exception_3_23;	// rob.scala:311:28
  reg              rob_exception_3_24;	// rob.scala:311:28
  reg              rob_exception_3_25;	// rob.scala:311:28
  reg              rob_exception_3_26;	// rob.scala:311:28
  reg              rob_exception_3_27;	// rob.scala:311:28
  reg              rob_exception_3_28;	// rob.scala:311:28
  reg              rob_exception_3_29;	// rob.scala:311:28
  reg              rob_exception_3_30;	// rob.scala:311:28
  reg              rob_exception_3_31;	// rob.scala:311:28
  reg              rob_predicated_3_0;	// rob.scala:312:29
  reg              rob_predicated_3_1;	// rob.scala:312:29
  reg              rob_predicated_3_2;	// rob.scala:312:29
  reg              rob_predicated_3_3;	// rob.scala:312:29
  reg              rob_predicated_3_4;	// rob.scala:312:29
  reg              rob_predicated_3_5;	// rob.scala:312:29
  reg              rob_predicated_3_6;	// rob.scala:312:29
  reg              rob_predicated_3_7;	// rob.scala:312:29
  reg              rob_predicated_3_8;	// rob.scala:312:29
  reg              rob_predicated_3_9;	// rob.scala:312:29
  reg              rob_predicated_3_10;	// rob.scala:312:29
  reg              rob_predicated_3_11;	// rob.scala:312:29
  reg              rob_predicated_3_12;	// rob.scala:312:29
  reg              rob_predicated_3_13;	// rob.scala:312:29
  reg              rob_predicated_3_14;	// rob.scala:312:29
  reg              rob_predicated_3_15;	// rob.scala:312:29
  reg              rob_predicated_3_16;	// rob.scala:312:29
  reg              rob_predicated_3_17;	// rob.scala:312:29
  reg              rob_predicated_3_18;	// rob.scala:312:29
  reg              rob_predicated_3_19;	// rob.scala:312:29
  reg              rob_predicated_3_20;	// rob.scala:312:29
  reg              rob_predicated_3_21;	// rob.scala:312:29
  reg              rob_predicated_3_22;	// rob.scala:312:29
  reg              rob_predicated_3_23;	// rob.scala:312:29
  reg              rob_predicated_3_24;	// rob.scala:312:29
  reg              rob_predicated_3_25;	// rob.scala:312:29
  reg              rob_predicated_3_26;	// rob.scala:312:29
  reg              rob_predicated_3_27;	// rob.scala:312:29
  reg              rob_predicated_3_28;	// rob.scala:312:29
  reg              rob_predicated_3_29;	// rob.scala:312:29
  reg              rob_predicated_3_30;	// rob.scala:312:29
  reg              rob_predicated_3_31;	// rob.scala:312:29
  wire [31:0]      _GEN_104 =
    {{rob_val_3_31},
     {rob_val_3_30},
     {rob_val_3_29},
     {rob_val_3_28},
     {rob_val_3_27},
     {rob_val_3_26},
     {rob_val_3_25},
     {rob_val_3_24},
     {rob_val_3_23},
     {rob_val_3_22},
     {rob_val_3_21},
     {rob_val_3_20},
     {rob_val_3_19},
     {rob_val_3_18},
     {rob_val_3_17},
     {rob_val_3_16},
     {rob_val_3_15},
     {rob_val_3_14},
     {rob_val_3_13},
     {rob_val_3_12},
     {rob_val_3_11},
     {rob_val_3_10},
     {rob_val_3_9},
     {rob_val_3_8},
     {rob_val_3_7},
     {rob_val_3_6},
     {rob_val_3_5},
     {rob_val_3_4},
     {rob_val_3_3},
     {rob_val_3_2},
     {rob_val_3_1},
     {rob_val_3_0}};	// rob.scala:307:32, :324:31
  wire             rob_tail_vals_3 = _GEN_104[rob_tail];	// rob.scala:228:29, :324:31
  wire             _GEN_105 =
    io_wb_resps_0_valid & (&(io_wb_resps_0_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_106 =
    io_wb_resps_1_valid & (&(io_wb_resps_1_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_107 =
    io_wb_resps_2_valid & (&(io_wb_resps_2_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_108 =
    io_wb_resps_3_valid & (&(io_wb_resps_3_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_109 =
    io_wb_resps_4_valid & (&(io_wb_resps_4_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_110 =
    io_wb_resps_5_valid & (&(io_wb_resps_5_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_111 =
    io_wb_resps_6_valid & (&(io_wb_resps_6_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_112 =
    io_wb_resps_7_valid & (&(io_wb_resps_7_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_113 =
    io_wb_resps_8_valid & (&(io_wb_resps_8_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_114 =
    io_wb_resps_9_valid & (&(io_wb_resps_9_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :346:27
  wire             _GEN_115 = io_lsu_clr_bsy_0_valid & (&(io_lsu_clr_bsy_0_bits[1:0]));	// rob.scala:272:36, :304:53, :361:31
  wire [31:0]      _GEN_116 =
    {{rob_bsy_3_31},
     {rob_bsy_3_30},
     {rob_bsy_3_29},
     {rob_bsy_3_28},
     {rob_bsy_3_27},
     {rob_bsy_3_26},
     {rob_bsy_3_25},
     {rob_bsy_3_24},
     {rob_bsy_3_23},
     {rob_bsy_3_22},
     {rob_bsy_3_21},
     {rob_bsy_3_20},
     {rob_bsy_3_19},
     {rob_bsy_3_18},
     {rob_bsy_3_17},
     {rob_bsy_3_16},
     {rob_bsy_3_15},
     {rob_bsy_3_14},
     {rob_bsy_3_13},
     {rob_bsy_3_12},
     {rob_bsy_3_11},
     {rob_bsy_3_10},
     {rob_bsy_3_9},
     {rob_bsy_3_8},
     {rob_bsy_3_7},
     {rob_bsy_3_6},
     {rob_bsy_3_5},
     {rob_bsy_3_4},
     {rob_bsy_3_3},
     {rob_bsy_3_2},
     {rob_bsy_3_1},
     {rob_bsy_3_0}};	// rob.scala:308:28, :366:31
  wire             _GEN_117 = io_lsu_clr_bsy_1_valid & (&(io_lsu_clr_bsy_1_bits[1:0]));	// rob.scala:272:36, :304:53, :361:31
  wire             _GEN_118 = io_lsu_clr_bsy_2_valid & (&(io_lsu_clr_bsy_2_bits[1:0]));	// rob.scala:272:36, :304:53, :361:31
  wire             _GEN_119 = io_lxcpt_valid & (&(io_lxcpt_bits_uop_rob_idx[1:0]));	// rob.scala:272:36, :304:53, :390:26
  wire [31:0]      _GEN_120 =
    {{rob_unsafe_3_31},
     {rob_unsafe_3_30},
     {rob_unsafe_3_29},
     {rob_unsafe_3_28},
     {rob_unsafe_3_27},
     {rob_unsafe_3_26},
     {rob_unsafe_3_25},
     {rob_unsafe_3_24},
     {rob_unsafe_3_23},
     {rob_unsafe_3_22},
     {rob_unsafe_3_21},
     {rob_unsafe_3_20},
     {rob_unsafe_3_19},
     {rob_unsafe_3_18},
     {rob_unsafe_3_17},
     {rob_unsafe_3_16},
     {rob_unsafe_3_15},
     {rob_unsafe_3_14},
     {rob_unsafe_3_13},
     {rob_unsafe_3_12},
     {rob_unsafe_3_11},
     {rob_unsafe_3_10},
     {rob_unsafe_3_9},
     {rob_unsafe_3_8},
     {rob_unsafe_3_7},
     {rob_unsafe_3_6},
     {rob_unsafe_3_5},
     {rob_unsafe_3_4},
     {rob_unsafe_3_3},
     {rob_unsafe_3_2},
     {rob_unsafe_3_1},
     {rob_unsafe_3_0}};	// rob.scala:309:28, :394:15
  wire             rob_head_vals_3 = _GEN_104[rob_head];	// rob.scala:224:29, :324:31, :398:49
  wire [31:0]      _GEN_121 =
    {{rob_exception_3_31},
     {rob_exception_3_30},
     {rob_exception_3_29},
     {rob_exception_3_28},
     {rob_exception_3_27},
     {rob_exception_3_26},
     {rob_exception_3_25},
     {rob_exception_3_24},
     {rob_exception_3_23},
     {rob_exception_3_22},
     {rob_exception_3_21},
     {rob_exception_3_20},
     {rob_exception_3_19},
     {rob_exception_3_18},
     {rob_exception_3_17},
     {rob_exception_3_16},
     {rob_exception_3_15},
     {rob_exception_3_14},
     {rob_exception_3_13},
     {rob_exception_3_12},
     {rob_exception_3_11},
     {rob_exception_3_10},
     {rob_exception_3_9},
     {rob_exception_3_8},
     {rob_exception_3_7},
     {rob_exception_3_6},
     {rob_exception_3_5},
     {rob_exception_3_4},
     {rob_exception_3_3},
     {rob_exception_3_2},
     {rob_exception_3_1},
     {rob_exception_3_0}};	// rob.scala:311:28, :398:49
  wire             can_throw_exception_3 = rob_head_vals_3 & _GEN_121[rob_head];	// rob.scala:224:29, :398:49
  wire [31:0]      _GEN_122 =
    {{rob_predicated_3_31},
     {rob_predicated_3_30},
     {rob_predicated_3_29},
     {rob_predicated_3_28},
     {rob_predicated_3_27},
     {rob_predicated_3_26},
     {rob_predicated_3_25},
     {rob_predicated_3_24},
     {rob_predicated_3_23},
     {rob_predicated_3_22},
     {rob_predicated_3_21},
     {rob_predicated_3_20},
     {rob_predicated_3_19},
     {rob_predicated_3_18},
     {rob_predicated_3_17},
     {rob_predicated_3_16},
     {rob_predicated_3_15},
     {rob_predicated_3_14},
     {rob_predicated_3_13},
     {rob_predicated_3_12},
     {rob_predicated_3_11},
     {rob_predicated_3_10},
     {rob_predicated_3_9},
     {rob_predicated_3_8},
     {rob_predicated_3_7},
     {rob_predicated_3_6},
     {rob_predicated_3_5},
     {rob_predicated_3_4},
     {rob_predicated_3_3},
     {rob_predicated_3_2},
     {rob_predicated_3_1},
     {rob_predicated_3_0}};	// rob.scala:312:29, :410:51
  wire [31:0][6:0] _GEN_123 =
    {{rob_uop_3_31_uopc},
     {rob_uop_3_30_uopc},
     {rob_uop_3_29_uopc},
     {rob_uop_3_28_uopc},
     {rob_uop_3_27_uopc},
     {rob_uop_3_26_uopc},
     {rob_uop_3_25_uopc},
     {rob_uop_3_24_uopc},
     {rob_uop_3_23_uopc},
     {rob_uop_3_22_uopc},
     {rob_uop_3_21_uopc},
     {rob_uop_3_20_uopc},
     {rob_uop_3_19_uopc},
     {rob_uop_3_18_uopc},
     {rob_uop_3_17_uopc},
     {rob_uop_3_16_uopc},
     {rob_uop_3_15_uopc},
     {rob_uop_3_14_uopc},
     {rob_uop_3_13_uopc},
     {rob_uop_3_12_uopc},
     {rob_uop_3_11_uopc},
     {rob_uop_3_10_uopc},
     {rob_uop_3_9_uopc},
     {rob_uop_3_8_uopc},
     {rob_uop_3_7_uopc},
     {rob_uop_3_6_uopc},
     {rob_uop_3_5_uopc},
     {rob_uop_3_4_uopc},
     {rob_uop_3_3_uopc},
     {rob_uop_3_2_uopc},
     {rob_uop_3_1_uopc},
     {rob_uop_3_0_uopc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_124 =
    {{rob_uop_3_31_is_rvc},
     {rob_uop_3_30_is_rvc},
     {rob_uop_3_29_is_rvc},
     {rob_uop_3_28_is_rvc},
     {rob_uop_3_27_is_rvc},
     {rob_uop_3_26_is_rvc},
     {rob_uop_3_25_is_rvc},
     {rob_uop_3_24_is_rvc},
     {rob_uop_3_23_is_rvc},
     {rob_uop_3_22_is_rvc},
     {rob_uop_3_21_is_rvc},
     {rob_uop_3_20_is_rvc},
     {rob_uop_3_19_is_rvc},
     {rob_uop_3_18_is_rvc},
     {rob_uop_3_17_is_rvc},
     {rob_uop_3_16_is_rvc},
     {rob_uop_3_15_is_rvc},
     {rob_uop_3_14_is_rvc},
     {rob_uop_3_13_is_rvc},
     {rob_uop_3_12_is_rvc},
     {rob_uop_3_11_is_rvc},
     {rob_uop_3_10_is_rvc},
     {rob_uop_3_9_is_rvc},
     {rob_uop_3_8_is_rvc},
     {rob_uop_3_7_is_rvc},
     {rob_uop_3_6_is_rvc},
     {rob_uop_3_5_is_rvc},
     {rob_uop_3_4_is_rvc},
     {rob_uop_3_3_is_rvc},
     {rob_uop_3_2_is_rvc},
     {rob_uop_3_1_is_rvc},
     {rob_uop_3_0_is_rvc}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_125 =
    {{rob_uop_3_31_ftq_idx},
     {rob_uop_3_30_ftq_idx},
     {rob_uop_3_29_ftq_idx},
     {rob_uop_3_28_ftq_idx},
     {rob_uop_3_27_ftq_idx},
     {rob_uop_3_26_ftq_idx},
     {rob_uop_3_25_ftq_idx},
     {rob_uop_3_24_ftq_idx},
     {rob_uop_3_23_ftq_idx},
     {rob_uop_3_22_ftq_idx},
     {rob_uop_3_21_ftq_idx},
     {rob_uop_3_20_ftq_idx},
     {rob_uop_3_19_ftq_idx},
     {rob_uop_3_18_ftq_idx},
     {rob_uop_3_17_ftq_idx},
     {rob_uop_3_16_ftq_idx},
     {rob_uop_3_15_ftq_idx},
     {rob_uop_3_14_ftq_idx},
     {rob_uop_3_13_ftq_idx},
     {rob_uop_3_12_ftq_idx},
     {rob_uop_3_11_ftq_idx},
     {rob_uop_3_10_ftq_idx},
     {rob_uop_3_9_ftq_idx},
     {rob_uop_3_8_ftq_idx},
     {rob_uop_3_7_ftq_idx},
     {rob_uop_3_6_ftq_idx},
     {rob_uop_3_5_ftq_idx},
     {rob_uop_3_4_ftq_idx},
     {rob_uop_3_3_ftq_idx},
     {rob_uop_3_2_ftq_idx},
     {rob_uop_3_1_ftq_idx},
     {rob_uop_3_0_ftq_idx}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_126 =
    {{rob_uop_3_31_edge_inst},
     {rob_uop_3_30_edge_inst},
     {rob_uop_3_29_edge_inst},
     {rob_uop_3_28_edge_inst},
     {rob_uop_3_27_edge_inst},
     {rob_uop_3_26_edge_inst},
     {rob_uop_3_25_edge_inst},
     {rob_uop_3_24_edge_inst},
     {rob_uop_3_23_edge_inst},
     {rob_uop_3_22_edge_inst},
     {rob_uop_3_21_edge_inst},
     {rob_uop_3_20_edge_inst},
     {rob_uop_3_19_edge_inst},
     {rob_uop_3_18_edge_inst},
     {rob_uop_3_17_edge_inst},
     {rob_uop_3_16_edge_inst},
     {rob_uop_3_15_edge_inst},
     {rob_uop_3_14_edge_inst},
     {rob_uop_3_13_edge_inst},
     {rob_uop_3_12_edge_inst},
     {rob_uop_3_11_edge_inst},
     {rob_uop_3_10_edge_inst},
     {rob_uop_3_9_edge_inst},
     {rob_uop_3_8_edge_inst},
     {rob_uop_3_7_edge_inst},
     {rob_uop_3_6_edge_inst},
     {rob_uop_3_5_edge_inst},
     {rob_uop_3_4_edge_inst},
     {rob_uop_3_3_edge_inst},
     {rob_uop_3_2_edge_inst},
     {rob_uop_3_1_edge_inst},
     {rob_uop_3_0_edge_inst}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_127 =
    {{rob_uop_3_31_pc_lob},
     {rob_uop_3_30_pc_lob},
     {rob_uop_3_29_pc_lob},
     {rob_uop_3_28_pc_lob},
     {rob_uop_3_27_pc_lob},
     {rob_uop_3_26_pc_lob},
     {rob_uop_3_25_pc_lob},
     {rob_uop_3_24_pc_lob},
     {rob_uop_3_23_pc_lob},
     {rob_uop_3_22_pc_lob},
     {rob_uop_3_21_pc_lob},
     {rob_uop_3_20_pc_lob},
     {rob_uop_3_19_pc_lob},
     {rob_uop_3_18_pc_lob},
     {rob_uop_3_17_pc_lob},
     {rob_uop_3_16_pc_lob},
     {rob_uop_3_15_pc_lob},
     {rob_uop_3_14_pc_lob},
     {rob_uop_3_13_pc_lob},
     {rob_uop_3_12_pc_lob},
     {rob_uop_3_11_pc_lob},
     {rob_uop_3_10_pc_lob},
     {rob_uop_3_9_pc_lob},
     {rob_uop_3_8_pc_lob},
     {rob_uop_3_7_pc_lob},
     {rob_uop_3_6_pc_lob},
     {rob_uop_3_5_pc_lob},
     {rob_uop_3_4_pc_lob},
     {rob_uop_3_3_pc_lob},
     {rob_uop_3_2_pc_lob},
     {rob_uop_3_1_pc_lob},
     {rob_uop_3_0_pc_lob}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_128 =
    {{rob_uop_3_31_pdst},
     {rob_uop_3_30_pdst},
     {rob_uop_3_29_pdst},
     {rob_uop_3_28_pdst},
     {rob_uop_3_27_pdst},
     {rob_uop_3_26_pdst},
     {rob_uop_3_25_pdst},
     {rob_uop_3_24_pdst},
     {rob_uop_3_23_pdst},
     {rob_uop_3_22_pdst},
     {rob_uop_3_21_pdst},
     {rob_uop_3_20_pdst},
     {rob_uop_3_19_pdst},
     {rob_uop_3_18_pdst},
     {rob_uop_3_17_pdst},
     {rob_uop_3_16_pdst},
     {rob_uop_3_15_pdst},
     {rob_uop_3_14_pdst},
     {rob_uop_3_13_pdst},
     {rob_uop_3_12_pdst},
     {rob_uop_3_11_pdst},
     {rob_uop_3_10_pdst},
     {rob_uop_3_9_pdst},
     {rob_uop_3_8_pdst},
     {rob_uop_3_7_pdst},
     {rob_uop_3_6_pdst},
     {rob_uop_3_5_pdst},
     {rob_uop_3_4_pdst},
     {rob_uop_3_3_pdst},
     {rob_uop_3_2_pdst},
     {rob_uop_3_1_pdst},
     {rob_uop_3_0_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_129 =
    {{rob_uop_3_31_stale_pdst},
     {rob_uop_3_30_stale_pdst},
     {rob_uop_3_29_stale_pdst},
     {rob_uop_3_28_stale_pdst},
     {rob_uop_3_27_stale_pdst},
     {rob_uop_3_26_stale_pdst},
     {rob_uop_3_25_stale_pdst},
     {rob_uop_3_24_stale_pdst},
     {rob_uop_3_23_stale_pdst},
     {rob_uop_3_22_stale_pdst},
     {rob_uop_3_21_stale_pdst},
     {rob_uop_3_20_stale_pdst},
     {rob_uop_3_19_stale_pdst},
     {rob_uop_3_18_stale_pdst},
     {rob_uop_3_17_stale_pdst},
     {rob_uop_3_16_stale_pdst},
     {rob_uop_3_15_stale_pdst},
     {rob_uop_3_14_stale_pdst},
     {rob_uop_3_13_stale_pdst},
     {rob_uop_3_12_stale_pdst},
     {rob_uop_3_11_stale_pdst},
     {rob_uop_3_10_stale_pdst},
     {rob_uop_3_9_stale_pdst},
     {rob_uop_3_8_stale_pdst},
     {rob_uop_3_7_stale_pdst},
     {rob_uop_3_6_stale_pdst},
     {rob_uop_3_5_stale_pdst},
     {rob_uop_3_4_stale_pdst},
     {rob_uop_3_3_stale_pdst},
     {rob_uop_3_2_stale_pdst},
     {rob_uop_3_1_stale_pdst},
     {rob_uop_3_0_stale_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_130 =
    {{rob_uop_3_31_is_fencei},
     {rob_uop_3_30_is_fencei},
     {rob_uop_3_29_is_fencei},
     {rob_uop_3_28_is_fencei},
     {rob_uop_3_27_is_fencei},
     {rob_uop_3_26_is_fencei},
     {rob_uop_3_25_is_fencei},
     {rob_uop_3_24_is_fencei},
     {rob_uop_3_23_is_fencei},
     {rob_uop_3_22_is_fencei},
     {rob_uop_3_21_is_fencei},
     {rob_uop_3_20_is_fencei},
     {rob_uop_3_19_is_fencei},
     {rob_uop_3_18_is_fencei},
     {rob_uop_3_17_is_fencei},
     {rob_uop_3_16_is_fencei},
     {rob_uop_3_15_is_fencei},
     {rob_uop_3_14_is_fencei},
     {rob_uop_3_13_is_fencei},
     {rob_uop_3_12_is_fencei},
     {rob_uop_3_11_is_fencei},
     {rob_uop_3_10_is_fencei},
     {rob_uop_3_9_is_fencei},
     {rob_uop_3_8_is_fencei},
     {rob_uop_3_7_is_fencei},
     {rob_uop_3_6_is_fencei},
     {rob_uop_3_5_is_fencei},
     {rob_uop_3_4_is_fencei},
     {rob_uop_3_3_is_fencei},
     {rob_uop_3_2_is_fencei},
     {rob_uop_3_1_is_fencei},
     {rob_uop_3_0_is_fencei}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_131 =
    {{rob_uop_3_31_uses_ldq},
     {rob_uop_3_30_uses_ldq},
     {rob_uop_3_29_uses_ldq},
     {rob_uop_3_28_uses_ldq},
     {rob_uop_3_27_uses_ldq},
     {rob_uop_3_26_uses_ldq},
     {rob_uop_3_25_uses_ldq},
     {rob_uop_3_24_uses_ldq},
     {rob_uop_3_23_uses_ldq},
     {rob_uop_3_22_uses_ldq},
     {rob_uop_3_21_uses_ldq},
     {rob_uop_3_20_uses_ldq},
     {rob_uop_3_19_uses_ldq},
     {rob_uop_3_18_uses_ldq},
     {rob_uop_3_17_uses_ldq},
     {rob_uop_3_16_uses_ldq},
     {rob_uop_3_15_uses_ldq},
     {rob_uop_3_14_uses_ldq},
     {rob_uop_3_13_uses_ldq},
     {rob_uop_3_12_uses_ldq},
     {rob_uop_3_11_uses_ldq},
     {rob_uop_3_10_uses_ldq},
     {rob_uop_3_9_uses_ldq},
     {rob_uop_3_8_uses_ldq},
     {rob_uop_3_7_uses_ldq},
     {rob_uop_3_6_uses_ldq},
     {rob_uop_3_5_uses_ldq},
     {rob_uop_3_4_uses_ldq},
     {rob_uop_3_3_uses_ldq},
     {rob_uop_3_2_uses_ldq},
     {rob_uop_3_1_uses_ldq},
     {rob_uop_3_0_uses_ldq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_132 =
    {{rob_uop_3_31_uses_stq},
     {rob_uop_3_30_uses_stq},
     {rob_uop_3_29_uses_stq},
     {rob_uop_3_28_uses_stq},
     {rob_uop_3_27_uses_stq},
     {rob_uop_3_26_uses_stq},
     {rob_uop_3_25_uses_stq},
     {rob_uop_3_24_uses_stq},
     {rob_uop_3_23_uses_stq},
     {rob_uop_3_22_uses_stq},
     {rob_uop_3_21_uses_stq},
     {rob_uop_3_20_uses_stq},
     {rob_uop_3_19_uses_stq},
     {rob_uop_3_18_uses_stq},
     {rob_uop_3_17_uses_stq},
     {rob_uop_3_16_uses_stq},
     {rob_uop_3_15_uses_stq},
     {rob_uop_3_14_uses_stq},
     {rob_uop_3_13_uses_stq},
     {rob_uop_3_12_uses_stq},
     {rob_uop_3_11_uses_stq},
     {rob_uop_3_10_uses_stq},
     {rob_uop_3_9_uses_stq},
     {rob_uop_3_8_uses_stq},
     {rob_uop_3_7_uses_stq},
     {rob_uop_3_6_uses_stq},
     {rob_uop_3_5_uses_stq},
     {rob_uop_3_4_uses_stq},
     {rob_uop_3_3_uses_stq},
     {rob_uop_3_2_uses_stq},
     {rob_uop_3_1_uses_stq},
     {rob_uop_3_0_uses_stq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_133 =
    {{rob_uop_3_31_is_sys_pc2epc},
     {rob_uop_3_30_is_sys_pc2epc},
     {rob_uop_3_29_is_sys_pc2epc},
     {rob_uop_3_28_is_sys_pc2epc},
     {rob_uop_3_27_is_sys_pc2epc},
     {rob_uop_3_26_is_sys_pc2epc},
     {rob_uop_3_25_is_sys_pc2epc},
     {rob_uop_3_24_is_sys_pc2epc},
     {rob_uop_3_23_is_sys_pc2epc},
     {rob_uop_3_22_is_sys_pc2epc},
     {rob_uop_3_21_is_sys_pc2epc},
     {rob_uop_3_20_is_sys_pc2epc},
     {rob_uop_3_19_is_sys_pc2epc},
     {rob_uop_3_18_is_sys_pc2epc},
     {rob_uop_3_17_is_sys_pc2epc},
     {rob_uop_3_16_is_sys_pc2epc},
     {rob_uop_3_15_is_sys_pc2epc},
     {rob_uop_3_14_is_sys_pc2epc},
     {rob_uop_3_13_is_sys_pc2epc},
     {rob_uop_3_12_is_sys_pc2epc},
     {rob_uop_3_11_is_sys_pc2epc},
     {rob_uop_3_10_is_sys_pc2epc},
     {rob_uop_3_9_is_sys_pc2epc},
     {rob_uop_3_8_is_sys_pc2epc},
     {rob_uop_3_7_is_sys_pc2epc},
     {rob_uop_3_6_is_sys_pc2epc},
     {rob_uop_3_5_is_sys_pc2epc},
     {rob_uop_3_4_is_sys_pc2epc},
     {rob_uop_3_3_is_sys_pc2epc},
     {rob_uop_3_2_is_sys_pc2epc},
     {rob_uop_3_1_is_sys_pc2epc},
     {rob_uop_3_0_is_sys_pc2epc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_134 =
    {{rob_uop_3_31_flush_on_commit},
     {rob_uop_3_30_flush_on_commit},
     {rob_uop_3_29_flush_on_commit},
     {rob_uop_3_28_flush_on_commit},
     {rob_uop_3_27_flush_on_commit},
     {rob_uop_3_26_flush_on_commit},
     {rob_uop_3_25_flush_on_commit},
     {rob_uop_3_24_flush_on_commit},
     {rob_uop_3_23_flush_on_commit},
     {rob_uop_3_22_flush_on_commit},
     {rob_uop_3_21_flush_on_commit},
     {rob_uop_3_20_flush_on_commit},
     {rob_uop_3_19_flush_on_commit},
     {rob_uop_3_18_flush_on_commit},
     {rob_uop_3_17_flush_on_commit},
     {rob_uop_3_16_flush_on_commit},
     {rob_uop_3_15_flush_on_commit},
     {rob_uop_3_14_flush_on_commit},
     {rob_uop_3_13_flush_on_commit},
     {rob_uop_3_12_flush_on_commit},
     {rob_uop_3_11_flush_on_commit},
     {rob_uop_3_10_flush_on_commit},
     {rob_uop_3_9_flush_on_commit},
     {rob_uop_3_8_flush_on_commit},
     {rob_uop_3_7_flush_on_commit},
     {rob_uop_3_6_flush_on_commit},
     {rob_uop_3_5_flush_on_commit},
     {rob_uop_3_4_flush_on_commit},
     {rob_uop_3_3_flush_on_commit},
     {rob_uop_3_2_flush_on_commit},
     {rob_uop_3_1_flush_on_commit},
     {rob_uop_3_0_flush_on_commit}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_135 =
    {{rob_uop_3_31_ldst},
     {rob_uop_3_30_ldst},
     {rob_uop_3_29_ldst},
     {rob_uop_3_28_ldst},
     {rob_uop_3_27_ldst},
     {rob_uop_3_26_ldst},
     {rob_uop_3_25_ldst},
     {rob_uop_3_24_ldst},
     {rob_uop_3_23_ldst},
     {rob_uop_3_22_ldst},
     {rob_uop_3_21_ldst},
     {rob_uop_3_20_ldst},
     {rob_uop_3_19_ldst},
     {rob_uop_3_18_ldst},
     {rob_uop_3_17_ldst},
     {rob_uop_3_16_ldst},
     {rob_uop_3_15_ldst},
     {rob_uop_3_14_ldst},
     {rob_uop_3_13_ldst},
     {rob_uop_3_12_ldst},
     {rob_uop_3_11_ldst},
     {rob_uop_3_10_ldst},
     {rob_uop_3_9_ldst},
     {rob_uop_3_8_ldst},
     {rob_uop_3_7_ldst},
     {rob_uop_3_6_ldst},
     {rob_uop_3_5_ldst},
     {rob_uop_3_4_ldst},
     {rob_uop_3_3_ldst},
     {rob_uop_3_2_ldst},
     {rob_uop_3_1_ldst},
     {rob_uop_3_0_ldst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_136 =
    {{rob_uop_3_31_ldst_val},
     {rob_uop_3_30_ldst_val},
     {rob_uop_3_29_ldst_val},
     {rob_uop_3_28_ldst_val},
     {rob_uop_3_27_ldst_val},
     {rob_uop_3_26_ldst_val},
     {rob_uop_3_25_ldst_val},
     {rob_uop_3_24_ldst_val},
     {rob_uop_3_23_ldst_val},
     {rob_uop_3_22_ldst_val},
     {rob_uop_3_21_ldst_val},
     {rob_uop_3_20_ldst_val},
     {rob_uop_3_19_ldst_val},
     {rob_uop_3_18_ldst_val},
     {rob_uop_3_17_ldst_val},
     {rob_uop_3_16_ldst_val},
     {rob_uop_3_15_ldst_val},
     {rob_uop_3_14_ldst_val},
     {rob_uop_3_13_ldst_val},
     {rob_uop_3_12_ldst_val},
     {rob_uop_3_11_ldst_val},
     {rob_uop_3_10_ldst_val},
     {rob_uop_3_9_ldst_val},
     {rob_uop_3_8_ldst_val},
     {rob_uop_3_7_ldst_val},
     {rob_uop_3_6_ldst_val},
     {rob_uop_3_5_ldst_val},
     {rob_uop_3_4_ldst_val},
     {rob_uop_3_3_ldst_val},
     {rob_uop_3_2_ldst_val},
     {rob_uop_3_1_ldst_val},
     {rob_uop_3_0_ldst_val}};	// rob.scala:310:28, :411:25
  wire [31:0][1:0] _GEN_137 =
    {{rob_uop_3_31_dst_rtype},
     {rob_uop_3_30_dst_rtype},
     {rob_uop_3_29_dst_rtype},
     {rob_uop_3_28_dst_rtype},
     {rob_uop_3_27_dst_rtype},
     {rob_uop_3_26_dst_rtype},
     {rob_uop_3_25_dst_rtype},
     {rob_uop_3_24_dst_rtype},
     {rob_uop_3_23_dst_rtype},
     {rob_uop_3_22_dst_rtype},
     {rob_uop_3_21_dst_rtype},
     {rob_uop_3_20_dst_rtype},
     {rob_uop_3_19_dst_rtype},
     {rob_uop_3_18_dst_rtype},
     {rob_uop_3_17_dst_rtype},
     {rob_uop_3_16_dst_rtype},
     {rob_uop_3_15_dst_rtype},
     {rob_uop_3_14_dst_rtype},
     {rob_uop_3_13_dst_rtype},
     {rob_uop_3_12_dst_rtype},
     {rob_uop_3_11_dst_rtype},
     {rob_uop_3_10_dst_rtype},
     {rob_uop_3_9_dst_rtype},
     {rob_uop_3_8_dst_rtype},
     {rob_uop_3_7_dst_rtype},
     {rob_uop_3_6_dst_rtype},
     {rob_uop_3_5_dst_rtype},
     {rob_uop_3_4_dst_rtype},
     {rob_uop_3_3_dst_rtype},
     {rob_uop_3_2_dst_rtype},
     {rob_uop_3_1_dst_rtype},
     {rob_uop_3_0_dst_rtype}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_138 =
    {{rob_uop_3_31_fp_val},
     {rob_uop_3_30_fp_val},
     {rob_uop_3_29_fp_val},
     {rob_uop_3_28_fp_val},
     {rob_uop_3_27_fp_val},
     {rob_uop_3_26_fp_val},
     {rob_uop_3_25_fp_val},
     {rob_uop_3_24_fp_val},
     {rob_uop_3_23_fp_val},
     {rob_uop_3_22_fp_val},
     {rob_uop_3_21_fp_val},
     {rob_uop_3_20_fp_val},
     {rob_uop_3_19_fp_val},
     {rob_uop_3_18_fp_val},
     {rob_uop_3_17_fp_val},
     {rob_uop_3_16_fp_val},
     {rob_uop_3_15_fp_val},
     {rob_uop_3_14_fp_val},
     {rob_uop_3_13_fp_val},
     {rob_uop_3_12_fp_val},
     {rob_uop_3_11_fp_val},
     {rob_uop_3_10_fp_val},
     {rob_uop_3_9_fp_val},
     {rob_uop_3_8_fp_val},
     {rob_uop_3_7_fp_val},
     {rob_uop_3_6_fp_val},
     {rob_uop_3_5_fp_val},
     {rob_uop_3_4_fp_val},
     {rob_uop_3_3_fp_val},
     {rob_uop_3_2_fp_val},
     {rob_uop_3_1_fp_val},
     {rob_uop_3_0_fp_val}};	// rob.scala:310:28, :411:25
  wire             rbk_row_3 = _io_commit_rollback_T_3 & ~full;	// rob.scala:236:31, :425:{44,47}, :787:39
  wire             _io_commit_rbk_valids_3_output = rbk_row_3 & _GEN_104[com_idx];	// rob.scala:236:20, :324:31, :425:44, :427:40
  reg              block_commit_REG;	// rob.scala:540:94
  reg              block_commit_REG_1;	// rob.scala:540:131
  reg              block_commit_REG_2;	// rob.scala:540:123
  wire             block_commit =
    rob_state != 2'h1 & rob_state != 2'h3 | block_commit_REG | block_commit_REG_2;	// rob.scala:221:26, :419:36, :540:{33,47,61,94,113,123}
  assign will_commit_0 = can_commit_0 & ~can_throw_exception_0 & ~block_commit;	// rob.scala:398:49, :404:64, :540:113, :545:55, :547:{46,70}
  wire             _GEN_139 =
    rob_head_vals_0 & (~can_commit_0 | can_throw_exception_0) | block_commit;	// rob.scala:398:49, :404:64, :540:113, :548:46, :549:{29,44,72}
  assign will_commit_1 = can_commit_1 & ~can_throw_exception_1 & ~_GEN_139;	// rob.scala:398:49, :404:64, :545:55, :547:{46,70}, :549:72
  wire             _GEN_140 =
    rob_head_vals_1 & (~can_commit_1 | can_throw_exception_1) | _GEN_139;	// rob.scala:398:49, :404:64, :548:46, :549:{29,44,72}
  assign will_commit_2 = can_commit_2 & ~can_throw_exception_2 & ~_GEN_140;	// rob.scala:398:49, :404:64, :545:55, :547:{46,70}, :549:72
  wire             _GEN_141 =
    rob_head_vals_2 & (~can_commit_2 | can_throw_exception_2) | _GEN_140;	// rob.scala:398:49, :404:64, :548:46, :549:{29,44,72}
  wire             exception_thrown =
    can_throw_exception_3 & ~_GEN_141 & ~will_commit_2 | can_throw_exception_2 & ~_GEN_140
    & ~will_commit_1 | can_throw_exception_1 & ~_GEN_139 & ~will_commit_0
    | can_throw_exception_0 & ~block_commit;	// rob.scala:398:49, :540:113, :545:{52,55,69,72,85}, :547:70, :549:72
  assign will_commit_3 =
    rob_head_vals_3 & ~_GEN_116[rob_head] & ~io_csr_stall & ~can_throw_exception_3
    & ~_GEN_141;	// rob.scala:224:29, :366:31, :398:49, :404:{43,67}, :545:55, :547:{46,70}, :549:72
  wire             _io_flush_bits_flush_typ_T = r_xcpt_uop_exc_cause != 64'h10;	// rob.scala:259:29, :556:50
  wire [5:0]       com_xcpt_uop_ftq_idx =
    rob_head_vals_0
      ? _GEN_20[com_idx]
      : rob_head_vals_1
          ? _GEN_55[com_idx]
          : rob_head_vals_2 ? _GEN_90[com_idx] : _GEN_125[com_idx];	// Mux.scala:47:69, rob.scala:236:20, :398:49, :411:25
  wire             com_xcpt_uop_edge_inst =
    rob_head_vals_0
      ? _GEN_21[com_idx]
      : rob_head_vals_1
          ? _GEN_56[com_idx]
          : rob_head_vals_2 ? _GEN_91[com_idx] : _GEN_126[com_idx];	// Mux.scala:47:69, rob.scala:236:20, :398:49, :411:25
  wire [5:0]       com_xcpt_uop_pc_lob =
    rob_head_vals_0
      ? _GEN_22[com_idx]
      : rob_head_vals_1
          ? _GEN_57[com_idx]
          : rob_head_vals_2 ? _GEN_92[com_idx] : _GEN_127[com_idx];	// Mux.scala:47:69, rob.scala:236:20, :398:49, :411:25
  wire             flush_commit_mask_0 = will_commit_0 & _GEN_29[com_idx];	// rob.scala:236:20, :411:25, :547:70, :571:75
  wire             flush_commit_mask_1 = will_commit_1 & _GEN_64[com_idx];	// rob.scala:236:20, :411:25, :547:70, :571:75
  wire             flush_commit_mask_2 = will_commit_2 & _GEN_99[com_idx];	// rob.scala:236:20, :411:25, :547:70, :571:75
  wire             flush_commit_mask_3 = will_commit_3 & _GEN_134[com_idx];	// rob.scala:236:20, :411:25, :547:70, :571:75
  wire             flush_commit =
    flush_commit_mask_0 | flush_commit_mask_1 | flush_commit_mask_2 | flush_commit_mask_3;	// rob.scala:571:75, :572:48
  wire             _io_flush_valid_output = exception_thrown | flush_commit;	// rob.scala:545:85, :572:48, :573:36
  wire             _fflags_val_0_T = will_commit_0 & _GEN_33[com_idx];	// rob.scala:236:20, :411:25, :547:70, :601:27
  wire             fflags_val_0 = _fflags_val_0_T & ~_GEN_27[com_idx];	// rob.scala:236:20, :411:25, :601:27, :602:32, :603:7
  wire             _fflags_val_1_T = will_commit_1 & _GEN_68[com_idx];	// rob.scala:236:20, :411:25, :547:70, :601:27
  wire             fflags_val_1 = _fflags_val_1_T & ~_GEN_62[com_idx];	// rob.scala:236:20, :411:25, :601:27, :602:32, :603:7
  wire             _fflags_val_2_T = will_commit_2 & _GEN_103[com_idx];	// rob.scala:236:20, :411:25, :547:70, :601:27
  wire             fflags_val_2 = _fflags_val_2_T & ~_GEN_97[com_idx];	// rob.scala:236:20, :411:25, :601:27, :602:32, :603:7
  wire             _fflags_val_3_T = will_commit_3 & _GEN_138[com_idx];	// rob.scala:236:20, :411:25, :547:70, :601:27
  wire             fflags_val_3 = _fflags_val_3_T & ~_GEN_132[com_idx];	// rob.scala:236:20, :411:25, :601:27, :602:32, :603:7
  reg              r_partial_row;	// rob.scala:677:30
  wire             _empty_T = rob_head == rob_tail;	// rob.scala:224:29, :228:29, :686:33
  wire             finished_committing_row =
    (|{will_commit_3, will_commit_2, will_commit_1, will_commit_0})
    & ({will_commit_3, will_commit_2, will_commit_1, will_commit_0}
       ^ {rob_head_vals_3, rob_head_vals_2, rob_head_vals_1, rob_head_vals_0}) == 4'h0
    & ~(r_partial_row & _empty_T & ~maybe_full);	// rob.scala:239:29, :287:15, :398:49, :547:70, :677:30, :684:{23,30}, :685:{19,26,42,50,59}, :686:{5,33,46,49}
  reg              pnr_maybe_at_tail;	// rob.scala:714:36
  wire             _io_ready_T = rob_state == 2'h1;	// rob.scala:221:26, :540:33, :716:33
  `ifndef SYNTHESIS	// rob.scala:333:14
    always @(posedge clock) begin	// rob.scala:333:14
      automatic logic [6:0] rob_pnr_idx;	// Cat.scala:30:58
      automatic logic       _GEN_142 = io_lxcpt_bits_cause != 5'h10;	// rob.scala:324:31, :392:33
      automatic logic       _GEN_143 =
        ~((will_commit_0 | will_commit_1 | will_commit_2 | will_commit_3)
          & (_io_commit_rbk_valids_0_output | _io_commit_rbk_valids_1_output
             | _io_commit_rbk_valids_2_output | _io_commit_rbk_valids_3_output)) | reset;	// rob.scala:427:40, :430:{12,13,40,45,77}, :547:70
      automatic logic       _GEN_144;	// util.scala:363:52
      automatic logic [2:0] _GEN_145 =
        {1'h0, {1'h0, flush_commit_mask_0} + {1'h0, flush_commit_mask_1}}
        + {1'h0, {1'h0, flush_commit_mask_2} + {1'h0, flush_commit_mask_3}};	// Bitwise.scala:47:55, rob.scala:370:{23,59}, :372:26, :381:32, :571:75
      rob_pnr_idx = {rob_pnr, rob_pnr_lsb};	// Cat.scala:30:58, rob.scala:232:29, :233:29
      _GEN_144 = rob_pnr_idx < rob_head_idx;	// Cat.scala:30:58, util.scala:363:52
      if (io_enq_valids_0 & ~(~rob_tail_vals_0 | reset)) begin	// rob.scala:324:31, :333:{14,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:333:14
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");	// rob.scala:333:14
        if (`STOP_COND_)	// rob.scala:333:14
          $fatal;	// rob.scala:333:14
      end
      if (io_enq_valids_0 & ~(io_enq_uops_0_rob_idx[6:2] == rob_tail | reset)) begin	// rob.scala:228:29, :334:{14,39,63}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:334:14
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");	// rob.scala:334:14
        if (`STOP_COND_)	// rob.scala:334:14
          $fatal;	// rob.scala:334:14
      end
      if (_GEN_10 & ~(_GEN[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_10 & ~(_GEN_11[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_12 & ~(_GEN[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_12 & ~(_GEN_11[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_13 & ~(_GEN[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_13 & ~(_GEN_11[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_14 & _GEN_142 & ~(_GEN_15[io_lxcpt_bits_uop_rob_idx[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :390:26, :392:33, :394:15
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:394:15
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");	// rob.scala:394:15
        if (`STOP_COND_)	// rob.scala:394:15
          $fatal;	// rob.scala:394:15
      end
      if (~_GEN_143) begin	// rob.scala:430:12
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:430:12
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");	// rob.scala:430:12
        if (`STOP_COND_)	// rob.scala:430:12
          $fatal;	// rob.scala:430:12
      end
      if (~(~(_GEN_0 & ~_GEN[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_0 & ~_GEN_11[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_0 & _GEN_31[io_wb_resps_0_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_0_bits_uop_rob_idx[6:2]] != io_wb_resps_0_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_1 & ~_GEN[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_1 & ~_GEN_11[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_1 & _GEN_31[io_wb_resps_1_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_1_bits_uop_rob_idx[6:2]] != io_wb_resps_1_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_2 & ~_GEN[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_2 & ~_GEN_11[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_2 & _GEN_31[io_wb_resps_2_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_2_bits_uop_rob_idx[6:2]] != io_wb_resps_2_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_3 & ~_GEN[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_3 & ~_GEN_11[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_3 & _GEN_31[io_wb_resps_3_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_3_bits_uop_rob_idx[6:2]] != io_wb_resps_3_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_4 & ~_GEN[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_4 & ~_GEN_11[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_4 & _GEN_31[io_wb_resps_4_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_4_bits_uop_rob_idx[6:2]] != io_wb_resps_4_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_5 & ~_GEN[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_5 & ~_GEN_11[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_5 & _GEN_31[io_wb_resps_5_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_5_bits_uop_rob_idx[6:2]] != io_wb_resps_5_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_6 & ~_GEN[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_6 & ~_GEN_11[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_6 & _GEN_31[io_wb_resps_6_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_6_bits_uop_rob_idx[6:2]] != io_wb_resps_6_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_7 & ~_GEN[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_7 & ~_GEN_11[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_7 & _GEN_31[io_wb_resps_7_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_7_bits_uop_rob_idx[6:2]] != io_wb_resps_7_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_8 & ~_GEN[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_8 & ~_GEN_11[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_8 & _GEN_31[io_wb_resps_8_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_8_bits_uop_rob_idx[6:2]] != io_wb_resps_8_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_9 & ~_GEN[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_9 & ~_GEN_11[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_9 & _GEN_31[io_wb_resps_9_bits_uop_rob_idx[6:2]]
              & _GEN_23[io_wb_resps_9_bits_uop_rob_idx[6:2]] != io_wb_resps_9_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (io_enq_valids_1 & ~(~rob_tail_vals_1 | reset)) begin	// rob.scala:324:31, :333:{14,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:333:14
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");	// rob.scala:333:14
        if (`STOP_COND_)	// rob.scala:333:14
          $fatal;	// rob.scala:333:14
      end
      if (io_enq_valids_1 & ~(io_enq_uops_1_rob_idx[6:2] == rob_tail | reset)) begin	// rob.scala:228:29, :334:{14,39,63}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:334:14
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");	// rob.scala:334:14
        if (`STOP_COND_)	// rob.scala:334:14
          $fatal;	// rob.scala:334:14
      end
      if (_GEN_45 & ~(_GEN_34[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_45 & ~(_GEN_46[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_47 & ~(_GEN_34[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_47 & ~(_GEN_46[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_48 & ~(_GEN_34[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_48 & ~(_GEN_46[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_49 & _GEN_142 & ~(_GEN_50[io_lxcpt_bits_uop_rob_idx[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :390:26, :392:33, :394:15
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:394:15
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");	// rob.scala:394:15
        if (`STOP_COND_)	// rob.scala:394:15
          $fatal;	// rob.scala:394:15
      end
      if (~_GEN_143) begin	// rob.scala:430:12
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:430:12
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");	// rob.scala:430:12
        if (`STOP_COND_)	// rob.scala:430:12
          $fatal;	// rob.scala:430:12
      end
      if (~(~(_GEN_35 & ~_GEN_34[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_35 & ~_GEN_46[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_35 & _GEN_66[io_wb_resps_0_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_0_bits_uop_rob_idx[6:2]] != io_wb_resps_0_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_36 & ~_GEN_34[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_36 & ~_GEN_46[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_36 & _GEN_66[io_wb_resps_1_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_1_bits_uop_rob_idx[6:2]] != io_wb_resps_1_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_37 & ~_GEN_34[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_37 & ~_GEN_46[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_37 & _GEN_66[io_wb_resps_2_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_2_bits_uop_rob_idx[6:2]] != io_wb_resps_2_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_38 & ~_GEN_34[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_38 & ~_GEN_46[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_38 & _GEN_66[io_wb_resps_3_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_3_bits_uop_rob_idx[6:2]] != io_wb_resps_3_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_39 & ~_GEN_34[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_39 & ~_GEN_46[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_39 & _GEN_66[io_wb_resps_4_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_4_bits_uop_rob_idx[6:2]] != io_wb_resps_4_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_40 & ~_GEN_34[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_40 & ~_GEN_46[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_40 & _GEN_66[io_wb_resps_5_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_5_bits_uop_rob_idx[6:2]] != io_wb_resps_5_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_41 & ~_GEN_34[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_41 & ~_GEN_46[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_41 & _GEN_66[io_wb_resps_6_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_6_bits_uop_rob_idx[6:2]] != io_wb_resps_6_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_42 & ~_GEN_34[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_42 & ~_GEN_46[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_42 & _GEN_66[io_wb_resps_7_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_7_bits_uop_rob_idx[6:2]] != io_wb_resps_7_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_43 & ~_GEN_34[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_43 & ~_GEN_46[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_43 & _GEN_66[io_wb_resps_8_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_8_bits_uop_rob_idx[6:2]] != io_wb_resps_8_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_44 & ~_GEN_34[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_44 & ~_GEN_46[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_44 & _GEN_66[io_wb_resps_9_bits_uop_rob_idx[6:2]]
              & _GEN_58[io_wb_resps_9_bits_uop_rob_idx[6:2]] != io_wb_resps_9_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (io_enq_valids_2 & ~(~rob_tail_vals_2 | reset)) begin	// rob.scala:324:31, :333:{14,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:333:14
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");	// rob.scala:333:14
        if (`STOP_COND_)	// rob.scala:333:14
          $fatal;	// rob.scala:333:14
      end
      if (io_enq_valids_2 & ~(io_enq_uops_2_rob_idx[6:2] == rob_tail | reset)) begin	// rob.scala:228:29, :334:{14,39,63}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:334:14
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");	// rob.scala:334:14
        if (`STOP_COND_)	// rob.scala:334:14
          $fatal;	// rob.scala:334:14
      end
      if (_GEN_80 & ~(_GEN_69[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_80 & ~(_GEN_81[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_82 & ~(_GEN_69[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_82 & ~(_GEN_81[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_83 & ~(_GEN_69[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_83 & ~(_GEN_81[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_84 & _GEN_142 & ~(_GEN_85[io_lxcpt_bits_uop_rob_idx[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :390:26, :392:33, :394:15
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:394:15
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");	// rob.scala:394:15
        if (`STOP_COND_)	// rob.scala:394:15
          $fatal;	// rob.scala:394:15
      end
      if (~_GEN_143) begin	// rob.scala:430:12
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:430:12
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");	// rob.scala:430:12
        if (`STOP_COND_)	// rob.scala:430:12
          $fatal;	// rob.scala:430:12
      end
      if (~(~(_GEN_70 & ~_GEN_69[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_70 & ~_GEN_81[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_70 & _GEN_101[io_wb_resps_0_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_0_bits_uop_rob_idx[6:2]] != io_wb_resps_0_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_71 & ~_GEN_69[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_71 & ~_GEN_81[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_71 & _GEN_101[io_wb_resps_1_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_1_bits_uop_rob_idx[6:2]] != io_wb_resps_1_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_72 & ~_GEN_69[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_72 & ~_GEN_81[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_72 & _GEN_101[io_wb_resps_2_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_2_bits_uop_rob_idx[6:2]] != io_wb_resps_2_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_73 & ~_GEN_69[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_73 & ~_GEN_81[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_73 & _GEN_101[io_wb_resps_3_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_3_bits_uop_rob_idx[6:2]] != io_wb_resps_3_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_74 & ~_GEN_69[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_74 & ~_GEN_81[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_74 & _GEN_101[io_wb_resps_4_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_4_bits_uop_rob_idx[6:2]] != io_wb_resps_4_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_75 & ~_GEN_69[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_75 & ~_GEN_81[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_75 & _GEN_101[io_wb_resps_5_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_5_bits_uop_rob_idx[6:2]] != io_wb_resps_5_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_76 & ~_GEN_69[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_76 & ~_GEN_81[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_76 & _GEN_101[io_wb_resps_6_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_6_bits_uop_rob_idx[6:2]] != io_wb_resps_6_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_77 & ~_GEN_69[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_77 & ~_GEN_81[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_77 & _GEN_101[io_wb_resps_7_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_7_bits_uop_rob_idx[6:2]] != io_wb_resps_7_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_78 & ~_GEN_69[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_78 & ~_GEN_81[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_78 & _GEN_101[io_wb_resps_8_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_8_bits_uop_rob_idx[6:2]] != io_wb_resps_8_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_79 & ~_GEN_69[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_79 & ~_GEN_81[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_79 & _GEN_101[io_wb_resps_9_bits_uop_rob_idx[6:2]]
              & _GEN_93[io_wb_resps_9_bits_uop_rob_idx[6:2]] != io_wb_resps_9_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (io_enq_valids_3 & ~(~rob_tail_vals_3 | reset)) begin	// rob.scala:324:31, :333:{14,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:333:14
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");	// rob.scala:333:14
        if (`STOP_COND_)	// rob.scala:333:14
          $fatal;	// rob.scala:333:14
      end
      if (io_enq_valids_3 & ~(io_enq_uops_3_rob_idx[6:2] == rob_tail | reset)) begin	// rob.scala:228:29, :334:{14,39,63}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:334:14
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");	// rob.scala:334:14
        if (`STOP_COND_)	// rob.scala:334:14
          $fatal;	// rob.scala:334:14
      end
      if (_GEN_115 & ~(_GEN_104[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_115 & ~(_GEN_116[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_117 & ~(_GEN_104[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_117 & ~(_GEN_116[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_118 & ~(_GEN_104[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_118 & ~(_GEN_116[io_lsu_clr_bsy_2_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_119 & _GEN_142 & ~(_GEN_120[io_lxcpt_bits_uop_rob_idx[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :390:26, :392:33, :394:15
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:394:15
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");	// rob.scala:394:15
        if (`STOP_COND_)	// rob.scala:394:15
          $fatal;	// rob.scala:394:15
      end
      if (~_GEN_143) begin	// rob.scala:430:12
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:430:12
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");	// rob.scala:430:12
        if (`STOP_COND_)	// rob.scala:430:12
          $fatal;	// rob.scala:430:12
      end
      if (~(~(_GEN_105 & ~_GEN_104[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_105 & ~_GEN_116[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_105 & _GEN_136[io_wb_resps_0_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_0_bits_uop_rob_idx[6:2]] != io_wb_resps_0_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_106 & ~_GEN_104[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_106 & ~_GEN_116[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_106 & _GEN_136[io_wb_resps_1_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_1_bits_uop_rob_idx[6:2]] != io_wb_resps_1_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_107 & ~_GEN_104[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_107 & ~_GEN_116[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_107 & _GEN_136[io_wb_resps_2_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_2_bits_uop_rob_idx[6:2]] != io_wb_resps_2_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_108 & ~_GEN_104[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_108 & ~_GEN_116[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_108 & _GEN_136[io_wb_resps_3_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_3_bits_uop_rob_idx[6:2]] != io_wb_resps_3_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_109 & ~_GEN_104[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_109 & ~_GEN_116[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_109 & _GEN_136[io_wb_resps_4_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_4_bits_uop_rob_idx[6:2]] != io_wb_resps_4_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_110 & ~_GEN_104[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_110 & ~_GEN_116[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_110 & _GEN_136[io_wb_resps_5_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_5_bits_uop_rob_idx[6:2]] != io_wb_resps_5_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_111 & ~_GEN_104[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_111 & ~_GEN_116[io_wb_resps_6_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_111 & _GEN_136[io_wb_resps_6_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_6_bits_uop_rob_idx[6:2]] != io_wb_resps_6_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_112 & ~_GEN_104[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_112 & ~_GEN_116[io_wb_resps_7_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_112 & _GEN_136[io_wb_resps_7_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_7_bits_uop_rob_idx[6:2]] != io_wb_resps_7_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_113 & ~_GEN_104[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_113 & ~_GEN_116[io_wb_resps_8_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_113 & _GEN_136[io_wb_resps_8_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_8_bits_uop_rob_idx[6:2]] != io_wb_resps_8_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_114 & ~_GEN_104[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_114 & ~_GEN_116[io_wb_resps_9_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_114 & _GEN_136[io_wb_resps_9_bits_uop_rob_idx[6:2]]
              & _GEN_128[io_wb_resps_9_bits_uop_rob_idx[6:2]] != io_wb_resps_9_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(_GEN_145[2:1] == 2'h0 | reset)) begin	// Bitwise.scala:47:55, rob.scala:221:26, :575:{9,40}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:575:9
          $error("Assertion failed: [rob] Can't commit multiple flush_on_commit instructions on one cycle\n    at rob.scala:575 assert(!(PopCount(flush_commit_mask) > 1.U),\n");	// rob.scala:575:9
        if (`STOP_COND_)	// rob.scala:575:9
          $fatal;	// rob.scala:575:9
      end
      if (~(~(will_commit_0 & ~_GEN_33[com_idx] & (|_rob_fflags_ext_R0_data))
            | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :547:70, :607:{12,13}, :608:{14,40}, :609:33
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:607:12
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n");	// rob.scala:607:12
        if (`STOP_COND_)	// rob.scala:607:12
          $fatal;	// rob.scala:607:12
      end
      if (~(~(_fflags_val_0_T & (_GEN_26[com_idx] | _GEN_27[com_idx])
              & (|_rob_fflags_ext_R0_data)) | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :601:27, :609:33, :611:{12,13}, :613:{42,73}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:611:12
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n");	// rob.scala:611:12
        if (`STOP_COND_)	// rob.scala:611:12
          $fatal;	// rob.scala:611:12
      end
      if (~(~(will_commit_1 & ~_GEN_68[com_idx] & (|_rob_fflags_1_ext_R0_data))
            | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :547:70, :607:{12,13}, :608:{14,40}, :609:33
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:607:12
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n");	// rob.scala:607:12
        if (`STOP_COND_)	// rob.scala:607:12
          $fatal;	// rob.scala:607:12
      end
      if (~(~(_fflags_val_1_T & (_GEN_61[com_idx] | _GEN_62[com_idx])
              & (|_rob_fflags_1_ext_R0_data)) | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :601:27, :609:33, :611:{12,13}, :613:{42,73}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:611:12
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n");	// rob.scala:611:12
        if (`STOP_COND_)	// rob.scala:611:12
          $fatal;	// rob.scala:611:12
      end
      if (~(~(will_commit_2 & ~_GEN_103[com_idx] & (|_rob_fflags_2_ext_R0_data))
            | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :547:70, :607:{12,13}, :608:{14,40}, :609:33
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:607:12
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n");	// rob.scala:607:12
        if (`STOP_COND_)	// rob.scala:607:12
          $fatal;	// rob.scala:607:12
      end
      if (~(~(_fflags_val_2_T & (_GEN_96[com_idx] | _GEN_97[com_idx])
              & (|_rob_fflags_2_ext_R0_data)) | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :601:27, :609:33, :611:{12,13}, :613:{42,73}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:611:12
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n");	// rob.scala:611:12
        if (`STOP_COND_)	// rob.scala:611:12
          $fatal;	// rob.scala:611:12
      end
      if (~(~(will_commit_3 & ~_GEN_138[com_idx] & (|_rob_fflags_3_ext_R0_data))
            | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :547:70, :607:{12,13}, :608:{14,40}, :609:33
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:607:12
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n");	// rob.scala:607:12
        if (`STOP_COND_)	// rob.scala:607:12
          $fatal;	// rob.scala:607:12
      end
      if (~(~(_fflags_val_3_T & (_GEN_131[com_idx] | _GEN_132[com_idx])
              & (|_rob_fflags_3_ext_R0_data)) | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :601:27, :609:33, :611:{12,13}, :613:{42,73}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:611:12
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n");	// rob.scala:611:12
        if (`STOP_COND_)	// rob.scala:611:12
          $fatal;	// rob.scala:611:12
      end
      if (~(~(exception_thrown & ~r_xcpt_val) | reset)) begin	// rob.scala:258:33, :545:85, :658:{10,11,30,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:658:10
          $error("Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:658 assert (!(exception_thrown && !r_xcpt_val),\n");	// rob.scala:658:10
        if (`STOP_COND_)	// rob.scala:658:10
          $fatal;	// rob.scala:658:10
      end
      if (~(~(empty & r_xcpt_val) | reset)) begin	// rob.scala:258:33, :661:{10,11,19}, :788:41
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:661:10
          $error("Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:661 assert (!(empty && r_xcpt_val),\n");	// rob.scala:661:10
        if (`STOP_COND_)	// rob.scala:661:10
          $fatal;	// rob.scala:661:10
      end
      if (~(~(exception_thrown & r_xcpt_uop_rob_idx[6:2] != rob_head) | reset)) begin	// rob.scala:224:29, :236:31, :259:29, :268:25, :545:85, :664:{10,11,34,68}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:664:10
          $error("Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:664 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n");	// rob.scala:664:10
        if (`STOP_COND_)	// rob.scala:664:10
          $fatal;	// rob.scala:664:10
      end
      if (~(_GEN_144 ^ rob_head_idx < rob_tail_idx ^ rob_pnr_idx >= rob_tail_idx
            | rob_pnr_idx == rob_tail_idx | reset)) begin	// Cat.scala:30:58, rob.scala:740:{9,10,75}, util.scala:363:{52,64,78}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:740:9
          $error("Assertion failed\n    at rob.scala:740 assert(!IsOlder(rob_pnr_idx, rob_head_idx, rob_tail_idx) || rob_pnr_idx === rob_tail_idx)\n");	// rob.scala:740:9
        if (`STOP_COND_)	// rob.scala:740:9
          $fatal;	// rob.scala:740:9
      end
      if (~(rob_tail_idx < rob_head_idx ^ _GEN_144 ^ rob_tail_idx >= rob_pnr_idx | full
            | reset)) begin	// Cat.scala:30:58, rob.scala:743:{9,10}, :787:39, util.scala:363:{52,64}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:743:9
          $error("Assertion failed\n    at rob.scala:743 assert(!IsOlder(rob_tail_idx, rob_pnr_idx, rob_head_idx) || full)\n");	// rob.scala:743:9
        if (`STOP_COND_)	// rob.scala:743:9
          $fatal;	// rob.scala:743:9
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire             _GEN_146 =
    _io_commit_rollback_T_3 & (rob_tail != rob_head | maybe_full);	// rob.scala:224:29, :228:29, :236:31, :239:29, :750:{34,47,60}
  wire             rob_deq = _GEN_146 | finished_committing_row;	// rob.scala:685:59, :688:34, :750:{34,76}, :754:13
  assign full = rob_tail == rob_head & maybe_full;	// rob.scala:224:29, :228:29, :239:29, :787:{26,39}
  assign empty =
    _empty_T
    & {rob_head_vals_3, rob_head_vals_2, rob_head_vals_1, rob_head_vals_0} == 4'h0;	// rob.scala:287:15, :398:49, :686:33, :788:{41,59,66}
  reg              REG;	// rob.scala:808:30
  reg              REG_1;	// rob.scala:808:22
  reg              REG_2;	// rob.scala:824:22
  reg              io_com_load_is_at_rob_head_REG;	// rob.scala:865:40
  always @(posedge clock) begin
    automatic logic             _GEN_147;	// rob.scala:324:31
    automatic logic             _GEN_148;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_149;	// rob.scala:324:31
    automatic logic             _GEN_150;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_151;	// rob.scala:324:31
    automatic logic             _GEN_152;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_153;	// rob.scala:324:31
    automatic logic             _GEN_154;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_155;	// rob.scala:324:31
    automatic logic             _GEN_156;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_157;	// rob.scala:324:31
    automatic logic             _GEN_158;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_159;	// rob.scala:324:31
    automatic logic             _GEN_160;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_161;	// rob.scala:324:31
    automatic logic             _GEN_162;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_163;	// rob.scala:324:31
    automatic logic             _GEN_164;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_165;	// rob.scala:324:31
    automatic logic             _GEN_166;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_167;	// rob.scala:324:31
    automatic logic             _GEN_168;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_169;	// rob.scala:324:31
    automatic logic             _GEN_170;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_171;	// rob.scala:324:31
    automatic logic             _GEN_172;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_173;	// rob.scala:324:31
    automatic logic             _GEN_174;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_175;	// rob.scala:324:31
    automatic logic             _GEN_176;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_177;	// rob.scala:324:31
    automatic logic             _GEN_178;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_179;	// rob.scala:324:31
    automatic logic             _GEN_180;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_181;	// rob.scala:324:31
    automatic logic             _GEN_182;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_183;	// rob.scala:324:31
    automatic logic             _GEN_184;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_185;	// rob.scala:324:31
    automatic logic             _GEN_186;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_187;	// rob.scala:324:31
    automatic logic             _GEN_188;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_189;	// rob.scala:324:31
    automatic logic             _GEN_190;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_191;	// rob.scala:324:31
    automatic logic             _GEN_192;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_193;	// rob.scala:324:31
    automatic logic             _GEN_194;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_195;	// rob.scala:324:31
    automatic logic             _GEN_196;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_197;	// rob.scala:324:31
    automatic logic             _GEN_198;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_199;	// rob.scala:324:31
    automatic logic             _GEN_200;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_201;	// rob.scala:324:31
    automatic logic             _GEN_202;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_203;	// rob.scala:324:31
    automatic logic             _GEN_204;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_205;	// rob.scala:324:31
    automatic logic             _GEN_206;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_207;	// rob.scala:324:31
    automatic logic             _GEN_208;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_209;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _rob_bsy_T =
      io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei;	// rob.scala:325:60
    automatic logic             _GEN_210;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_211;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_212;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_213;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_214;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_215;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_216;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_217;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_218;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_219;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_220;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_221;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_222;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_223;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_224;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_225;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_226;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_227;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_228;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_229;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_230;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_231;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_232;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_233;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_234;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_235;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_236;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_237;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_238;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_239;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_240;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_241;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _rob_unsafe_T_4 =
      io_enq_uops_0_uses_ldq | io_enq_uops_0_uses_stq & ~io_enq_uops_0_is_fence
      | io_enq_uops_0_is_br | io_enq_uops_0_is_jalr;	// micro-op.scala:152:{48,51,71}
    automatic logic             _GEN_242;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_243;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_244;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_245;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_246;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_247;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_248;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_249;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_250;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_251;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_252;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_253;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_254;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_255;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_256;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_257;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_258;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_259;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_260;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_261;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_262;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_263;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_264;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_265;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_266;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_267;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_268;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_269;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_270;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_271;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_272;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_273;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_274 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_275 = _GEN_0 & _GEN_274;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_276 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_277 = _GEN_0 & _GEN_276;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_278 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_279 = _GEN_0 & _GEN_278;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_280 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_281 = _GEN_0 & _GEN_280;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_282 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_283 = _GEN_0 & _GEN_282;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_284 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_285 = _GEN_0 & _GEN_284;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_286 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_287 = _GEN_0 & _GEN_286;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_288 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_289 = _GEN_0 & _GEN_288;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_290 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_291 = _GEN_0 & _GEN_290;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_292 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_293 = _GEN_0 & _GEN_292;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_294 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_295 = _GEN_0 & _GEN_294;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_296 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_297 = _GEN_0 & _GEN_296;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_298 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_299 = _GEN_0 & _GEN_298;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_300 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_301 = _GEN_0 & _GEN_300;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_302 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_303 = _GEN_0 & _GEN_302;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_304 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_305 = _GEN_0 & _GEN_304;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_306 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_307 = _GEN_0 & _GEN_306;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_308 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_309 = _GEN_0 & _GEN_308;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_310 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_311 = _GEN_0 & _GEN_310;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_312 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_313 = _GEN_0 & _GEN_312;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_314 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_315 = _GEN_0 & _GEN_314;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_316 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_317 = _GEN_0 & _GEN_316;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_318 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_319 = _GEN_0 & _GEN_318;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_320 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_321 = _GEN_0 & _GEN_320;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_322 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_323 = _GEN_0 & _GEN_322;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_324 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_325 = _GEN_0 & _GEN_324;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_326 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_327 = _GEN_0 & _GEN_326;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_328 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_329 = _GEN_0 & _GEN_328;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_330 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_331 = _GEN_0 & _GEN_330;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_332 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_333 = _GEN_0 & _GEN_332;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_334 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_335 = _GEN_0 & _GEN_334;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_336 =
      _GEN_0 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_337 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_338 = _GEN_337 | _GEN_275;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_339;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_340 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_341 = _GEN_340 | _GEN_277;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_342;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_343 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_344 = _GEN_343 | _GEN_279;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_345;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_346 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_347 = _GEN_346 | _GEN_281;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_348;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_349 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_350 = _GEN_349 | _GEN_283;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_351;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_352 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_353 = _GEN_352 | _GEN_285;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_354;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_355 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_356 = _GEN_355 | _GEN_287;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_357;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_358 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_359 = _GEN_358 | _GEN_289;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_360;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_361 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_362 = _GEN_361 | _GEN_291;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_363;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_364 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_365 = _GEN_364 | _GEN_293;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_366;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_367 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_368 = _GEN_367 | _GEN_295;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_369;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_370 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_371 = _GEN_370 | _GEN_297;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_372;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_373 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_374 = _GEN_373 | _GEN_299;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_375;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_376 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_377 = _GEN_376 | _GEN_301;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_378;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_379 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_380 = _GEN_379 | _GEN_303;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_381;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_382 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_383 = _GEN_382 | _GEN_305;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_384;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_385 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_386 = _GEN_385 | _GEN_307;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_387;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_388 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_389 = _GEN_388 | _GEN_309;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_390;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_391 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_392 = _GEN_391 | _GEN_311;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_393;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_394 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_395 = _GEN_394 | _GEN_313;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_396;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_397 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_398 = _GEN_397 | _GEN_315;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_399;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_400 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_401 = _GEN_400 | _GEN_317;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_402;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_403 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_404 = _GEN_403 | _GEN_319;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_405;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_406 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_407 = _GEN_406 | _GEN_321;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_408;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_409 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_410 = _GEN_409 | _GEN_323;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_411;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_412 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_413 = _GEN_412 | _GEN_325;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_414;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_415 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_416 = _GEN_415 | _GEN_327;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_417;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_418 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_419 = _GEN_418 | _GEN_329;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_420;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_421 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_422 = _GEN_421 | _GEN_331;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_423;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_424 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_425 = _GEN_424 | _GEN_333;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_426;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_427 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_428 = _GEN_427 | _GEN_335;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_429;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_430 =
      (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_336;	// rob.scala:236:31, :268:25, :323:29, :346:69, :347:31
    automatic logic             _GEN_431;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_432;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_433;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_434;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_435;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_436;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_437;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_438;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_439;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_440;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_441;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_442;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_443;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_444;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_445;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_446;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_447;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_448;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_449;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_450;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_451;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_452;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_453;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_454;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_455;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_456;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_457;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_458;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_459;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_460;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_461;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_462;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_463;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_464 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_465 = _GEN_2 & _GEN_464;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_466 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_467 = _GEN_2 & _GEN_466;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_468 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_469 = _GEN_2 & _GEN_468;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_470 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_471 = _GEN_2 & _GEN_470;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_472 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_473 = _GEN_2 & _GEN_472;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_474 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_475 = _GEN_2 & _GEN_474;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_476 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_477 = _GEN_2 & _GEN_476;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_478 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_479 = _GEN_2 & _GEN_478;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_480 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_481 = _GEN_2 & _GEN_480;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_482 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_483 = _GEN_2 & _GEN_482;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_484 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_485 = _GEN_2 & _GEN_484;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_486 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_487 = _GEN_2 & _GEN_486;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_488 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_489 = _GEN_2 & _GEN_488;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_490 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_491 = _GEN_2 & _GEN_490;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_492 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_493 = _GEN_2 & _GEN_492;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_494 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_495 = _GEN_2 & _GEN_494;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_496 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_497 = _GEN_2 & _GEN_496;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_498 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_499 = _GEN_2 & _GEN_498;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_500 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_501 = _GEN_2 & _GEN_500;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_502 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_503 = _GEN_2 & _GEN_502;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_504 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_505 = _GEN_2 & _GEN_504;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_506 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_507 = _GEN_2 & _GEN_506;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_508 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_509 = _GEN_2 & _GEN_508;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_510 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_511 = _GEN_2 & _GEN_510;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_512 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_513 = _GEN_2 & _GEN_512;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_514 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_515 = _GEN_2 & _GEN_514;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_516 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_517 = _GEN_2 & _GEN_516;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_518 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_519 = _GEN_2 & _GEN_518;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_520 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_521 = _GEN_2 & _GEN_520;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_522 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_523 = _GEN_2 & _GEN_522;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_524 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_525 = _GEN_2 & _GEN_524;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_526 =
      _GEN_2 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_527 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_528 = _GEN_527 | _GEN_465;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_529;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_530 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_531 = _GEN_530 | _GEN_467;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_532;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_533 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_534 = _GEN_533 | _GEN_469;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_535;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_536 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_537 = _GEN_536 | _GEN_471;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_538;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_539 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_540 = _GEN_539 | _GEN_473;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_541;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_542 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_543 = _GEN_542 | _GEN_475;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_544;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_545 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_546 = _GEN_545 | _GEN_477;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_547;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_548 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_549 = _GEN_548 | _GEN_479;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_550;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_551 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_552 = _GEN_551 | _GEN_481;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_553;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_554 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_555 = _GEN_554 | _GEN_483;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_556;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_557 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_558 = _GEN_557 | _GEN_485;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_559;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_560 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_561 = _GEN_560 | _GEN_487;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_562;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_563 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_564 = _GEN_563 | _GEN_489;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_565;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_566 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_567 = _GEN_566 | _GEN_491;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_568;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_569 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_570 = _GEN_569 | _GEN_493;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_571;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_572 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_573 = _GEN_572 | _GEN_495;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_574;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_575 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_576 = _GEN_575 | _GEN_497;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_577;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_578 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_579 = _GEN_578 | _GEN_499;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_580;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_581 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_582 = _GEN_581 | _GEN_501;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_583;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_584 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_585 = _GEN_584 | _GEN_503;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_586;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_587 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_588 = _GEN_587 | _GEN_505;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_589;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_590 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_591 = _GEN_590 | _GEN_507;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_592;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_593 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_594 = _GEN_593 | _GEN_509;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_595;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_596 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_597 = _GEN_596 | _GEN_511;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_598;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_599 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_600 = _GEN_599 | _GEN_513;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_601;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_602 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_603 = _GEN_602 | _GEN_515;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_604;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_605 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_606 = _GEN_605 | _GEN_517;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_607;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_608 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_609 = _GEN_608 | _GEN_519;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_610;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_611 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_612 = _GEN_611 | _GEN_521;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_613;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_614 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_615 = _GEN_614 | _GEN_523;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_616;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_617 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_618 = _GEN_617 | _GEN_525;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_619;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_620 =
      (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_526;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_621;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_622;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_623;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_624;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_625;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_626;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_627;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_628;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_629;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_630;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_631;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_632;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_633;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_634;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_635;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_636;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_637;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_638;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_639;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_640;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_641;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_642;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_643;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_644;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_645;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_646;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_647;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_648;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_649;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_650;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_651;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_652;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_653;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_654 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_655 = _GEN_4 & _GEN_654;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_656 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_657 = _GEN_4 & _GEN_656;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_658 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_659 = _GEN_4 & _GEN_658;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_660 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_661 = _GEN_4 & _GEN_660;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_662 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_663 = _GEN_4 & _GEN_662;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_664 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_665 = _GEN_4 & _GEN_664;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_666 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_667 = _GEN_4 & _GEN_666;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_668 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_669 = _GEN_4 & _GEN_668;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_670 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_671 = _GEN_4 & _GEN_670;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_672 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_673 = _GEN_4 & _GEN_672;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_674 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_675 = _GEN_4 & _GEN_674;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_676 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_677 = _GEN_4 & _GEN_676;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_678 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_679 = _GEN_4 & _GEN_678;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_680 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_681 = _GEN_4 & _GEN_680;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_682 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_683 = _GEN_4 & _GEN_682;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_684 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_685 = _GEN_4 & _GEN_684;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_686 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_687 = _GEN_4 & _GEN_686;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_688 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_689 = _GEN_4 & _GEN_688;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_690 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_691 = _GEN_4 & _GEN_690;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_692 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_693 = _GEN_4 & _GEN_692;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_694 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_695 = _GEN_4 & _GEN_694;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_696 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_697 = _GEN_4 & _GEN_696;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_698 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_699 = _GEN_4 & _GEN_698;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_700 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_701 = _GEN_4 & _GEN_700;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_702 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_703 = _GEN_4 & _GEN_702;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_704 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_705 = _GEN_4 & _GEN_704;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_706 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_707 = _GEN_4 & _GEN_706;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_708 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_709 = _GEN_4 & _GEN_708;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_710 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_711 = _GEN_4 & _GEN_710;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_712 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_713 = _GEN_4 & _GEN_712;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_714 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_715 = _GEN_4 & _GEN_714;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_716 =
      _GEN_4 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_717 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_718 = _GEN_717 | _GEN_655;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_719;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_720 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_721 = _GEN_720 | _GEN_657;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_722;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_723 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_724 = _GEN_723 | _GEN_659;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_725;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_726 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_727 = _GEN_726 | _GEN_661;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_728;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_729 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_730 = _GEN_729 | _GEN_663;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_731;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_732 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_733 = _GEN_732 | _GEN_665;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_734;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_735 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_736 = _GEN_735 | _GEN_667;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_737;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_738 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_739 = _GEN_738 | _GEN_669;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_740;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_741 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_742 = _GEN_741 | _GEN_671;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_743;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_744 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_745 = _GEN_744 | _GEN_673;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_746;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_747 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_748 = _GEN_747 | _GEN_675;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_749;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_750 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_751 = _GEN_750 | _GEN_677;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_752;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_753 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_754 = _GEN_753 | _GEN_679;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_755;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_756 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_757 = _GEN_756 | _GEN_681;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_758;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_759 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_760 = _GEN_759 | _GEN_683;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_761;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_762 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_763 = _GEN_762 | _GEN_685;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_764;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_765 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_766 = _GEN_765 | _GEN_687;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_767;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_768 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_769 = _GEN_768 | _GEN_689;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_770;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_771 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_772 = _GEN_771 | _GEN_691;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_773;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_774 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_775 = _GEN_774 | _GEN_693;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_776;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_777 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_778 = _GEN_777 | _GEN_695;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_779;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_780 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_781 = _GEN_780 | _GEN_697;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_782;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_783 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_784 = _GEN_783 | _GEN_699;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_785;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_786 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_787 = _GEN_786 | _GEN_701;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_788;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_789 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_790 = _GEN_789 | _GEN_703;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_791;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_792 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_793 = _GEN_792 | _GEN_705;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_794;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_795 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_796 = _GEN_795 | _GEN_707;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_797;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_798 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_799 = _GEN_798 | _GEN_709;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_800;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_801 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_802 = _GEN_801 | _GEN_711;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_803;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_804 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_805 = _GEN_804 | _GEN_713;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_806;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_807 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_808 = _GEN_807 | _GEN_715;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_809;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_810 =
      (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_716;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_811;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_812;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_813;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_814;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_815;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_816;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_817;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_818;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_819;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_820;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_821;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_822;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_823;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_824;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_825;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_826;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_827;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_828;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_829;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_830;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_831;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_832;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_833;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_834;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_835;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_836;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_837;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_838;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_839;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_840;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_841;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_842;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_843;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_844 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_845 = _GEN_6 & _GEN_844;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_846 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_847 = _GEN_6 & _GEN_846;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_848 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_849 = _GEN_6 & _GEN_848;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_850 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_851 = _GEN_6 & _GEN_850;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_852 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_853 = _GEN_6 & _GEN_852;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_854 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_855 = _GEN_6 & _GEN_854;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_856 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_857 = _GEN_6 & _GEN_856;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_858 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_859 = _GEN_6 & _GEN_858;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_860 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_861 = _GEN_6 & _GEN_860;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_862 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_863 = _GEN_6 & _GEN_862;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_864 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_865 = _GEN_6 & _GEN_864;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_866 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_867 = _GEN_6 & _GEN_866;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_868 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_869 = _GEN_6 & _GEN_868;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_870 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_871 = _GEN_6 & _GEN_870;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_872 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_873 = _GEN_6 & _GEN_872;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_874 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_875 = _GEN_6 & _GEN_874;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_876 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_877 = _GEN_6 & _GEN_876;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_878 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_879 = _GEN_6 & _GEN_878;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_880 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_881 = _GEN_6 & _GEN_880;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_882 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_883 = _GEN_6 & _GEN_882;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_884 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_885 = _GEN_6 & _GEN_884;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_886 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_887 = _GEN_6 & _GEN_886;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_888 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_889 = _GEN_6 & _GEN_888;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_890 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_891 = _GEN_6 & _GEN_890;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_892 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_893 = _GEN_6 & _GEN_892;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_894 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_895 = _GEN_6 & _GEN_894;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_896 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_897 = _GEN_6 & _GEN_896;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_898 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_899 = _GEN_6 & _GEN_898;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_900 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_901 = _GEN_6 & _GEN_900;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_902 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_903 = _GEN_6 & _GEN_902;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_904 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_905 = _GEN_6 & _GEN_904;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_906 =
      _GEN_6 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_907 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_908 = _GEN_907 | _GEN_845;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_909;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_910 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_911 = _GEN_910 | _GEN_847;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_912;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_913 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_914 = _GEN_913 | _GEN_849;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_915;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_916 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_917 = _GEN_916 | _GEN_851;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_918;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_919 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_920 = _GEN_919 | _GEN_853;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_921;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_922 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_923 = _GEN_922 | _GEN_855;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_924;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_925 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_926 = _GEN_925 | _GEN_857;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_927;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_928 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_929 = _GEN_928 | _GEN_859;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_930;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_931 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_932 = _GEN_931 | _GEN_861;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_933;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_934 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_935 = _GEN_934 | _GEN_863;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_936;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_937 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_938 = _GEN_937 | _GEN_865;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_939;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_940 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_941 = _GEN_940 | _GEN_867;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_942;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_943 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_944 = _GEN_943 | _GEN_869;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_945;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_946 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_947 = _GEN_946 | _GEN_871;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_948;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_949 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_950 = _GEN_949 | _GEN_873;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_951;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_952 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_953 = _GEN_952 | _GEN_875;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_954;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_955 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_956 = _GEN_955 | _GEN_877;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_957;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_958 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_959 = _GEN_958 | _GEN_879;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_960;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_961 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_962 = _GEN_961 | _GEN_881;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_963;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_964 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_965 = _GEN_964 | _GEN_883;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_966;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_967 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_968 = _GEN_967 | _GEN_885;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_969;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_970 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_971 = _GEN_970 | _GEN_887;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_972;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_973 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_974 = _GEN_973 | _GEN_889;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_975;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_976 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_977 = _GEN_976 | _GEN_891;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_978;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_979 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_980 = _GEN_979 | _GEN_893;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_981;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_982 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_983 = _GEN_982 | _GEN_895;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_984;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_985 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_986 = _GEN_985 | _GEN_897;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_987;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_988 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_989 = _GEN_988 | _GEN_899;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_990;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_991 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_992 = _GEN_991 | _GEN_901;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_993;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_994 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_995 = _GEN_994 | _GEN_903;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_996;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_997 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_998 = _GEN_997 | _GEN_905;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_999;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1000 =
      (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_906;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_1001;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1002;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1003;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1004;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1005;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1006;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1007;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1008;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1009;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1010;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1011;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1012;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1013;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1014;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1015;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1016;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1017;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1018;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1019;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1020;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1021;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1022;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1023;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1024;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1025;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1026;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1027;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1028;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1029;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1030;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1031;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1032;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1033;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1034 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_1035 = _GEN_8 & _GEN_1034;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1036 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1037 = _GEN_8 & _GEN_1036;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1038 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1039 = _GEN_8 & _GEN_1038;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1040 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1041 = _GEN_8 & _GEN_1040;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1042 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1043 = _GEN_8 & _GEN_1042;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1044 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1045 = _GEN_8 & _GEN_1044;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1046 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1047 = _GEN_8 & _GEN_1046;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1048 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1049 = _GEN_8 & _GEN_1048;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1050 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1051 = _GEN_8 & _GEN_1050;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1052 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1053 = _GEN_8 & _GEN_1052;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1054 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1055 = _GEN_8 & _GEN_1054;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1056 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1057 = _GEN_8 & _GEN_1056;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1058 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1059 = _GEN_8 & _GEN_1058;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1060 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1061 = _GEN_8 & _GEN_1060;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1062 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1063 = _GEN_8 & _GEN_1062;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1064 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1065 = _GEN_8 & _GEN_1064;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1066 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1067 = _GEN_8 & _GEN_1066;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1068 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1069 = _GEN_8 & _GEN_1068;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1070 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1071 = _GEN_8 & _GEN_1070;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1072 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1073 = _GEN_8 & _GEN_1072;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1074 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1075 = _GEN_8 & _GEN_1074;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1076 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1077 = _GEN_8 & _GEN_1076;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1078 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1079 = _GEN_8 & _GEN_1078;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1080 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1081 = _GEN_8 & _GEN_1080;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1082 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1083 = _GEN_8 & _GEN_1082;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1084 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1085 = _GEN_8 & _GEN_1084;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1086 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1087 = _GEN_8 & _GEN_1086;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1088 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1089 = _GEN_8 & _GEN_1088;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1090 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1091 = _GEN_8 & _GEN_1090;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1092 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1093 = _GEN_8 & _GEN_1092;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1094 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1095 = _GEN_8 & _GEN_1094;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1096 =
      _GEN_8 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_1097 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :347:31
    automatic logic             _GEN_1098 = _GEN_1097 | _GEN_1035;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1099;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1100 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1101 = _GEN_1100 | _GEN_1037;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1102;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1103 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1104 = _GEN_1103 | _GEN_1039;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1105;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1106 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1107 = _GEN_1106 | _GEN_1041;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1108;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1109 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1110 = _GEN_1109 | _GEN_1043;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1111;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1112 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1113 = _GEN_1112 | _GEN_1045;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1114;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1115 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1116 = _GEN_1115 | _GEN_1047;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1117;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1118 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1119 = _GEN_1118 | _GEN_1049;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1120;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1121 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1122 = _GEN_1121 | _GEN_1051;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1123;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1124 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1125 = _GEN_1124 | _GEN_1053;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1126;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1127 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1128 = _GEN_1127 | _GEN_1055;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1129;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1130 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1131 = _GEN_1130 | _GEN_1057;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1132;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1133 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1134 = _GEN_1133 | _GEN_1059;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1135;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1136 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1137 = _GEN_1136 | _GEN_1061;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1138;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1139 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1140 = _GEN_1139 | _GEN_1063;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1141;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1142 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1143 = _GEN_1142 | _GEN_1065;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1144;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1145 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1146 = _GEN_1145 | _GEN_1067;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1147;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1148 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1149 = _GEN_1148 | _GEN_1069;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1150;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1151 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1152 = _GEN_1151 | _GEN_1071;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1153;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1154 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1155 = _GEN_1154 | _GEN_1073;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1156;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1157 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1158 = _GEN_1157 | _GEN_1075;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1159;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1160 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1161 = _GEN_1160 | _GEN_1077;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1162;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1163 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1164 = _GEN_1163 | _GEN_1079;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1165;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1166 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1167 = _GEN_1166 | _GEN_1081;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1168;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1169 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1170 = _GEN_1169 | _GEN_1083;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1171;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1172 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1173 = _GEN_1172 | _GEN_1085;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1174;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1175 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1176 = _GEN_1175 | _GEN_1087;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1177;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1178 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1179 = _GEN_1178 | _GEN_1089;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1180;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1181 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1182 = _GEN_1181 | _GEN_1091;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1183;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1184 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1185 = _GEN_1184 | _GEN_1093;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1186;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1187 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_1188 = _GEN_1187 | _GEN_1095;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1189;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1190 =
      (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1096;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_1191;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1192;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1193;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1194;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1195;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1196;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1197;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1198;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1199;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1200;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1201;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1202;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1203;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1204;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1205;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1206;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1207;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1208;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1209;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1210;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1211;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1212;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1213;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1214;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1215;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1216;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1217;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1218;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1219;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1220;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1221;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1222;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1223;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1224 = io_lsu_clr_bsy_0_bits[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :363:26
    automatic logic             _GEN_1225 = _GEN_10 & _GEN_1224;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1226 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1227 = _GEN_10 & _GEN_1226;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1228 = io_lsu_clr_bsy_0_bits[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1229 = _GEN_10 & _GEN_1228;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1230 = io_lsu_clr_bsy_0_bits[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1231 = _GEN_10 & _GEN_1230;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1232 = io_lsu_clr_bsy_0_bits[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1233 = _GEN_10 & _GEN_1232;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1234 = io_lsu_clr_bsy_0_bits[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1235 = _GEN_10 & _GEN_1234;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1236 = io_lsu_clr_bsy_0_bits[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1237 = _GEN_10 & _GEN_1236;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1238 = io_lsu_clr_bsy_0_bits[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1239 = _GEN_10 & _GEN_1238;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1240 = io_lsu_clr_bsy_0_bits[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1241 = _GEN_10 & _GEN_1240;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1242 = io_lsu_clr_bsy_0_bits[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1243 = _GEN_10 & _GEN_1242;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1244 = io_lsu_clr_bsy_0_bits[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1245 = _GEN_10 & _GEN_1244;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1246 = io_lsu_clr_bsy_0_bits[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1247 = _GEN_10 & _GEN_1246;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1248 = io_lsu_clr_bsy_0_bits[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1249 = _GEN_10 & _GEN_1248;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1250 = io_lsu_clr_bsy_0_bits[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1251 = _GEN_10 & _GEN_1250;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1252 = io_lsu_clr_bsy_0_bits[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1253 = _GEN_10 & _GEN_1252;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1254 = io_lsu_clr_bsy_0_bits[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1255 = _GEN_10 & _GEN_1254;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1256 = io_lsu_clr_bsy_0_bits[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1257 = _GEN_10 & _GEN_1256;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1258 = io_lsu_clr_bsy_0_bits[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1259 = _GEN_10 & _GEN_1258;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1260 = io_lsu_clr_bsy_0_bits[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1261 = _GEN_10 & _GEN_1260;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1262 = io_lsu_clr_bsy_0_bits[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1263 = _GEN_10 & _GEN_1262;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1264 = io_lsu_clr_bsy_0_bits[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1265 = _GEN_10 & _GEN_1264;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1266 = io_lsu_clr_bsy_0_bits[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1267 = _GEN_10 & _GEN_1266;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1268 = io_lsu_clr_bsy_0_bits[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1269 = _GEN_10 & _GEN_1268;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1270 = io_lsu_clr_bsy_0_bits[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1271 = _GEN_10 & _GEN_1270;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1272 = io_lsu_clr_bsy_0_bits[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1273 = _GEN_10 & _GEN_1272;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1274 = io_lsu_clr_bsy_0_bits[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1275 = _GEN_10 & _GEN_1274;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1276 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1277 = _GEN_10 & _GEN_1276;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1278 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1279 = _GEN_10 & _GEN_1278;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1280 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1281 = _GEN_10 & _GEN_1280;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1282 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1283 = _GEN_10 & _GEN_1282;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1284 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1285 = _GEN_10 & _GEN_1284;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1286 = _GEN_10 & (&(io_lsu_clr_bsy_0_bits[6:2]));	// rob.scala:236:31, :268:25, :346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_1287 = io_lsu_clr_bsy_1_bits[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :363:26
    automatic logic             _GEN_1288 = _GEN_1287 | _GEN_1225;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1289 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1290 = _GEN_1289 | _GEN_1227;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1291 = io_lsu_clr_bsy_1_bits[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1292 = _GEN_1291 | _GEN_1229;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1293 = io_lsu_clr_bsy_1_bits[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1294 = _GEN_1293 | _GEN_1231;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1295 = io_lsu_clr_bsy_1_bits[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1296 = _GEN_1295 | _GEN_1233;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1297 = io_lsu_clr_bsy_1_bits[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1298 = _GEN_1297 | _GEN_1235;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1299 = io_lsu_clr_bsy_1_bits[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1300 = _GEN_1299 | _GEN_1237;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1301 = io_lsu_clr_bsy_1_bits[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1302 = _GEN_1301 | _GEN_1239;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1303 = io_lsu_clr_bsy_1_bits[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1304 = _GEN_1303 | _GEN_1241;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1305 = io_lsu_clr_bsy_1_bits[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1306 = _GEN_1305 | _GEN_1243;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1307 = io_lsu_clr_bsy_1_bits[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1308 = _GEN_1307 | _GEN_1245;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1309 = io_lsu_clr_bsy_1_bits[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1310 = _GEN_1309 | _GEN_1247;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1311 = io_lsu_clr_bsy_1_bits[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1312 = _GEN_1311 | _GEN_1249;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1313 = io_lsu_clr_bsy_1_bits[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1314 = _GEN_1313 | _GEN_1251;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1315 = io_lsu_clr_bsy_1_bits[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1316 = _GEN_1315 | _GEN_1253;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1317 = io_lsu_clr_bsy_1_bits[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1318 = _GEN_1317 | _GEN_1255;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1319 = io_lsu_clr_bsy_1_bits[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1320 = _GEN_1319 | _GEN_1257;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1321 = io_lsu_clr_bsy_1_bits[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1322 = _GEN_1321 | _GEN_1259;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1323 = io_lsu_clr_bsy_1_bits[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1324 = _GEN_1323 | _GEN_1261;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1325 = io_lsu_clr_bsy_1_bits[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1326 = _GEN_1325 | _GEN_1263;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1327 = io_lsu_clr_bsy_1_bits[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1328 = _GEN_1327 | _GEN_1265;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1329 = io_lsu_clr_bsy_1_bits[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1330 = _GEN_1329 | _GEN_1267;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1331 = io_lsu_clr_bsy_1_bits[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1332 = _GEN_1331 | _GEN_1269;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1333 = io_lsu_clr_bsy_1_bits[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1334 = _GEN_1333 | _GEN_1271;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1335 = io_lsu_clr_bsy_1_bits[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1336 = _GEN_1335 | _GEN_1273;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1337 = io_lsu_clr_bsy_1_bits[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1338 = _GEN_1337 | _GEN_1275;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1339 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1340 = _GEN_1339 | _GEN_1277;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1341 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1342 = _GEN_1341 | _GEN_1279;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1343 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1344 = _GEN_1343 | _GEN_1281;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1345 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1346 = _GEN_1345 | _GEN_1283;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1347 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1348 = _GEN_1347 | _GEN_1285;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1349 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_1286;	// rob.scala:236:31, :268:25, :346:69, :361:75, :363:26
    automatic logic             _GEN_1350 = io_lsu_clr_bsy_2_bits[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :363:26
    automatic logic             _GEN_1351 = _GEN_13 & _GEN_1350;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1352 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1353 = _GEN_13 & _GEN_1352;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1354 = io_lsu_clr_bsy_2_bits[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1355 = _GEN_13 & _GEN_1354;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1356 = io_lsu_clr_bsy_2_bits[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1357 = _GEN_13 & _GEN_1356;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1358 = io_lsu_clr_bsy_2_bits[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1359 = _GEN_13 & _GEN_1358;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1360 = io_lsu_clr_bsy_2_bits[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1361 = _GEN_13 & _GEN_1360;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1362 = io_lsu_clr_bsy_2_bits[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1363 = _GEN_13 & _GEN_1362;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1364 = io_lsu_clr_bsy_2_bits[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1365 = _GEN_13 & _GEN_1364;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1366 = io_lsu_clr_bsy_2_bits[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1367 = _GEN_13 & _GEN_1366;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1368 = io_lsu_clr_bsy_2_bits[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1369 = _GEN_13 & _GEN_1368;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1370 = io_lsu_clr_bsy_2_bits[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1371 = _GEN_13 & _GEN_1370;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1372 = io_lsu_clr_bsy_2_bits[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1373 = _GEN_13 & _GEN_1372;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1374 = io_lsu_clr_bsy_2_bits[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1375 = _GEN_13 & _GEN_1374;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1376 = io_lsu_clr_bsy_2_bits[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1377 = _GEN_13 & _GEN_1376;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1378 = io_lsu_clr_bsy_2_bits[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1379 = _GEN_13 & _GEN_1378;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1380 = io_lsu_clr_bsy_2_bits[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1381 = _GEN_13 & _GEN_1380;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1382 = io_lsu_clr_bsy_2_bits[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1383 = _GEN_13 & _GEN_1382;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1384 = io_lsu_clr_bsy_2_bits[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1385 = _GEN_13 & _GEN_1384;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1386 = io_lsu_clr_bsy_2_bits[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1387 = _GEN_13 & _GEN_1386;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1388 = io_lsu_clr_bsy_2_bits[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1389 = _GEN_13 & _GEN_1388;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1390 = io_lsu_clr_bsy_2_bits[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1391 = _GEN_13 & _GEN_1390;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1392 = io_lsu_clr_bsy_2_bits[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1393 = _GEN_13 & _GEN_1392;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1394 = io_lsu_clr_bsy_2_bits[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1395 = _GEN_13 & _GEN_1394;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1396 = io_lsu_clr_bsy_2_bits[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1397 = _GEN_13 & _GEN_1396;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1398 = io_lsu_clr_bsy_2_bits[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1399 = _GEN_13 & _GEN_1398;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1400 = io_lsu_clr_bsy_2_bits[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1401 = _GEN_13 & _GEN_1400;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1402 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1403 = _GEN_13 & _GEN_1402;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1404 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1405 = _GEN_13 & _GEN_1404;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1406 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1407 = _GEN_13 & _GEN_1406;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1408 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1409 = _GEN_13 & _GEN_1408;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1410 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_1411 = _GEN_13 & _GEN_1410;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_1412 = _GEN_13 & (&(io_lsu_clr_bsy_2_bits[6:2]));	// rob.scala:236:31, :268:25, :361:{31,75}, :363:26
    automatic logic             _GEN_1413 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:236:31, :268:25, :391:59
    automatic logic             _GEN_1414 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1415 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1416 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1417 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1418 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1419 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1420 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1421 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1422 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1423 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1424 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1425 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1426 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1427 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1428 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1429 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1430 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1431 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1432 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1433 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1434 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1435 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1436 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1437 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1438 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1439 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1440 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1441 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1442 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1443 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_1444 = com_idx == 5'h0;	// rob.scala:236:{20,31}, :268:25, :434:30
    automatic logic             _GEN_1445;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1446 = com_idx == 5'h1;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1447;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1448 = com_idx == 5'h2;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1449;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1450 = com_idx == 5'h3;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1451;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1452 = com_idx == 5'h4;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1453;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1454 = com_idx == 5'h5;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1455;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1456 = com_idx == 5'h6;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1457;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1458 = com_idx == 5'h7;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1459;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1460 = com_idx == 5'h8;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1461;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1462 = com_idx == 5'h9;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1463;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1464 = com_idx == 5'hA;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1465;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1466 = com_idx == 5'hB;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1467;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1468 = com_idx == 5'hC;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1469;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1470 = com_idx == 5'hD;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1471;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1472 = com_idx == 5'hE;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1473;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1474 = com_idx == 5'hF;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1475;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1476 = com_idx == 5'h10;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1477;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1478 = com_idx == 5'h11;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1479;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1480 = com_idx == 5'h12;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1481;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1482 = com_idx == 5'h13;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1483;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1484 = com_idx == 5'h14;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1485;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1486 = com_idx == 5'h15;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1487;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1488 = com_idx == 5'h16;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1489;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1490 = com_idx == 5'h17;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1491;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1492 = com_idx == 5'h18;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1493;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1494 = com_idx == 5'h19;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1495;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1496 = com_idx == 5'h1A;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1497;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1498 = com_idx == 5'h1B;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1499;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1500 = com_idx == 5'h1C;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1501;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1502 = com_idx == 5'h1D;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1503;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1504 = com_idx == 5'h1E;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_1505;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1506;	// rob.scala:323:29, :433:20, :434:30
    automatic logic [19:0]      _GEN_1507;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1508;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1509;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1510;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1511;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1512;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1513;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1514;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1515;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1516;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1517;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1518;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1519;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1520;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1521;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1522;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1523;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1524;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1525;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1526;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1527;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1528;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1529;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1530;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1531;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1532;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1533;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1534;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1535;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1536;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1537;	// util.scala:118:51
    automatic logic [19:0]      _GEN_1538;	// util.scala:118:51
    automatic logic             _GEN_1539;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1540;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1541;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1542;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1543;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1544;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1545;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1546;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1547;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1548;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1549;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1550;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1551;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1552;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1553;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1554;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1555;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1556;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1557;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1558;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1559;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1560;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1561;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1562;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1563;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1564;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1565;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1566;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1567;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1568;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1569;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1570;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _rob_bsy_T_2 =
      io_enq_uops_1_is_fence | io_enq_uops_1_is_fencei;	// rob.scala:325:60
    automatic logic             _GEN_1571;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1572;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1573;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1574;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1575;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1576;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1577;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1578;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1579;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1580;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1581;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1582;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1583;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1584;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1585;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1586;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1587;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1588;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1589;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1590;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1591;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1592;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1593;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1594;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1595;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1596;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1597;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1598;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1599;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1600;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1601;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1602;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _rob_unsafe_T_9 =
      io_enq_uops_1_uses_ldq | io_enq_uops_1_uses_stq & ~io_enq_uops_1_is_fence
      | io_enq_uops_1_is_br | io_enq_uops_1_is_jalr;	// micro-op.scala:152:{48,51,71}
    automatic logic             _GEN_1603;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1604;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1605;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1606;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1607;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1608;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1609;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1610;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1611;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1612;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1613;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1614;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1615;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1616;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1617;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1618;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1619;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1620;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1621;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1622;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1623;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1624;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1625;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1626;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1627;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1628;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1629;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1630;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1631;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1632;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1633;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1634;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1635 = _GEN_35 & _GEN_274;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1636 = _GEN_35 & _GEN_276;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1637 = _GEN_35 & _GEN_278;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1638 = _GEN_35 & _GEN_280;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1639 = _GEN_35 & _GEN_282;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1640 = _GEN_35 & _GEN_284;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1641 = _GEN_35 & _GEN_286;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1642 = _GEN_35 & _GEN_288;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1643 = _GEN_35 & _GEN_290;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1644 = _GEN_35 & _GEN_292;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1645 = _GEN_35 & _GEN_294;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1646 = _GEN_35 & _GEN_296;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1647 = _GEN_35 & _GEN_298;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1648 = _GEN_35 & _GEN_300;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1649 = _GEN_35 & _GEN_302;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1650 = _GEN_35 & _GEN_304;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1651 = _GEN_35 & _GEN_306;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1652 = _GEN_35 & _GEN_308;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1653 = _GEN_35 & _GEN_310;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1654 = _GEN_35 & _GEN_312;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1655 = _GEN_35 & _GEN_314;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1656 = _GEN_35 & _GEN_316;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1657 = _GEN_35 & _GEN_318;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1658 = _GEN_35 & _GEN_320;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1659 = _GEN_35 & _GEN_322;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1660 = _GEN_35 & _GEN_324;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1661 = _GEN_35 & _GEN_326;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1662 = _GEN_35 & _GEN_328;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1663 = _GEN_35 & _GEN_330;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1664 = _GEN_35 & _GEN_332;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1665 = _GEN_35 & _GEN_334;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1666 =
      _GEN_35 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1667 = _GEN_337 | _GEN_1635;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1668;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1669 = _GEN_340 | _GEN_1636;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1670;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1671 = _GEN_343 | _GEN_1637;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1672;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1673 = _GEN_346 | _GEN_1638;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1674;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1675 = _GEN_349 | _GEN_1639;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1676;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1677 = _GEN_352 | _GEN_1640;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1678;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1679 = _GEN_355 | _GEN_1641;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1680;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1681 = _GEN_358 | _GEN_1642;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1682;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1683 = _GEN_361 | _GEN_1643;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1684;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1685 = _GEN_364 | _GEN_1644;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1686;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1687 = _GEN_367 | _GEN_1645;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1688;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1689 = _GEN_370 | _GEN_1646;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1690;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1691 = _GEN_373 | _GEN_1647;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1692;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1693 = _GEN_376 | _GEN_1648;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1694;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1695 = _GEN_379 | _GEN_1649;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1696;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1697 = _GEN_382 | _GEN_1650;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1698;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1699 = _GEN_385 | _GEN_1651;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1700;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1701 = _GEN_388 | _GEN_1652;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1702;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1703 = _GEN_391 | _GEN_1653;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1704;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1705 = _GEN_394 | _GEN_1654;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1706;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1707 = _GEN_397 | _GEN_1655;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1708;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1709 = _GEN_400 | _GEN_1656;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1710;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1711 = _GEN_403 | _GEN_1657;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1712;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1713 = _GEN_406 | _GEN_1658;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1714;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1715 = _GEN_409 | _GEN_1659;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1716;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1717 = _GEN_412 | _GEN_1660;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1718;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1719 = _GEN_415 | _GEN_1661;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1720;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1721 = _GEN_418 | _GEN_1662;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1722;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1723 = _GEN_421 | _GEN_1663;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1724;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1725 = _GEN_424 | _GEN_1664;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1726;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1727 = _GEN_427 | _GEN_1665;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1728;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1729 =
      (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_1666;	// rob.scala:236:31, :268:25, :323:29, :346:69, :347:31
    automatic logic             _GEN_1730;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1731;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1732;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1733;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1734;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1735;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1736;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1737;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1738;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1739;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1740;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1741;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1742;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1743;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1744;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1745;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1746;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1747;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1748;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1749;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1750;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1751;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1752;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1753;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1754;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1755;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1756;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1757;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1758;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1759;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1760;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1761;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1762;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1763 = _GEN_37 & _GEN_464;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1764 = _GEN_37 & _GEN_466;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1765 = _GEN_37 & _GEN_468;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1766 = _GEN_37 & _GEN_470;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1767 = _GEN_37 & _GEN_472;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1768 = _GEN_37 & _GEN_474;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1769 = _GEN_37 & _GEN_476;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1770 = _GEN_37 & _GEN_478;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1771 = _GEN_37 & _GEN_480;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1772 = _GEN_37 & _GEN_482;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1773 = _GEN_37 & _GEN_484;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1774 = _GEN_37 & _GEN_486;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1775 = _GEN_37 & _GEN_488;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1776 = _GEN_37 & _GEN_490;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1777 = _GEN_37 & _GEN_492;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1778 = _GEN_37 & _GEN_494;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1779 = _GEN_37 & _GEN_496;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1780 = _GEN_37 & _GEN_498;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1781 = _GEN_37 & _GEN_500;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1782 = _GEN_37 & _GEN_502;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1783 = _GEN_37 & _GEN_504;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1784 = _GEN_37 & _GEN_506;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1785 = _GEN_37 & _GEN_508;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1786 = _GEN_37 & _GEN_510;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1787 = _GEN_37 & _GEN_512;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1788 = _GEN_37 & _GEN_514;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1789 = _GEN_37 & _GEN_516;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1790 = _GEN_37 & _GEN_518;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1791 = _GEN_37 & _GEN_520;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1792 = _GEN_37 & _GEN_522;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1793 = _GEN_37 & _GEN_524;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1794 =
      _GEN_37 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_1795 = _GEN_527 | _GEN_1763;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1796;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1797 = _GEN_530 | _GEN_1764;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1798;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1799 = _GEN_533 | _GEN_1765;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1800;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1801 = _GEN_536 | _GEN_1766;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1802;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1803 = _GEN_539 | _GEN_1767;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1804;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1805 = _GEN_542 | _GEN_1768;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1806;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1807 = _GEN_545 | _GEN_1769;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1808;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1809 = _GEN_548 | _GEN_1770;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1810;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1811 = _GEN_551 | _GEN_1771;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1812;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1813 = _GEN_554 | _GEN_1772;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1814;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1815 = _GEN_557 | _GEN_1773;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1816;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1817 = _GEN_560 | _GEN_1774;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1818;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1819 = _GEN_563 | _GEN_1775;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1820;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1821 = _GEN_566 | _GEN_1776;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1822;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1823 = _GEN_569 | _GEN_1777;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1824;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1825 = _GEN_572 | _GEN_1778;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1826;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1827 = _GEN_575 | _GEN_1779;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1828;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1829 = _GEN_578 | _GEN_1780;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1830;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1831 = _GEN_581 | _GEN_1781;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1832;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1833 = _GEN_584 | _GEN_1782;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1834;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1835 = _GEN_587 | _GEN_1783;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1836;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1837 = _GEN_590 | _GEN_1784;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1838;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1839 = _GEN_593 | _GEN_1785;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1840;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1841 = _GEN_596 | _GEN_1786;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1842;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1843 = _GEN_599 | _GEN_1787;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1844;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1845 = _GEN_602 | _GEN_1788;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1846;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1847 = _GEN_605 | _GEN_1789;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1848;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1849 = _GEN_608 | _GEN_1790;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1850;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1851 = _GEN_611 | _GEN_1791;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1852;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1853 = _GEN_614 | _GEN_1792;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1854;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1855 = _GEN_617 | _GEN_1793;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1856;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1857 =
      (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1794;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_1858;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1859;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1860;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1861;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1862;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1863;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1864;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1865;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1866;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1867;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1868;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1869;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1870;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1871;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1872;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1873;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1874;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1875;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1876;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1877;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1878;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1879;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1880;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1881;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1882;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1883;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1884;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1885;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1886;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1887;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1888;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1889;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1890;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1891 = _GEN_39 & _GEN_654;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1892 = _GEN_39 & _GEN_656;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1893 = _GEN_39 & _GEN_658;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1894 = _GEN_39 & _GEN_660;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1895 = _GEN_39 & _GEN_662;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1896 = _GEN_39 & _GEN_664;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1897 = _GEN_39 & _GEN_666;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1898 = _GEN_39 & _GEN_668;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1899 = _GEN_39 & _GEN_670;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1900 = _GEN_39 & _GEN_672;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1901 = _GEN_39 & _GEN_674;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1902 = _GEN_39 & _GEN_676;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1903 = _GEN_39 & _GEN_678;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1904 = _GEN_39 & _GEN_680;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1905 = _GEN_39 & _GEN_682;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1906 = _GEN_39 & _GEN_684;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1907 = _GEN_39 & _GEN_686;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1908 = _GEN_39 & _GEN_688;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1909 = _GEN_39 & _GEN_690;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1910 = _GEN_39 & _GEN_692;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1911 = _GEN_39 & _GEN_694;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1912 = _GEN_39 & _GEN_696;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1913 = _GEN_39 & _GEN_698;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1914 = _GEN_39 & _GEN_700;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1915 = _GEN_39 & _GEN_702;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1916 = _GEN_39 & _GEN_704;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1917 = _GEN_39 & _GEN_706;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1918 = _GEN_39 & _GEN_708;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1919 = _GEN_39 & _GEN_710;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1920 = _GEN_39 & _GEN_712;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1921 = _GEN_39 & _GEN_714;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1922 =
      _GEN_39 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_1923 = _GEN_717 | _GEN_1891;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1924;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1925 = _GEN_720 | _GEN_1892;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1926;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1927 = _GEN_723 | _GEN_1893;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1928;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1929 = _GEN_726 | _GEN_1894;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1930;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1931 = _GEN_729 | _GEN_1895;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1932;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1933 = _GEN_732 | _GEN_1896;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1934;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1935 = _GEN_735 | _GEN_1897;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1936;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1937 = _GEN_738 | _GEN_1898;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1938;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1939 = _GEN_741 | _GEN_1899;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1940;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1941 = _GEN_744 | _GEN_1900;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1942;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1943 = _GEN_747 | _GEN_1901;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1944;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1945 = _GEN_750 | _GEN_1902;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1946;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1947 = _GEN_753 | _GEN_1903;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1948;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1949 = _GEN_756 | _GEN_1904;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1950;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1951 = _GEN_759 | _GEN_1905;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1952;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1953 = _GEN_762 | _GEN_1906;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1954;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1955 = _GEN_765 | _GEN_1907;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1956;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1957 = _GEN_768 | _GEN_1908;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1958;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1959 = _GEN_771 | _GEN_1909;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1960;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1961 = _GEN_774 | _GEN_1910;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1962;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1963 = _GEN_777 | _GEN_1911;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1964;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1965 = _GEN_780 | _GEN_1912;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1966;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1967 = _GEN_783 | _GEN_1913;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1968;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1969 = _GEN_786 | _GEN_1914;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1970;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1971 = _GEN_789 | _GEN_1915;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1972;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1973 = _GEN_792 | _GEN_1916;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1974;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1975 = _GEN_795 | _GEN_1917;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1976;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1977 = _GEN_798 | _GEN_1918;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1978;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1979 = _GEN_801 | _GEN_1919;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1980;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1981 = _GEN_804 | _GEN_1920;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1982;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1983 = _GEN_807 | _GEN_1921;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1984;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1985 =
      (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1922;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_1986;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1987;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1988;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1989;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1990;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1991;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1992;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1993;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1994;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1995;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1996;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1997;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1998;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1999;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2000;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2001;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2002;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2003;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2004;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2005;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2006;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2007;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2008;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2009;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2010;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2011;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2012;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2013;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2014;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2015;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2016;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2017;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2018;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2019 = _GEN_41 & _GEN_844;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2020 = _GEN_41 & _GEN_846;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2021 = _GEN_41 & _GEN_848;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2022 = _GEN_41 & _GEN_850;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2023 = _GEN_41 & _GEN_852;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2024 = _GEN_41 & _GEN_854;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2025 = _GEN_41 & _GEN_856;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2026 = _GEN_41 & _GEN_858;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2027 = _GEN_41 & _GEN_860;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2028 = _GEN_41 & _GEN_862;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2029 = _GEN_41 & _GEN_864;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2030 = _GEN_41 & _GEN_866;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2031 = _GEN_41 & _GEN_868;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2032 = _GEN_41 & _GEN_870;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2033 = _GEN_41 & _GEN_872;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2034 = _GEN_41 & _GEN_874;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2035 = _GEN_41 & _GEN_876;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2036 = _GEN_41 & _GEN_878;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2037 = _GEN_41 & _GEN_880;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2038 = _GEN_41 & _GEN_882;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2039 = _GEN_41 & _GEN_884;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2040 = _GEN_41 & _GEN_886;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2041 = _GEN_41 & _GEN_888;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2042 = _GEN_41 & _GEN_890;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2043 = _GEN_41 & _GEN_892;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2044 = _GEN_41 & _GEN_894;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2045 = _GEN_41 & _GEN_896;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2046 = _GEN_41 & _GEN_898;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2047 = _GEN_41 & _GEN_900;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2048 = _GEN_41 & _GEN_902;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2049 = _GEN_41 & _GEN_904;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2050 =
      _GEN_41 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_2051 = _GEN_907 | _GEN_2019;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2052;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2053 = _GEN_910 | _GEN_2020;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2054;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2055 = _GEN_913 | _GEN_2021;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2056;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2057 = _GEN_916 | _GEN_2022;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2058;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2059 = _GEN_919 | _GEN_2023;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2060;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2061 = _GEN_922 | _GEN_2024;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2062;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2063 = _GEN_925 | _GEN_2025;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2064;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2065 = _GEN_928 | _GEN_2026;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2066;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2067 = _GEN_931 | _GEN_2027;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2068;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2069 = _GEN_934 | _GEN_2028;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2070;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2071 = _GEN_937 | _GEN_2029;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2072;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2073 = _GEN_940 | _GEN_2030;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2074;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2075 = _GEN_943 | _GEN_2031;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2076;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2077 = _GEN_946 | _GEN_2032;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2078;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2079 = _GEN_949 | _GEN_2033;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2080;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2081 = _GEN_952 | _GEN_2034;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2082;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2083 = _GEN_955 | _GEN_2035;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2084;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2085 = _GEN_958 | _GEN_2036;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2086;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2087 = _GEN_961 | _GEN_2037;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2088;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2089 = _GEN_964 | _GEN_2038;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2090;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2091 = _GEN_967 | _GEN_2039;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2092;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2093 = _GEN_970 | _GEN_2040;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2094;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2095 = _GEN_973 | _GEN_2041;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2096;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2097 = _GEN_976 | _GEN_2042;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2098;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2099 = _GEN_979 | _GEN_2043;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2100;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2101 = _GEN_982 | _GEN_2044;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2102;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2103 = _GEN_985 | _GEN_2045;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2104;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2105 = _GEN_988 | _GEN_2046;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2106;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2107 = _GEN_991 | _GEN_2047;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2108;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2109 = _GEN_994 | _GEN_2048;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2110;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2111 = _GEN_997 | _GEN_2049;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2112;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2113 =
      (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_2050;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_2114;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2115;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2116;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2117;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2118;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2119;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2120;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2121;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2122;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2123;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2124;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2125;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2126;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2127;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2128;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2129;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2130;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2131;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2132;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2133;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2134;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2135;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2136;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2137;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2138;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2139;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2140;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2141;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2142;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2143;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2144;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2145;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2146;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2147 = _GEN_43 & _GEN_1034;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2148 = _GEN_43 & _GEN_1036;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2149 = _GEN_43 & _GEN_1038;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2150 = _GEN_43 & _GEN_1040;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2151 = _GEN_43 & _GEN_1042;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2152 = _GEN_43 & _GEN_1044;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2153 = _GEN_43 & _GEN_1046;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2154 = _GEN_43 & _GEN_1048;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2155 = _GEN_43 & _GEN_1050;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2156 = _GEN_43 & _GEN_1052;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2157 = _GEN_43 & _GEN_1054;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2158 = _GEN_43 & _GEN_1056;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2159 = _GEN_43 & _GEN_1058;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2160 = _GEN_43 & _GEN_1060;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2161 = _GEN_43 & _GEN_1062;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2162 = _GEN_43 & _GEN_1064;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2163 = _GEN_43 & _GEN_1066;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2164 = _GEN_43 & _GEN_1068;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2165 = _GEN_43 & _GEN_1070;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2166 = _GEN_43 & _GEN_1072;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2167 = _GEN_43 & _GEN_1074;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2168 = _GEN_43 & _GEN_1076;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2169 = _GEN_43 & _GEN_1078;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2170 = _GEN_43 & _GEN_1080;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2171 = _GEN_43 & _GEN_1082;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2172 = _GEN_43 & _GEN_1084;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2173 = _GEN_43 & _GEN_1086;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2174 = _GEN_43 & _GEN_1088;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2175 = _GEN_43 & _GEN_1090;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2176 = _GEN_43 & _GEN_1092;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2177 = _GEN_43 & _GEN_1094;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2178 =
      _GEN_43 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_2179 = _GEN_1097 | _GEN_2147;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2180;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2181 = _GEN_1100 | _GEN_2148;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2182;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2183 = _GEN_1103 | _GEN_2149;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2184;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2185 = _GEN_1106 | _GEN_2150;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2186;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2187 = _GEN_1109 | _GEN_2151;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2188;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2189 = _GEN_1112 | _GEN_2152;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2190;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2191 = _GEN_1115 | _GEN_2153;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2192;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2193 = _GEN_1118 | _GEN_2154;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2194;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2195 = _GEN_1121 | _GEN_2155;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2196;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2197 = _GEN_1124 | _GEN_2156;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2198;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2199 = _GEN_1127 | _GEN_2157;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2200;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2201 = _GEN_1130 | _GEN_2158;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2202;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2203 = _GEN_1133 | _GEN_2159;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2204;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2205 = _GEN_1136 | _GEN_2160;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2206;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2207 = _GEN_1139 | _GEN_2161;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2208;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2209 = _GEN_1142 | _GEN_2162;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2210;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2211 = _GEN_1145 | _GEN_2163;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2212;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2213 = _GEN_1148 | _GEN_2164;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2214;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2215 = _GEN_1151 | _GEN_2165;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2216;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2217 = _GEN_1154 | _GEN_2166;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2218;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2219 = _GEN_1157 | _GEN_2167;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2220;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2221 = _GEN_1160 | _GEN_2168;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2222;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2223 = _GEN_1163 | _GEN_2169;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2224;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2225 = _GEN_1166 | _GEN_2170;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2226;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2227 = _GEN_1169 | _GEN_2171;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2228;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2229 = _GEN_1172 | _GEN_2172;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2230;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2231 = _GEN_1175 | _GEN_2173;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2232;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2233 = _GEN_1178 | _GEN_2174;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2234;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2235 = _GEN_1181 | _GEN_2175;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2236;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2237 = _GEN_1184 | _GEN_2176;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2238;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2239 = _GEN_1187 | _GEN_2177;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2240;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2241 =
      (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_2178;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_2242;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2243;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2244;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2245;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2246;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2247;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2248;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2249;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2250;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2251;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2252;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2253;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2254;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2255;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2256;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2257;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2258;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2259;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2260;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2261;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2262;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2263;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2264;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2265;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2266;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2267;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2268;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2269;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2270;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2271;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2272;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2273;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2274;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2275 = _GEN_45 & _GEN_1224;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2276 = _GEN_45 & _GEN_1226;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2277 = _GEN_45 & _GEN_1228;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2278 = _GEN_45 & _GEN_1230;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2279 = _GEN_45 & _GEN_1232;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2280 = _GEN_45 & _GEN_1234;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2281 = _GEN_45 & _GEN_1236;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2282 = _GEN_45 & _GEN_1238;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2283 = _GEN_45 & _GEN_1240;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2284 = _GEN_45 & _GEN_1242;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2285 = _GEN_45 & _GEN_1244;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2286 = _GEN_45 & _GEN_1246;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2287 = _GEN_45 & _GEN_1248;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2288 = _GEN_45 & _GEN_1250;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2289 = _GEN_45 & _GEN_1252;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2290 = _GEN_45 & _GEN_1254;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2291 = _GEN_45 & _GEN_1256;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2292 = _GEN_45 & _GEN_1258;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2293 = _GEN_45 & _GEN_1260;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2294 = _GEN_45 & _GEN_1262;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2295 = _GEN_45 & _GEN_1264;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2296 = _GEN_45 & _GEN_1266;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2297 = _GEN_45 & _GEN_1268;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2298 = _GEN_45 & _GEN_1270;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2299 = _GEN_45 & _GEN_1272;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2300 = _GEN_45 & _GEN_1274;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2301 = _GEN_45 & _GEN_1276;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2302 = _GEN_45 & _GEN_1278;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2303 = _GEN_45 & _GEN_1280;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2304 = _GEN_45 & _GEN_1282;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2305 = _GEN_45 & _GEN_1284;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2306 = _GEN_45 & (&(io_lsu_clr_bsy_0_bits[6:2]));	// rob.scala:236:31, :268:25, :346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_2307 = _GEN_1287 | _GEN_2275;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2308 = _GEN_1289 | _GEN_2276;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2309 = _GEN_1291 | _GEN_2277;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2310 = _GEN_1293 | _GEN_2278;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2311 = _GEN_1295 | _GEN_2279;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2312 = _GEN_1297 | _GEN_2280;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2313 = _GEN_1299 | _GEN_2281;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2314 = _GEN_1301 | _GEN_2282;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2315 = _GEN_1303 | _GEN_2283;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2316 = _GEN_1305 | _GEN_2284;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2317 = _GEN_1307 | _GEN_2285;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2318 = _GEN_1309 | _GEN_2286;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2319 = _GEN_1311 | _GEN_2287;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2320 = _GEN_1313 | _GEN_2288;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2321 = _GEN_1315 | _GEN_2289;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2322 = _GEN_1317 | _GEN_2290;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2323 = _GEN_1319 | _GEN_2291;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2324 = _GEN_1321 | _GEN_2292;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2325 = _GEN_1323 | _GEN_2293;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2326 = _GEN_1325 | _GEN_2294;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2327 = _GEN_1327 | _GEN_2295;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2328 = _GEN_1329 | _GEN_2296;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2329 = _GEN_1331 | _GEN_2297;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2330 = _GEN_1333 | _GEN_2298;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2331 = _GEN_1335 | _GEN_2299;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2332 = _GEN_1337 | _GEN_2300;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2333 = _GEN_1339 | _GEN_2301;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2334 = _GEN_1341 | _GEN_2302;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2335 = _GEN_1343 | _GEN_2303;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2336 = _GEN_1345 | _GEN_2304;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2337 = _GEN_1347 | _GEN_2305;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2338 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_2306;	// rob.scala:236:31, :268:25, :346:69, :361:75, :363:26
    automatic logic             _GEN_2339 = _GEN_48 & _GEN_1350;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2340 = _GEN_48 & _GEN_1352;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2341 = _GEN_48 & _GEN_1354;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2342 = _GEN_48 & _GEN_1356;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2343 = _GEN_48 & _GEN_1358;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2344 = _GEN_48 & _GEN_1360;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2345 = _GEN_48 & _GEN_1362;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2346 = _GEN_48 & _GEN_1364;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2347 = _GEN_48 & _GEN_1366;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2348 = _GEN_48 & _GEN_1368;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2349 = _GEN_48 & _GEN_1370;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2350 = _GEN_48 & _GEN_1372;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2351 = _GEN_48 & _GEN_1374;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2352 = _GEN_48 & _GEN_1376;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2353 = _GEN_48 & _GEN_1378;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2354 = _GEN_48 & _GEN_1380;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2355 = _GEN_48 & _GEN_1382;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2356 = _GEN_48 & _GEN_1384;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2357 = _GEN_48 & _GEN_1386;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2358 = _GEN_48 & _GEN_1388;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2359 = _GEN_48 & _GEN_1390;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2360 = _GEN_48 & _GEN_1392;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2361 = _GEN_48 & _GEN_1394;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2362 = _GEN_48 & _GEN_1396;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2363 = _GEN_48 & _GEN_1398;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2364 = _GEN_48 & _GEN_1400;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2365 = _GEN_48 & _GEN_1402;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2366 = _GEN_48 & _GEN_1404;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2367 = _GEN_48 & _GEN_1406;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2368 = _GEN_48 & _GEN_1408;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2369 = _GEN_48 & _GEN_1410;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_2370 = _GEN_48 & (&(io_lsu_clr_bsy_2_bits[6:2]));	// rob.scala:236:31, :268:25, :361:{31,75}, :363:26
    automatic logic             _GEN_2371;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2372;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2373;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2374;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2375;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2376;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2377;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2378;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2379;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2380;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2381;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2382;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2383;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2384;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2385;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2386;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2387;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2388;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2389;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2390;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2391;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2392;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2393;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2394;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2395;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2396;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2397;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2398;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2399;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2400;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2401;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2402;	// rob.scala:323:29, :433:20, :434:30
    automatic logic [19:0]      _GEN_2403;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2404;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2405;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2406;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2407;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2408;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2409;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2410;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2411;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2412;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2413;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2414;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2415;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2416;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2417;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2418;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2419;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2420;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2421;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2422;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2423;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2424;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2425;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2426;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2427;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2428;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2429;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2430;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2431;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2432;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2433;	// util.scala:118:51
    automatic logic [19:0]      _GEN_2434;	// util.scala:118:51
    automatic logic             _GEN_2435;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2436;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2437;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2438;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2439;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2440;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2441;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2442;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2443;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2444;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2445;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2446;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2447;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2448;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2449;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2450;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2451;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2452;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2453;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2454;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2455;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2456;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2457;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2458;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2459;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2460;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2461;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2462;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2463;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2464;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2465;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_2466;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _rob_bsy_T_4 =
      io_enq_uops_2_is_fence | io_enq_uops_2_is_fencei;	// rob.scala:325:60
    automatic logic             _GEN_2467;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2468;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2469;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2470;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2471;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2472;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2473;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2474;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2475;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2476;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2477;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2478;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2479;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2480;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2481;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2482;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2483;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2484;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2485;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2486;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2487;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2488;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2489;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2490;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2491;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2492;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2493;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2494;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2495;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2496;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2497;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_2498;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _rob_unsafe_T_14 =
      io_enq_uops_2_uses_ldq | io_enq_uops_2_uses_stq & ~io_enq_uops_2_is_fence
      | io_enq_uops_2_is_br | io_enq_uops_2_is_jalr;	// micro-op.scala:152:{48,51,71}
    automatic logic             _GEN_2499;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2500;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2501;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2502;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2503;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2504;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2505;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2506;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2507;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2508;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2509;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2510;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2511;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2512;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2513;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2514;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2515;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2516;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2517;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2518;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2519;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2520;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2521;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2522;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2523;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2524;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2525;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2526;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2527;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2528;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2529;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2530;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_2531 = _GEN_70 & _GEN_274;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2532 = _GEN_70 & _GEN_276;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2533 = _GEN_70 & _GEN_278;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2534 = _GEN_70 & _GEN_280;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2535 = _GEN_70 & _GEN_282;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2536 = _GEN_70 & _GEN_284;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2537 = _GEN_70 & _GEN_286;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2538 = _GEN_70 & _GEN_288;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2539 = _GEN_70 & _GEN_290;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2540 = _GEN_70 & _GEN_292;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2541 = _GEN_70 & _GEN_294;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2542 = _GEN_70 & _GEN_296;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2543 = _GEN_70 & _GEN_298;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2544 = _GEN_70 & _GEN_300;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2545 = _GEN_70 & _GEN_302;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2546 = _GEN_70 & _GEN_304;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2547 = _GEN_70 & _GEN_306;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2548 = _GEN_70 & _GEN_308;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2549 = _GEN_70 & _GEN_310;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2550 = _GEN_70 & _GEN_312;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2551 = _GEN_70 & _GEN_314;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2552 = _GEN_70 & _GEN_316;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2553 = _GEN_70 & _GEN_318;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2554 = _GEN_70 & _GEN_320;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2555 = _GEN_70 & _GEN_322;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2556 = _GEN_70 & _GEN_324;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2557 = _GEN_70 & _GEN_326;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2558 = _GEN_70 & _GEN_328;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2559 = _GEN_70 & _GEN_330;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2560 = _GEN_70 & _GEN_332;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2561 = _GEN_70 & _GEN_334;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2562 =
      _GEN_70 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_2563 = _GEN_337 | _GEN_2531;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2564;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2565 = _GEN_340 | _GEN_2532;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2566;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2567 = _GEN_343 | _GEN_2533;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2568;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2569 = _GEN_346 | _GEN_2534;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2570;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2571 = _GEN_349 | _GEN_2535;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2572;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2573 = _GEN_352 | _GEN_2536;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2574;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2575 = _GEN_355 | _GEN_2537;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2576;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2577 = _GEN_358 | _GEN_2538;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2578;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2579 = _GEN_361 | _GEN_2539;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2580;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2581 = _GEN_364 | _GEN_2540;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2582;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2583 = _GEN_367 | _GEN_2541;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2584;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2585 = _GEN_370 | _GEN_2542;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2586;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2587 = _GEN_373 | _GEN_2543;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2588;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2589 = _GEN_376 | _GEN_2544;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2590;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2591 = _GEN_379 | _GEN_2545;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2592;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2593 = _GEN_382 | _GEN_2546;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2594;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2595 = _GEN_385 | _GEN_2547;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2596;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2597 = _GEN_388 | _GEN_2548;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2598;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2599 = _GEN_391 | _GEN_2549;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2600;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2601 = _GEN_394 | _GEN_2550;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2602;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2603 = _GEN_397 | _GEN_2551;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2604;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2605 = _GEN_400 | _GEN_2552;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2606;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2607 = _GEN_403 | _GEN_2553;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2608;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2609 = _GEN_406 | _GEN_2554;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2610;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2611 = _GEN_409 | _GEN_2555;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2612;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2613 = _GEN_412 | _GEN_2556;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2614;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2615 = _GEN_415 | _GEN_2557;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2616;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2617 = _GEN_418 | _GEN_2558;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2618;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2619 = _GEN_421 | _GEN_2559;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2620;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2621 = _GEN_424 | _GEN_2560;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2622;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2623 = _GEN_427 | _GEN_2561;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_2624;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2625 =
      (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_2562;	// rob.scala:236:31, :268:25, :323:29, :346:69, :347:31
    automatic logic             _GEN_2626;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2627;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2628;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2629;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2630;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2631;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2632;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2633;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2634;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2635;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2636;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2637;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2638;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2639;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2640;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2641;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2642;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2643;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2644;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2645;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2646;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2647;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2648;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2649;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2650;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2651;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2652;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2653;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2654;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2655;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2656;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2657;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2658;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2659 = _GEN_72 & _GEN_464;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2660 = _GEN_72 & _GEN_466;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2661 = _GEN_72 & _GEN_468;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2662 = _GEN_72 & _GEN_470;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2663 = _GEN_72 & _GEN_472;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2664 = _GEN_72 & _GEN_474;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2665 = _GEN_72 & _GEN_476;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2666 = _GEN_72 & _GEN_478;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2667 = _GEN_72 & _GEN_480;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2668 = _GEN_72 & _GEN_482;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2669 = _GEN_72 & _GEN_484;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2670 = _GEN_72 & _GEN_486;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2671 = _GEN_72 & _GEN_488;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2672 = _GEN_72 & _GEN_490;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2673 = _GEN_72 & _GEN_492;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2674 = _GEN_72 & _GEN_494;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2675 = _GEN_72 & _GEN_496;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2676 = _GEN_72 & _GEN_498;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2677 = _GEN_72 & _GEN_500;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2678 = _GEN_72 & _GEN_502;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2679 = _GEN_72 & _GEN_504;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2680 = _GEN_72 & _GEN_506;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2681 = _GEN_72 & _GEN_508;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2682 = _GEN_72 & _GEN_510;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2683 = _GEN_72 & _GEN_512;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2684 = _GEN_72 & _GEN_514;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2685 = _GEN_72 & _GEN_516;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2686 = _GEN_72 & _GEN_518;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2687 = _GEN_72 & _GEN_520;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2688 = _GEN_72 & _GEN_522;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2689 = _GEN_72 & _GEN_524;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2690 =
      _GEN_72 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_2691 = _GEN_527 | _GEN_2659;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2692;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2693 = _GEN_530 | _GEN_2660;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2694;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2695 = _GEN_533 | _GEN_2661;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2696;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2697 = _GEN_536 | _GEN_2662;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2698;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2699 = _GEN_539 | _GEN_2663;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2700;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2701 = _GEN_542 | _GEN_2664;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2702;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2703 = _GEN_545 | _GEN_2665;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2704;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2705 = _GEN_548 | _GEN_2666;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2706;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2707 = _GEN_551 | _GEN_2667;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2708;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2709 = _GEN_554 | _GEN_2668;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2710;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2711 = _GEN_557 | _GEN_2669;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2712;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2713 = _GEN_560 | _GEN_2670;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2714;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2715 = _GEN_563 | _GEN_2671;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2716;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2717 = _GEN_566 | _GEN_2672;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2718;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2719 = _GEN_569 | _GEN_2673;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2720;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2721 = _GEN_572 | _GEN_2674;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2722;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2723 = _GEN_575 | _GEN_2675;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2724;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2725 = _GEN_578 | _GEN_2676;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2726;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2727 = _GEN_581 | _GEN_2677;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2728;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2729 = _GEN_584 | _GEN_2678;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2730;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2731 = _GEN_587 | _GEN_2679;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2732;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2733 = _GEN_590 | _GEN_2680;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2734;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2735 = _GEN_593 | _GEN_2681;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2736;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2737 = _GEN_596 | _GEN_2682;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2738;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2739 = _GEN_599 | _GEN_2683;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2740;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2741 = _GEN_602 | _GEN_2684;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2742;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2743 = _GEN_605 | _GEN_2685;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2744;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2745 = _GEN_608 | _GEN_2686;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2746;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2747 = _GEN_611 | _GEN_2687;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2748;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2749 = _GEN_614 | _GEN_2688;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2750;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2751 = _GEN_617 | _GEN_2689;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2752;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2753 =
      (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_2690;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_2754;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2755;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2756;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2757;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2758;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2759;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2760;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2761;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2762;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2763;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2764;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2765;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2766;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2767;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2768;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2769;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2770;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2771;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2772;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2773;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2774;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2775;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2776;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2777;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2778;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2779;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2780;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2781;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2782;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2783;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2784;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2785;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2786;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2787 = _GEN_74 & _GEN_654;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2788 = _GEN_74 & _GEN_656;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2789 = _GEN_74 & _GEN_658;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2790 = _GEN_74 & _GEN_660;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2791 = _GEN_74 & _GEN_662;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2792 = _GEN_74 & _GEN_664;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2793 = _GEN_74 & _GEN_666;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2794 = _GEN_74 & _GEN_668;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2795 = _GEN_74 & _GEN_670;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2796 = _GEN_74 & _GEN_672;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2797 = _GEN_74 & _GEN_674;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2798 = _GEN_74 & _GEN_676;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2799 = _GEN_74 & _GEN_678;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2800 = _GEN_74 & _GEN_680;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2801 = _GEN_74 & _GEN_682;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2802 = _GEN_74 & _GEN_684;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2803 = _GEN_74 & _GEN_686;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2804 = _GEN_74 & _GEN_688;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2805 = _GEN_74 & _GEN_690;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2806 = _GEN_74 & _GEN_692;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2807 = _GEN_74 & _GEN_694;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2808 = _GEN_74 & _GEN_696;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2809 = _GEN_74 & _GEN_698;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2810 = _GEN_74 & _GEN_700;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2811 = _GEN_74 & _GEN_702;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2812 = _GEN_74 & _GEN_704;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2813 = _GEN_74 & _GEN_706;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2814 = _GEN_74 & _GEN_708;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2815 = _GEN_74 & _GEN_710;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2816 = _GEN_74 & _GEN_712;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2817 = _GEN_74 & _GEN_714;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2818 =
      _GEN_74 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_2819 = _GEN_717 | _GEN_2787;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2820;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2821 = _GEN_720 | _GEN_2788;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2822;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2823 = _GEN_723 | _GEN_2789;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2824;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2825 = _GEN_726 | _GEN_2790;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2826;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2827 = _GEN_729 | _GEN_2791;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2828;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2829 = _GEN_732 | _GEN_2792;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2830;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2831 = _GEN_735 | _GEN_2793;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2832;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2833 = _GEN_738 | _GEN_2794;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2834;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2835 = _GEN_741 | _GEN_2795;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2836;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2837 = _GEN_744 | _GEN_2796;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2838;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2839 = _GEN_747 | _GEN_2797;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2840;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2841 = _GEN_750 | _GEN_2798;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2842;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2843 = _GEN_753 | _GEN_2799;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2844;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2845 = _GEN_756 | _GEN_2800;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2846;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2847 = _GEN_759 | _GEN_2801;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2848;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2849 = _GEN_762 | _GEN_2802;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2850;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2851 = _GEN_765 | _GEN_2803;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2852;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2853 = _GEN_768 | _GEN_2804;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2854;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2855 = _GEN_771 | _GEN_2805;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2856;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2857 = _GEN_774 | _GEN_2806;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2858;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2859 = _GEN_777 | _GEN_2807;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2860;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2861 = _GEN_780 | _GEN_2808;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2862;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2863 = _GEN_783 | _GEN_2809;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2864;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2865 = _GEN_786 | _GEN_2810;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2866;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2867 = _GEN_789 | _GEN_2811;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2868;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2869 = _GEN_792 | _GEN_2812;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2870;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2871 = _GEN_795 | _GEN_2813;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2872;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2873 = _GEN_798 | _GEN_2814;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2874;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2875 = _GEN_801 | _GEN_2815;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2876;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2877 = _GEN_804 | _GEN_2816;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2878;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2879 = _GEN_807 | _GEN_2817;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2880;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2881 =
      (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2818;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_2882;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2883;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2884;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2885;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2886;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2887;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2888;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2889;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2890;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2891;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2892;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2893;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2894;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2895;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2896;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2897;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2898;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2899;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2900;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2901;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2902;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2903;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2904;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2905;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2906;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2907;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2908;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2909;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2910;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2911;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2912;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2913;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2914;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2915 = _GEN_76 & _GEN_844;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2916 = _GEN_76 & _GEN_846;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2917 = _GEN_76 & _GEN_848;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2918 = _GEN_76 & _GEN_850;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2919 = _GEN_76 & _GEN_852;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2920 = _GEN_76 & _GEN_854;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2921 = _GEN_76 & _GEN_856;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2922 = _GEN_76 & _GEN_858;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2923 = _GEN_76 & _GEN_860;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2924 = _GEN_76 & _GEN_862;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2925 = _GEN_76 & _GEN_864;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2926 = _GEN_76 & _GEN_866;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2927 = _GEN_76 & _GEN_868;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2928 = _GEN_76 & _GEN_870;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2929 = _GEN_76 & _GEN_872;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2930 = _GEN_76 & _GEN_874;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2931 = _GEN_76 & _GEN_876;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2932 = _GEN_76 & _GEN_878;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2933 = _GEN_76 & _GEN_880;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2934 = _GEN_76 & _GEN_882;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2935 = _GEN_76 & _GEN_884;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2936 = _GEN_76 & _GEN_886;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2937 = _GEN_76 & _GEN_888;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2938 = _GEN_76 & _GEN_890;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2939 = _GEN_76 & _GEN_892;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2940 = _GEN_76 & _GEN_894;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2941 = _GEN_76 & _GEN_896;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2942 = _GEN_76 & _GEN_898;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2943 = _GEN_76 & _GEN_900;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2944 = _GEN_76 & _GEN_902;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2945 = _GEN_76 & _GEN_904;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_2946 =
      _GEN_76 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_2947 = _GEN_907 | _GEN_2915;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2948;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2949 = _GEN_910 | _GEN_2916;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2950;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2951 = _GEN_913 | _GEN_2917;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2952;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2953 = _GEN_916 | _GEN_2918;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2954;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2955 = _GEN_919 | _GEN_2919;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2956;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2957 = _GEN_922 | _GEN_2920;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2958;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2959 = _GEN_925 | _GEN_2921;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2960;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2961 = _GEN_928 | _GEN_2922;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2962;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2963 = _GEN_931 | _GEN_2923;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2964;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2965 = _GEN_934 | _GEN_2924;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2966;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2967 = _GEN_937 | _GEN_2925;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2968;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2969 = _GEN_940 | _GEN_2926;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2970;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2971 = _GEN_943 | _GEN_2927;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2972;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2973 = _GEN_946 | _GEN_2928;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2974;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2975 = _GEN_949 | _GEN_2929;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2976;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2977 = _GEN_952 | _GEN_2930;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2978;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2979 = _GEN_955 | _GEN_2931;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2980;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2981 = _GEN_958 | _GEN_2932;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2982;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2983 = _GEN_961 | _GEN_2933;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2984;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2985 = _GEN_964 | _GEN_2934;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2986;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2987 = _GEN_967 | _GEN_2935;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2988;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2989 = _GEN_970 | _GEN_2936;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2990;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2991 = _GEN_973 | _GEN_2937;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2992;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2993 = _GEN_976 | _GEN_2938;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2994;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2995 = _GEN_979 | _GEN_2939;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2996;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2997 = _GEN_982 | _GEN_2940;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2998;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2999 = _GEN_985 | _GEN_2941;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3000;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3001 = _GEN_988 | _GEN_2942;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3002;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3003 = _GEN_991 | _GEN_2943;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3004;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3005 = _GEN_994 | _GEN_2944;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3006;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3007 = _GEN_997 | _GEN_2945;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3008;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3009 =
      (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_2946;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_3010;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3011;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3012;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3013;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3014;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3015;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3016;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3017;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3018;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3019;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3020;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3021;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3022;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3023;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3024;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3025;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3026;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3027;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3028;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3029;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3030;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3031;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3032;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3033;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3034;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3035;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3036;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3037;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3038;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3039;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3040;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3041;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3042;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3043 = _GEN_78 & _GEN_1034;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3044 = _GEN_78 & _GEN_1036;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3045 = _GEN_78 & _GEN_1038;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3046 = _GEN_78 & _GEN_1040;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3047 = _GEN_78 & _GEN_1042;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3048 = _GEN_78 & _GEN_1044;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3049 = _GEN_78 & _GEN_1046;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3050 = _GEN_78 & _GEN_1048;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3051 = _GEN_78 & _GEN_1050;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3052 = _GEN_78 & _GEN_1052;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3053 = _GEN_78 & _GEN_1054;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3054 = _GEN_78 & _GEN_1056;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3055 = _GEN_78 & _GEN_1058;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3056 = _GEN_78 & _GEN_1060;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3057 = _GEN_78 & _GEN_1062;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3058 = _GEN_78 & _GEN_1064;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3059 = _GEN_78 & _GEN_1066;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3060 = _GEN_78 & _GEN_1068;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3061 = _GEN_78 & _GEN_1070;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3062 = _GEN_78 & _GEN_1072;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3063 = _GEN_78 & _GEN_1074;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3064 = _GEN_78 & _GEN_1076;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3065 = _GEN_78 & _GEN_1078;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3066 = _GEN_78 & _GEN_1080;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3067 = _GEN_78 & _GEN_1082;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3068 = _GEN_78 & _GEN_1084;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3069 = _GEN_78 & _GEN_1086;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3070 = _GEN_78 & _GEN_1088;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3071 = _GEN_78 & _GEN_1090;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3072 = _GEN_78 & _GEN_1092;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3073 = _GEN_78 & _GEN_1094;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3074 =
      _GEN_78 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_3075 = _GEN_1097 | _GEN_3043;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3076;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3077 = _GEN_1100 | _GEN_3044;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3078;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3079 = _GEN_1103 | _GEN_3045;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3080;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3081 = _GEN_1106 | _GEN_3046;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3082;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3083 = _GEN_1109 | _GEN_3047;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3084;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3085 = _GEN_1112 | _GEN_3048;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3086;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3087 = _GEN_1115 | _GEN_3049;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3088;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3089 = _GEN_1118 | _GEN_3050;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3090;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3091 = _GEN_1121 | _GEN_3051;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3092;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3093 = _GEN_1124 | _GEN_3052;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3094;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3095 = _GEN_1127 | _GEN_3053;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3096;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3097 = _GEN_1130 | _GEN_3054;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3098;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3099 = _GEN_1133 | _GEN_3055;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3100;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3101 = _GEN_1136 | _GEN_3056;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3102;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3103 = _GEN_1139 | _GEN_3057;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3104;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3105 = _GEN_1142 | _GEN_3058;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3106;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3107 = _GEN_1145 | _GEN_3059;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3108;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3109 = _GEN_1148 | _GEN_3060;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3110;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3111 = _GEN_1151 | _GEN_3061;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3112;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3113 = _GEN_1154 | _GEN_3062;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3114;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3115 = _GEN_1157 | _GEN_3063;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3116;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3117 = _GEN_1160 | _GEN_3064;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3118;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3119 = _GEN_1163 | _GEN_3065;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3120;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3121 = _GEN_1166 | _GEN_3066;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3122;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3123 = _GEN_1169 | _GEN_3067;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3124;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3125 = _GEN_1172 | _GEN_3068;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3126;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3127 = _GEN_1175 | _GEN_3069;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3128;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3129 = _GEN_1178 | _GEN_3070;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3130;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3131 = _GEN_1181 | _GEN_3071;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3132;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3133 = _GEN_1184 | _GEN_3072;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3134;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3135 = _GEN_1187 | _GEN_3073;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3136;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3137 =
      (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_3074;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_3138;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3139;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3140;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3141;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3142;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3143;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3144;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3145;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3146;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3147;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3148;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3149;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3150;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3151;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3152;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3153;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3154;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3155;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3156;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3157;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3158;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3159;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3160;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3161;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3162;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3163;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3164;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3165;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3166;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3167;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3168;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3169;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3170;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3171 = _GEN_80 & _GEN_1224;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3172 = _GEN_80 & _GEN_1226;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3173 = _GEN_80 & _GEN_1228;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3174 = _GEN_80 & _GEN_1230;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3175 = _GEN_80 & _GEN_1232;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3176 = _GEN_80 & _GEN_1234;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3177 = _GEN_80 & _GEN_1236;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3178 = _GEN_80 & _GEN_1238;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3179 = _GEN_80 & _GEN_1240;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3180 = _GEN_80 & _GEN_1242;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3181 = _GEN_80 & _GEN_1244;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3182 = _GEN_80 & _GEN_1246;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3183 = _GEN_80 & _GEN_1248;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3184 = _GEN_80 & _GEN_1250;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3185 = _GEN_80 & _GEN_1252;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3186 = _GEN_80 & _GEN_1254;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3187 = _GEN_80 & _GEN_1256;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3188 = _GEN_80 & _GEN_1258;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3189 = _GEN_80 & _GEN_1260;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3190 = _GEN_80 & _GEN_1262;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3191 = _GEN_80 & _GEN_1264;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3192 = _GEN_80 & _GEN_1266;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3193 = _GEN_80 & _GEN_1268;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3194 = _GEN_80 & _GEN_1270;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3195 = _GEN_80 & _GEN_1272;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3196 = _GEN_80 & _GEN_1274;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3197 = _GEN_80 & _GEN_1276;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3198 = _GEN_80 & _GEN_1278;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3199 = _GEN_80 & _GEN_1280;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3200 = _GEN_80 & _GEN_1282;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3201 = _GEN_80 & _GEN_1284;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3202 = _GEN_80 & (&(io_lsu_clr_bsy_0_bits[6:2]));	// rob.scala:236:31, :268:25, :346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_3203 = _GEN_1287 | _GEN_3171;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3204 = _GEN_1289 | _GEN_3172;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3205 = _GEN_1291 | _GEN_3173;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3206 = _GEN_1293 | _GEN_3174;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3207 = _GEN_1295 | _GEN_3175;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3208 = _GEN_1297 | _GEN_3176;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3209 = _GEN_1299 | _GEN_3177;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3210 = _GEN_1301 | _GEN_3178;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3211 = _GEN_1303 | _GEN_3179;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3212 = _GEN_1305 | _GEN_3180;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3213 = _GEN_1307 | _GEN_3181;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3214 = _GEN_1309 | _GEN_3182;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3215 = _GEN_1311 | _GEN_3183;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3216 = _GEN_1313 | _GEN_3184;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3217 = _GEN_1315 | _GEN_3185;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3218 = _GEN_1317 | _GEN_3186;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3219 = _GEN_1319 | _GEN_3187;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3220 = _GEN_1321 | _GEN_3188;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3221 = _GEN_1323 | _GEN_3189;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3222 = _GEN_1325 | _GEN_3190;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3223 = _GEN_1327 | _GEN_3191;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3224 = _GEN_1329 | _GEN_3192;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3225 = _GEN_1331 | _GEN_3193;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3226 = _GEN_1333 | _GEN_3194;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3227 = _GEN_1335 | _GEN_3195;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3228 = _GEN_1337 | _GEN_3196;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3229 = _GEN_1339 | _GEN_3197;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3230 = _GEN_1341 | _GEN_3198;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3231 = _GEN_1343 | _GEN_3199;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3232 = _GEN_1345 | _GEN_3200;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3233 = _GEN_1347 | _GEN_3201;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_3234 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_3202;	// rob.scala:236:31, :268:25, :346:69, :361:75, :363:26
    automatic logic             _GEN_3235 = _GEN_83 & _GEN_1350;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3236 = _GEN_83 & _GEN_1352;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3237 = _GEN_83 & _GEN_1354;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3238 = _GEN_83 & _GEN_1356;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3239 = _GEN_83 & _GEN_1358;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3240 = _GEN_83 & _GEN_1360;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3241 = _GEN_83 & _GEN_1362;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3242 = _GEN_83 & _GEN_1364;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3243 = _GEN_83 & _GEN_1366;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3244 = _GEN_83 & _GEN_1368;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3245 = _GEN_83 & _GEN_1370;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3246 = _GEN_83 & _GEN_1372;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3247 = _GEN_83 & _GEN_1374;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3248 = _GEN_83 & _GEN_1376;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3249 = _GEN_83 & _GEN_1378;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3250 = _GEN_83 & _GEN_1380;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3251 = _GEN_83 & _GEN_1382;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3252 = _GEN_83 & _GEN_1384;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3253 = _GEN_83 & _GEN_1386;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3254 = _GEN_83 & _GEN_1388;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3255 = _GEN_83 & _GEN_1390;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3256 = _GEN_83 & _GEN_1392;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3257 = _GEN_83 & _GEN_1394;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3258 = _GEN_83 & _GEN_1396;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3259 = _GEN_83 & _GEN_1398;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3260 = _GEN_83 & _GEN_1400;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3261 = _GEN_83 & _GEN_1402;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3262 = _GEN_83 & _GEN_1404;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3263 = _GEN_83 & _GEN_1406;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3264 = _GEN_83 & _GEN_1408;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3265 = _GEN_83 & _GEN_1410;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_3266 = _GEN_83 & (&(io_lsu_clr_bsy_2_bits[6:2]));	// rob.scala:236:31, :268:25, :361:{31,75}, :363:26
    automatic logic             _GEN_3267;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3268;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3269;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3270;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3271;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3272;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3273;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3274;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3275;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3276;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3277;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3278;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3279;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3280;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3281;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3282;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3283;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3284;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3285;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3286;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3287;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3288;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3289;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3290;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3291;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3292;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3293;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3294;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3295;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3296;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3297;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_3298;	// rob.scala:323:29, :433:20, :434:30
    automatic logic [19:0]      _GEN_3299;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3300;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3301;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3302;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3303;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3304;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3305;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3306;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3307;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3308;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3309;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3310;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3311;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3312;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3313;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3314;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3315;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3316;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3317;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3318;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3319;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3320;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3321;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3322;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3323;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3324;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3325;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3326;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3327;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3328;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3329;	// util.scala:118:51
    automatic logic [19:0]      _GEN_3330;	// util.scala:118:51
    automatic logic             _GEN_3331;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3332;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3333;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3334;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3335;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3336;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3337;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3338;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3339;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3340;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3341;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3342;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3343;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3344;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3345;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3346;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3347;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3348;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3349;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3350;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3351;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3352;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3353;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3354;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3355;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3356;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3357;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3358;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3359;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3360;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3361;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_3362;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _rob_bsy_T_6 =
      io_enq_uops_3_is_fence | io_enq_uops_3_is_fencei;	// rob.scala:325:60
    automatic logic             _GEN_3363;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3364;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3365;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3366;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3367;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3368;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3369;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3370;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3371;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3372;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3373;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3374;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3375;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3376;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3377;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3378;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3379;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3380;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3381;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3382;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3383;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3384;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3385;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3386;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3387;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3388;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3389;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3390;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3391;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3392;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3393;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_3394;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _rob_unsafe_T_19 =
      io_enq_uops_3_uses_ldq | io_enq_uops_3_uses_stq & ~io_enq_uops_3_is_fence
      | io_enq_uops_3_is_br | io_enq_uops_3_is_jalr;	// micro-op.scala:152:{48,51,71}
    automatic logic             _GEN_3395;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3396;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3397;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3398;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3399;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3400;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3401;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3402;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3403;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3404;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3405;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3406;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3407;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3408;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3409;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3410;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3411;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3412;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3413;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3414;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3415;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3416;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3417;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3418;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3419;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3420;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3421;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3422;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3423;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3424;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3425;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3426;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_3427 = _GEN_105 & _GEN_274;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3428 = _GEN_105 & _GEN_276;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3429 = _GEN_105 & _GEN_278;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3430 = _GEN_105 & _GEN_280;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3431 = _GEN_105 & _GEN_282;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3432 = _GEN_105 & _GEN_284;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3433 = _GEN_105 & _GEN_286;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3434 = _GEN_105 & _GEN_288;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3435 = _GEN_105 & _GEN_290;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3436 = _GEN_105 & _GEN_292;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3437 = _GEN_105 & _GEN_294;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3438 = _GEN_105 & _GEN_296;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3439 = _GEN_105 & _GEN_298;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3440 = _GEN_105 & _GEN_300;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3441 = _GEN_105 & _GEN_302;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3442 = _GEN_105 & _GEN_304;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3443 = _GEN_105 & _GEN_306;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3444 = _GEN_105 & _GEN_308;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3445 = _GEN_105 & _GEN_310;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3446 = _GEN_105 & _GEN_312;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3447 = _GEN_105 & _GEN_314;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3448 = _GEN_105 & _GEN_316;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3449 = _GEN_105 & _GEN_318;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3450 = _GEN_105 & _GEN_320;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3451 = _GEN_105 & _GEN_322;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3452 = _GEN_105 & _GEN_324;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3453 = _GEN_105 & _GEN_326;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3454 = _GEN_105 & _GEN_328;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3455 = _GEN_105 & _GEN_330;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3456 = _GEN_105 & _GEN_332;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3457 = _GEN_105 & _GEN_334;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3458 =
      _GEN_105 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_3459 = _GEN_337 | _GEN_3427;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3460;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3461 = _GEN_340 | _GEN_3428;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3462;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3463 = _GEN_343 | _GEN_3429;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3464;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3465 = _GEN_346 | _GEN_3430;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3466;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3467 = _GEN_349 | _GEN_3431;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3468;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3469 = _GEN_352 | _GEN_3432;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3470;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3471 = _GEN_355 | _GEN_3433;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3472;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3473 = _GEN_358 | _GEN_3434;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3474;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3475 = _GEN_361 | _GEN_3435;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3476;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3477 = _GEN_364 | _GEN_3436;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3478;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3479 = _GEN_367 | _GEN_3437;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3480;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3481 = _GEN_370 | _GEN_3438;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3482;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3483 = _GEN_373 | _GEN_3439;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3484;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3485 = _GEN_376 | _GEN_3440;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3486;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3487 = _GEN_379 | _GEN_3441;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3488;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3489 = _GEN_382 | _GEN_3442;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3490;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3491 = _GEN_385 | _GEN_3443;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3492;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3493 = _GEN_388 | _GEN_3444;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3494;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3495 = _GEN_391 | _GEN_3445;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3496;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3497 = _GEN_394 | _GEN_3446;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3498;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3499 = _GEN_397 | _GEN_3447;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3500;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3501 = _GEN_400 | _GEN_3448;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3502;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3503 = _GEN_403 | _GEN_3449;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3504;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3505 = _GEN_406 | _GEN_3450;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3506;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3507 = _GEN_409 | _GEN_3451;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3508;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3509 = _GEN_412 | _GEN_3452;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3510;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3511 = _GEN_415 | _GEN_3453;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3512;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3513 = _GEN_418 | _GEN_3454;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3514;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3515 = _GEN_421 | _GEN_3455;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3516;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3517 = _GEN_424 | _GEN_3456;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3518;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3519 = _GEN_427 | _GEN_3457;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_3520;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3521 =
      (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_3458;	// rob.scala:236:31, :268:25, :323:29, :346:69, :347:31
    automatic logic             _GEN_3522;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3523;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3524;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3525;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3526;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3527;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3528;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3529;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3530;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3531;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3532;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3533;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3534;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3535;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3536;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3537;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3538;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3539;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3540;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3541;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3542;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3543;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3544;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3545;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3546;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3547;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3548;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3549;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3550;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3551;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3552;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3553;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3554;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3555 = _GEN_107 & _GEN_464;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3556 = _GEN_107 & _GEN_466;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3557 = _GEN_107 & _GEN_468;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3558 = _GEN_107 & _GEN_470;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3559 = _GEN_107 & _GEN_472;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3560 = _GEN_107 & _GEN_474;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3561 = _GEN_107 & _GEN_476;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3562 = _GEN_107 & _GEN_478;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3563 = _GEN_107 & _GEN_480;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3564 = _GEN_107 & _GEN_482;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3565 = _GEN_107 & _GEN_484;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3566 = _GEN_107 & _GEN_486;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3567 = _GEN_107 & _GEN_488;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3568 = _GEN_107 & _GEN_490;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3569 = _GEN_107 & _GEN_492;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3570 = _GEN_107 & _GEN_494;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3571 = _GEN_107 & _GEN_496;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3572 = _GEN_107 & _GEN_498;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3573 = _GEN_107 & _GEN_500;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3574 = _GEN_107 & _GEN_502;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3575 = _GEN_107 & _GEN_504;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3576 = _GEN_107 & _GEN_506;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3577 = _GEN_107 & _GEN_508;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3578 = _GEN_107 & _GEN_510;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3579 = _GEN_107 & _GEN_512;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3580 = _GEN_107 & _GEN_514;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3581 = _GEN_107 & _GEN_516;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3582 = _GEN_107 & _GEN_518;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3583 = _GEN_107 & _GEN_520;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3584 = _GEN_107 & _GEN_522;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3585 = _GEN_107 & _GEN_524;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3586 =
      _GEN_107 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_3587 = _GEN_527 | _GEN_3555;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3588;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3589 = _GEN_530 | _GEN_3556;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3590;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3591 = _GEN_533 | _GEN_3557;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3592;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3593 = _GEN_536 | _GEN_3558;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3594;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3595 = _GEN_539 | _GEN_3559;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3596;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3597 = _GEN_542 | _GEN_3560;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3598;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3599 = _GEN_545 | _GEN_3561;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3600;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3601 = _GEN_548 | _GEN_3562;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3602;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3603 = _GEN_551 | _GEN_3563;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3604;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3605 = _GEN_554 | _GEN_3564;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3606;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3607 = _GEN_557 | _GEN_3565;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3608;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3609 = _GEN_560 | _GEN_3566;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3610;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3611 = _GEN_563 | _GEN_3567;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3612;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3613 = _GEN_566 | _GEN_3568;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3614;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3615 = _GEN_569 | _GEN_3569;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3616;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3617 = _GEN_572 | _GEN_3570;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3618;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3619 = _GEN_575 | _GEN_3571;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3620;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3621 = _GEN_578 | _GEN_3572;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3622;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3623 = _GEN_581 | _GEN_3573;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3624;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3625 = _GEN_584 | _GEN_3574;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3626;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3627 = _GEN_587 | _GEN_3575;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3628;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3629 = _GEN_590 | _GEN_3576;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3630;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3631 = _GEN_593 | _GEN_3577;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3632;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3633 = _GEN_596 | _GEN_3578;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3634;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3635 = _GEN_599 | _GEN_3579;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3636;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3637 = _GEN_602 | _GEN_3580;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3638;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3639 = _GEN_605 | _GEN_3581;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3640;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3641 = _GEN_608 | _GEN_3582;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3642;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3643 = _GEN_611 | _GEN_3583;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3644;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3645 = _GEN_614 | _GEN_3584;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3646;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3647 = _GEN_617 | _GEN_3585;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3648;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3649 =
      (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_3586;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_3650;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3651;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3652;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3653;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3654;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3655;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3656;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3657;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3658;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3659;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3660;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3661;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3662;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3663;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3664;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3665;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3666;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3667;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3668;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3669;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3670;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3671;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3672;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3673;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3674;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3675;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3676;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3677;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3678;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3679;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3680;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3681;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3682;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3683 = _GEN_109 & _GEN_654;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3684 = _GEN_109 & _GEN_656;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3685 = _GEN_109 & _GEN_658;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3686 = _GEN_109 & _GEN_660;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3687 = _GEN_109 & _GEN_662;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3688 = _GEN_109 & _GEN_664;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3689 = _GEN_109 & _GEN_666;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3690 = _GEN_109 & _GEN_668;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3691 = _GEN_109 & _GEN_670;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3692 = _GEN_109 & _GEN_672;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3693 = _GEN_109 & _GEN_674;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3694 = _GEN_109 & _GEN_676;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3695 = _GEN_109 & _GEN_678;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3696 = _GEN_109 & _GEN_680;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3697 = _GEN_109 & _GEN_682;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3698 = _GEN_109 & _GEN_684;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3699 = _GEN_109 & _GEN_686;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3700 = _GEN_109 & _GEN_688;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3701 = _GEN_109 & _GEN_690;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3702 = _GEN_109 & _GEN_692;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3703 = _GEN_109 & _GEN_694;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3704 = _GEN_109 & _GEN_696;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3705 = _GEN_109 & _GEN_698;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3706 = _GEN_109 & _GEN_700;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3707 = _GEN_109 & _GEN_702;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3708 = _GEN_109 & _GEN_704;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3709 = _GEN_109 & _GEN_706;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3710 = _GEN_109 & _GEN_708;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3711 = _GEN_109 & _GEN_710;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3712 = _GEN_109 & _GEN_712;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3713 = _GEN_109 & _GEN_714;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3714 =
      _GEN_109 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_3715 = _GEN_717 | _GEN_3683;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3716;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3717 = _GEN_720 | _GEN_3684;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3718;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3719 = _GEN_723 | _GEN_3685;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3720;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3721 = _GEN_726 | _GEN_3686;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3722;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3723 = _GEN_729 | _GEN_3687;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3724;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3725 = _GEN_732 | _GEN_3688;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3726;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3727 = _GEN_735 | _GEN_3689;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3728;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3729 = _GEN_738 | _GEN_3690;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3730;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3731 = _GEN_741 | _GEN_3691;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3732;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3733 = _GEN_744 | _GEN_3692;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3734;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3735 = _GEN_747 | _GEN_3693;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3736;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3737 = _GEN_750 | _GEN_3694;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3738;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3739 = _GEN_753 | _GEN_3695;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3740;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3741 = _GEN_756 | _GEN_3696;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3742;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3743 = _GEN_759 | _GEN_3697;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3744;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3745 = _GEN_762 | _GEN_3698;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3746;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3747 = _GEN_765 | _GEN_3699;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3748;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3749 = _GEN_768 | _GEN_3700;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3750;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3751 = _GEN_771 | _GEN_3701;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3752;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3753 = _GEN_774 | _GEN_3702;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3754;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3755 = _GEN_777 | _GEN_3703;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3756;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3757 = _GEN_780 | _GEN_3704;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3758;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3759 = _GEN_783 | _GEN_3705;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3760;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3761 = _GEN_786 | _GEN_3706;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3762;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3763 = _GEN_789 | _GEN_3707;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3764;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3765 = _GEN_792 | _GEN_3708;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3766;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3767 = _GEN_795 | _GEN_3709;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3768;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3769 = _GEN_798 | _GEN_3710;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3770;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3771 = _GEN_801 | _GEN_3711;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3772;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3773 = _GEN_804 | _GEN_3712;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3774;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3775 = _GEN_807 | _GEN_3713;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3776;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3777 =
      (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_3714;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_3778;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3779;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3780;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3781;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3782;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3783;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3784;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3785;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3786;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3787;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3788;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3789;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3790;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3791;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3792;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3793;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3794;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3795;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3796;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3797;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3798;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3799;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3800;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3801;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3802;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3803;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3804;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3805;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3806;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3807;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3808;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3809;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3810;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3811 = _GEN_111 & _GEN_844;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3812 = _GEN_111 & _GEN_846;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3813 = _GEN_111 & _GEN_848;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3814 = _GEN_111 & _GEN_850;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3815 = _GEN_111 & _GEN_852;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3816 = _GEN_111 & _GEN_854;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3817 = _GEN_111 & _GEN_856;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3818 = _GEN_111 & _GEN_858;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3819 = _GEN_111 & _GEN_860;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3820 = _GEN_111 & _GEN_862;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3821 = _GEN_111 & _GEN_864;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3822 = _GEN_111 & _GEN_866;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3823 = _GEN_111 & _GEN_868;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3824 = _GEN_111 & _GEN_870;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3825 = _GEN_111 & _GEN_872;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3826 = _GEN_111 & _GEN_874;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3827 = _GEN_111 & _GEN_876;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3828 = _GEN_111 & _GEN_878;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3829 = _GEN_111 & _GEN_880;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3830 = _GEN_111 & _GEN_882;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3831 = _GEN_111 & _GEN_884;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3832 = _GEN_111 & _GEN_886;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3833 = _GEN_111 & _GEN_888;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3834 = _GEN_111 & _GEN_890;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3835 = _GEN_111 & _GEN_892;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3836 = _GEN_111 & _GEN_894;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3837 = _GEN_111 & _GEN_896;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3838 = _GEN_111 & _GEN_898;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3839 = _GEN_111 & _GEN_900;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3840 = _GEN_111 & _GEN_902;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3841 = _GEN_111 & _GEN_904;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3842 =
      _GEN_111 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_3843 = _GEN_907 | _GEN_3811;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3844;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3845 = _GEN_910 | _GEN_3812;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3846;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3847 = _GEN_913 | _GEN_3813;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3848;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3849 = _GEN_916 | _GEN_3814;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3850;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3851 = _GEN_919 | _GEN_3815;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3852;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3853 = _GEN_922 | _GEN_3816;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3854;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3855 = _GEN_925 | _GEN_3817;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3856;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3857 = _GEN_928 | _GEN_3818;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3858;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3859 = _GEN_931 | _GEN_3819;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3860;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3861 = _GEN_934 | _GEN_3820;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3862;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3863 = _GEN_937 | _GEN_3821;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3864;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3865 = _GEN_940 | _GEN_3822;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3866;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3867 = _GEN_943 | _GEN_3823;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3868;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3869 = _GEN_946 | _GEN_3824;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3870;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3871 = _GEN_949 | _GEN_3825;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3872;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3873 = _GEN_952 | _GEN_3826;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3874;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3875 = _GEN_955 | _GEN_3827;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3876;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3877 = _GEN_958 | _GEN_3828;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3878;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3879 = _GEN_961 | _GEN_3829;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3880;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3881 = _GEN_964 | _GEN_3830;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3882;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3883 = _GEN_967 | _GEN_3831;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3884;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3885 = _GEN_970 | _GEN_3832;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3886;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3887 = _GEN_973 | _GEN_3833;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3888;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3889 = _GEN_976 | _GEN_3834;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3890;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3891 = _GEN_979 | _GEN_3835;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3892;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3893 = _GEN_982 | _GEN_3836;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3894;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3895 = _GEN_985 | _GEN_3837;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3896;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3897 = _GEN_988 | _GEN_3838;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3898;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3899 = _GEN_991 | _GEN_3839;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3900;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3901 = _GEN_994 | _GEN_3840;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3902;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3903 = _GEN_997 | _GEN_3841;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3904;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3905 =
      (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_3842;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_3906;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3907;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3908;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3909;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3910;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3911;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3912;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3913;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3914;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3915;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3916;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3917;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3918;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3919;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3920;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3921;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3922;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3923;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3924;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3925;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3926;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3927;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3928;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3929;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3930;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3931;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3932;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3933;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3934;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3935;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3936;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3937;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3938;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_3939 = _GEN_113 & _GEN_1034;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3940 = _GEN_113 & _GEN_1036;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3941 = _GEN_113 & _GEN_1038;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3942 = _GEN_113 & _GEN_1040;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3943 = _GEN_113 & _GEN_1042;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3944 = _GEN_113 & _GEN_1044;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3945 = _GEN_113 & _GEN_1046;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3946 = _GEN_113 & _GEN_1048;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3947 = _GEN_113 & _GEN_1050;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3948 = _GEN_113 & _GEN_1052;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3949 = _GEN_113 & _GEN_1054;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3950 = _GEN_113 & _GEN_1056;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3951 = _GEN_113 & _GEN_1058;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3952 = _GEN_113 & _GEN_1060;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3953 = _GEN_113 & _GEN_1062;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3954 = _GEN_113 & _GEN_1064;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3955 = _GEN_113 & _GEN_1066;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3956 = _GEN_113 & _GEN_1068;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3957 = _GEN_113 & _GEN_1070;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3958 = _GEN_113 & _GEN_1072;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3959 = _GEN_113 & _GEN_1074;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3960 = _GEN_113 & _GEN_1076;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3961 = _GEN_113 & _GEN_1078;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3962 = _GEN_113 & _GEN_1080;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3963 = _GEN_113 & _GEN_1082;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3964 = _GEN_113 & _GEN_1084;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3965 = _GEN_113 & _GEN_1086;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3966 = _GEN_113 & _GEN_1088;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3967 = _GEN_113 & _GEN_1090;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3968 = _GEN_113 & _GEN_1092;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3969 = _GEN_113 & _GEN_1094;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_3970 =
      _GEN_113 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_3971 = _GEN_1097 | _GEN_3939;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3972;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3973 = _GEN_1100 | _GEN_3940;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3974;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3975 = _GEN_1103 | _GEN_3941;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3976;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3977 = _GEN_1106 | _GEN_3942;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3978;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3979 = _GEN_1109 | _GEN_3943;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3980;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3981 = _GEN_1112 | _GEN_3944;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3982;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3983 = _GEN_1115 | _GEN_3945;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3984;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3985 = _GEN_1118 | _GEN_3946;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3986;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3987 = _GEN_1121 | _GEN_3947;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3988;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3989 = _GEN_1124 | _GEN_3948;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3990;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3991 = _GEN_1127 | _GEN_3949;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3992;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3993 = _GEN_1130 | _GEN_3950;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3994;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3995 = _GEN_1133 | _GEN_3951;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3996;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3997 = _GEN_1136 | _GEN_3952;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3998;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_3999 = _GEN_1139 | _GEN_3953;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4000;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4001 = _GEN_1142 | _GEN_3954;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4002;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4003 = _GEN_1145 | _GEN_3955;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4004;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4005 = _GEN_1148 | _GEN_3956;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4006;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4007 = _GEN_1151 | _GEN_3957;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4008;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4009 = _GEN_1154 | _GEN_3958;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4010;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4011 = _GEN_1157 | _GEN_3959;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4012;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4013 = _GEN_1160 | _GEN_3960;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4014;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4015 = _GEN_1163 | _GEN_3961;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4016;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4017 = _GEN_1166 | _GEN_3962;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4018;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4019 = _GEN_1169 | _GEN_3963;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4020;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4021 = _GEN_1172 | _GEN_3964;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4022;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4023 = _GEN_1175 | _GEN_3965;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4024;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4025 = _GEN_1178 | _GEN_3966;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4026;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4027 = _GEN_1181 | _GEN_3967;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4028;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4029 = _GEN_1184 | _GEN_3968;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4030;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4031 = _GEN_1187 | _GEN_3969;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4032;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4033 =
      (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_3970;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_4034;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_4035;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4036;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4037;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4038;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4039;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4040;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4041;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4042;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4043;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4044;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4045;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4046;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4047;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4048;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4049;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4050;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4051;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4052;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4053;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4054;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4055;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4056;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4057;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4058;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4059;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4060;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4061;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4062;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4063;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4064;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4065;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4066;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_4067 = _GEN_115 & _GEN_1224;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4068 = _GEN_115 & _GEN_1226;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4069 = _GEN_115 & _GEN_1228;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4070 = _GEN_115 & _GEN_1230;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4071 = _GEN_115 & _GEN_1232;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4072 = _GEN_115 & _GEN_1234;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4073 = _GEN_115 & _GEN_1236;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4074 = _GEN_115 & _GEN_1238;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4075 = _GEN_115 & _GEN_1240;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4076 = _GEN_115 & _GEN_1242;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4077 = _GEN_115 & _GEN_1244;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4078 = _GEN_115 & _GEN_1246;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4079 = _GEN_115 & _GEN_1248;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4080 = _GEN_115 & _GEN_1250;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4081 = _GEN_115 & _GEN_1252;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4082 = _GEN_115 & _GEN_1254;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4083 = _GEN_115 & _GEN_1256;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4084 = _GEN_115 & _GEN_1258;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4085 = _GEN_115 & _GEN_1260;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4086 = _GEN_115 & _GEN_1262;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4087 = _GEN_115 & _GEN_1264;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4088 = _GEN_115 & _GEN_1266;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4089 = _GEN_115 & _GEN_1268;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4090 = _GEN_115 & _GEN_1270;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4091 = _GEN_115 & _GEN_1272;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4092 = _GEN_115 & _GEN_1274;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4093 = _GEN_115 & _GEN_1276;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4094 = _GEN_115 & _GEN_1278;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4095 = _GEN_115 & _GEN_1280;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4096 = _GEN_115 & _GEN_1282;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4097 = _GEN_115 & _GEN_1284;	// rob.scala:346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4098 = _GEN_115 & (&(io_lsu_clr_bsy_0_bits[6:2]));	// rob.scala:236:31, :268:25, :346:69, :361:{31,75}, :363:26
    automatic logic             _GEN_4099 = _GEN_1287 | _GEN_4067;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4100 = _GEN_1289 | _GEN_4068;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4101 = _GEN_1291 | _GEN_4069;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4102 = _GEN_1293 | _GEN_4070;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4103 = _GEN_1295 | _GEN_4071;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4104 = _GEN_1297 | _GEN_4072;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4105 = _GEN_1299 | _GEN_4073;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4106 = _GEN_1301 | _GEN_4074;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4107 = _GEN_1303 | _GEN_4075;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4108 = _GEN_1305 | _GEN_4076;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4109 = _GEN_1307 | _GEN_4077;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4110 = _GEN_1309 | _GEN_4078;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4111 = _GEN_1311 | _GEN_4079;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4112 = _GEN_1313 | _GEN_4080;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4113 = _GEN_1315 | _GEN_4081;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4114 = _GEN_1317 | _GEN_4082;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4115 = _GEN_1319 | _GEN_4083;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4116 = _GEN_1321 | _GEN_4084;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4117 = _GEN_1323 | _GEN_4085;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4118 = _GEN_1325 | _GEN_4086;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4119 = _GEN_1327 | _GEN_4087;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4120 = _GEN_1329 | _GEN_4088;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4121 = _GEN_1331 | _GEN_4089;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4122 = _GEN_1333 | _GEN_4090;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4123 = _GEN_1335 | _GEN_4091;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4124 = _GEN_1337 | _GEN_4092;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4125 = _GEN_1339 | _GEN_4093;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4126 = _GEN_1341 | _GEN_4094;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4127 = _GEN_1343 | _GEN_4095;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4128 = _GEN_1345 | _GEN_4096;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4129 = _GEN_1347 | _GEN_4097;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_4130 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_4098;	// rob.scala:236:31, :268:25, :346:69, :361:75, :363:26
    automatic logic             _GEN_4131 = _GEN_118 & _GEN_1350;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4132 = _GEN_118 & _GEN_1352;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4133 = _GEN_118 & _GEN_1354;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4134 = _GEN_118 & _GEN_1356;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4135 = _GEN_118 & _GEN_1358;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4136 = _GEN_118 & _GEN_1360;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4137 = _GEN_118 & _GEN_1362;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4138 = _GEN_118 & _GEN_1364;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4139 = _GEN_118 & _GEN_1366;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4140 = _GEN_118 & _GEN_1368;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4141 = _GEN_118 & _GEN_1370;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4142 = _GEN_118 & _GEN_1372;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4143 = _GEN_118 & _GEN_1374;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4144 = _GEN_118 & _GEN_1376;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4145 = _GEN_118 & _GEN_1378;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4146 = _GEN_118 & _GEN_1380;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4147 = _GEN_118 & _GEN_1382;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4148 = _GEN_118 & _GEN_1384;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4149 = _GEN_118 & _GEN_1386;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4150 = _GEN_118 & _GEN_1388;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4151 = _GEN_118 & _GEN_1390;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4152 = _GEN_118 & _GEN_1392;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4153 = _GEN_118 & _GEN_1394;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4154 = _GEN_118 & _GEN_1396;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4155 = _GEN_118 & _GEN_1398;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4156 = _GEN_118 & _GEN_1400;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4157 = _GEN_118 & _GEN_1402;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4158 = _GEN_118 & _GEN_1404;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4159 = _GEN_118 & _GEN_1406;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4160 = _GEN_118 & _GEN_1408;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4161 = _GEN_118 & _GEN_1410;	// rob.scala:361:{31,75}, :363:26
    automatic logic             _GEN_4162 = _GEN_118 & (&(io_lsu_clr_bsy_2_bits[6:2]));	// rob.scala:236:31, :268:25, :361:{31,75}, :363:26
    automatic logic             _GEN_4163;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4164;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4165;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4166;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4167;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4168;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4169;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4170;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4171;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4172;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4173;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4174;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4175;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4176;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4177;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4178;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4179;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4180;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4181;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4182;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4183;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4184;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4185;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4186;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4187;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4188;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4189;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4190;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4191;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4192;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4193;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_4194;	// rob.scala:323:29, :433:20, :434:30
    automatic logic [19:0]      _GEN_4195;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4196;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4197;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4198;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4199;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4200;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4201;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4202;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4203;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4204;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4205;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4206;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4207;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4208;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4209;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4210;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4211;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4212;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4213;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4214;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4215;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4216;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4217;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4218;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4219;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4220;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4221;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4222;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4223;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4224;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4225;	// util.scala:118:51
    automatic logic [19:0]      _GEN_4226;	// util.scala:118:51
    automatic logic             enq_xcpts_0 = io_enq_valids_0 & io_enq_uops_0_exception;	// rob.scala:628:38
    automatic logic             enq_xcpts_1 = io_enq_valids_1 & io_enq_uops_1_exception;	// rob.scala:628:38
    automatic logic             enq_xcpts_2 = io_enq_valids_2 & io_enq_uops_2_exception;	// rob.scala:628:38
    automatic logic             _GEN_4227;	// rob.scala:631:47
    automatic logic             _GEN_4228;	// rob.scala:635:25
    automatic logic             _GEN_4229;	// rob.scala:641:30
    automatic logic [1:0]       idx;	// rob.scala:642:37
    automatic logic [3:0][19:0] _GEN_4230 =
      {{io_enq_uops_3_br_mask},
       {io_enq_uops_2_br_mask},
       {io_enq_uops_1_br_mask},
       {io_enq_uops_0_br_mask}};	// rob.scala:646:23
    automatic logic [19:0]      next_xcpt_uop_br_mask;	// rob.scala:625:17, :631:76, :632:27
    automatic logic [3:0]       _GEN_4231;	// rob.scala:865:98
    _GEN_147 = rob_tail == 5'h0;	// rob.scala:228:29, :236:31, :268:25, :324:31
    _GEN_148 = io_enq_valids_0 & _GEN_147;	// rob.scala:307:32, :323:29, :324:31
    _GEN_149 = rob_tail == 5'h1;	// rob.scala:228:29, :324:31
    _GEN_150 = io_enq_valids_0 & _GEN_149;	// rob.scala:307:32, :323:29, :324:31
    _GEN_151 = rob_tail == 5'h2;	// rob.scala:228:29, :324:31
    _GEN_152 = io_enq_valids_0 & _GEN_151;	// rob.scala:307:32, :323:29, :324:31
    _GEN_153 = rob_tail == 5'h3;	// rob.scala:228:29, :324:31
    _GEN_154 = io_enq_valids_0 & _GEN_153;	// rob.scala:307:32, :323:29, :324:31
    _GEN_155 = rob_tail == 5'h4;	// rob.scala:228:29, :324:31
    _GEN_156 = io_enq_valids_0 & _GEN_155;	// rob.scala:307:32, :323:29, :324:31
    _GEN_157 = rob_tail == 5'h5;	// rob.scala:228:29, :324:31
    _GEN_158 = io_enq_valids_0 & _GEN_157;	// rob.scala:307:32, :323:29, :324:31
    _GEN_159 = rob_tail == 5'h6;	// rob.scala:228:29, :324:31
    _GEN_160 = io_enq_valids_0 & _GEN_159;	// rob.scala:307:32, :323:29, :324:31
    _GEN_161 = rob_tail == 5'h7;	// rob.scala:228:29, :324:31
    _GEN_162 = io_enq_valids_0 & _GEN_161;	// rob.scala:307:32, :323:29, :324:31
    _GEN_163 = rob_tail == 5'h8;	// rob.scala:228:29, :324:31
    _GEN_164 = io_enq_valids_0 & _GEN_163;	// rob.scala:307:32, :323:29, :324:31
    _GEN_165 = rob_tail == 5'h9;	// rob.scala:228:29, :324:31
    _GEN_166 = io_enq_valids_0 & _GEN_165;	// rob.scala:307:32, :323:29, :324:31
    _GEN_167 = rob_tail == 5'hA;	// rob.scala:228:29, :324:31
    _GEN_168 = io_enq_valids_0 & _GEN_167;	// rob.scala:307:32, :323:29, :324:31
    _GEN_169 = rob_tail == 5'hB;	// rob.scala:228:29, :324:31
    _GEN_170 = io_enq_valids_0 & _GEN_169;	// rob.scala:307:32, :323:29, :324:31
    _GEN_171 = rob_tail == 5'hC;	// rob.scala:228:29, :324:31
    _GEN_172 = io_enq_valids_0 & _GEN_171;	// rob.scala:307:32, :323:29, :324:31
    _GEN_173 = rob_tail == 5'hD;	// rob.scala:228:29, :324:31
    _GEN_174 = io_enq_valids_0 & _GEN_173;	// rob.scala:307:32, :323:29, :324:31
    _GEN_175 = rob_tail == 5'hE;	// rob.scala:228:29, :324:31
    _GEN_176 = io_enq_valids_0 & _GEN_175;	// rob.scala:307:32, :323:29, :324:31
    _GEN_177 = rob_tail == 5'hF;	// rob.scala:228:29, :324:31
    _GEN_178 = io_enq_valids_0 & _GEN_177;	// rob.scala:307:32, :323:29, :324:31
    _GEN_179 = rob_tail == 5'h10;	// rob.scala:228:29, :324:31
    _GEN_180 = io_enq_valids_0 & _GEN_179;	// rob.scala:307:32, :323:29, :324:31
    _GEN_181 = rob_tail == 5'h11;	// rob.scala:228:29, :324:31
    _GEN_182 = io_enq_valids_0 & _GEN_181;	// rob.scala:307:32, :323:29, :324:31
    _GEN_183 = rob_tail == 5'h12;	// rob.scala:228:29, :324:31
    _GEN_184 = io_enq_valids_0 & _GEN_183;	// rob.scala:307:32, :323:29, :324:31
    _GEN_185 = rob_tail == 5'h13;	// rob.scala:228:29, :324:31
    _GEN_186 = io_enq_valids_0 & _GEN_185;	// rob.scala:307:32, :323:29, :324:31
    _GEN_187 = rob_tail == 5'h14;	// rob.scala:228:29, :324:31
    _GEN_188 = io_enq_valids_0 & _GEN_187;	// rob.scala:307:32, :323:29, :324:31
    _GEN_189 = rob_tail == 5'h15;	// rob.scala:228:29, :324:31
    _GEN_190 = io_enq_valids_0 & _GEN_189;	// rob.scala:307:32, :323:29, :324:31
    _GEN_191 = rob_tail == 5'h16;	// rob.scala:228:29, :324:31
    _GEN_192 = io_enq_valids_0 & _GEN_191;	// rob.scala:307:32, :323:29, :324:31
    _GEN_193 = rob_tail == 5'h17;	// rob.scala:228:29, :324:31
    _GEN_194 = io_enq_valids_0 & _GEN_193;	// rob.scala:307:32, :323:29, :324:31
    _GEN_195 = rob_tail == 5'h18;	// rob.scala:228:29, :324:31
    _GEN_196 = io_enq_valids_0 & _GEN_195;	// rob.scala:307:32, :323:29, :324:31
    _GEN_197 = rob_tail == 5'h19;	// rob.scala:228:29, :324:31
    _GEN_198 = io_enq_valids_0 & _GEN_197;	// rob.scala:307:32, :323:29, :324:31
    _GEN_199 = rob_tail == 5'h1A;	// rob.scala:228:29, :324:31
    _GEN_200 = io_enq_valids_0 & _GEN_199;	// rob.scala:307:32, :323:29, :324:31
    _GEN_201 = rob_tail == 5'h1B;	// rob.scala:228:29, :324:31
    _GEN_202 = io_enq_valids_0 & _GEN_201;	// rob.scala:307:32, :323:29, :324:31
    _GEN_203 = rob_tail == 5'h1C;	// rob.scala:228:29, :324:31
    _GEN_204 = io_enq_valids_0 & _GEN_203;	// rob.scala:307:32, :323:29, :324:31
    _GEN_205 = rob_tail == 5'h1D;	// rob.scala:228:29, :324:31
    _GEN_206 = io_enq_valids_0 & _GEN_205;	// rob.scala:307:32, :323:29, :324:31
    _GEN_207 = rob_tail == 5'h1E;	// rob.scala:228:29, :324:31
    _GEN_208 = io_enq_valids_0 & _GEN_207;	// rob.scala:307:32, :323:29, :324:31
    _GEN_209 = io_enq_valids_0 & (&rob_tail);	// rob.scala:228:29, :307:32, :323:29, :324:31
    _GEN_210 = _GEN_148 ? ~_rob_bsy_T : rob_bsy_0;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_211 = _GEN_150 ? ~_rob_bsy_T : rob_bsy_1;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_212 = _GEN_152 ? ~_rob_bsy_T : rob_bsy_2;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_213 = _GEN_154 ? ~_rob_bsy_T : rob_bsy_3;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_214 = _GEN_156 ? ~_rob_bsy_T : rob_bsy_4;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_215 = _GEN_158 ? ~_rob_bsy_T : rob_bsy_5;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_216 = _GEN_160 ? ~_rob_bsy_T : rob_bsy_6;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_217 = _GEN_162 ? ~_rob_bsy_T : rob_bsy_7;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_218 = _GEN_164 ? ~_rob_bsy_T : rob_bsy_8;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_219 = _GEN_166 ? ~_rob_bsy_T : rob_bsy_9;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_220 = _GEN_168 ? ~_rob_bsy_T : rob_bsy_10;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_221 = _GEN_170 ? ~_rob_bsy_T : rob_bsy_11;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_222 = _GEN_172 ? ~_rob_bsy_T : rob_bsy_12;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_223 = _GEN_174 ? ~_rob_bsy_T : rob_bsy_13;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_224 = _GEN_176 ? ~_rob_bsy_T : rob_bsy_14;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_225 = _GEN_178 ? ~_rob_bsy_T : rob_bsy_15;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_226 = _GEN_180 ? ~_rob_bsy_T : rob_bsy_16;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_227 = _GEN_182 ? ~_rob_bsy_T : rob_bsy_17;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_228 = _GEN_184 ? ~_rob_bsy_T : rob_bsy_18;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_229 = _GEN_186 ? ~_rob_bsy_T : rob_bsy_19;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_230 = _GEN_188 ? ~_rob_bsy_T : rob_bsy_20;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_231 = _GEN_190 ? ~_rob_bsy_T : rob_bsy_21;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_232 = _GEN_192 ? ~_rob_bsy_T : rob_bsy_22;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_233 = _GEN_194 ? ~_rob_bsy_T : rob_bsy_23;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_234 = _GEN_196 ? ~_rob_bsy_T : rob_bsy_24;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_235 = _GEN_198 ? ~_rob_bsy_T : rob_bsy_25;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_236 = _GEN_200 ? ~_rob_bsy_T : rob_bsy_26;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_237 = _GEN_202 ? ~_rob_bsy_T : rob_bsy_27;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_238 = _GEN_204 ? ~_rob_bsy_T : rob_bsy_28;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_239 = _GEN_206 ? ~_rob_bsy_T : rob_bsy_29;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_240 = _GEN_208 ? ~_rob_bsy_T : rob_bsy_30;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_241 = _GEN_209 ? ~_rob_bsy_T : rob_bsy_31;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_242 = _GEN_148 ? _rob_unsafe_T_4 : rob_unsafe_0;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_243 = _GEN_150 ? _rob_unsafe_T_4 : rob_unsafe_1;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_244 = _GEN_152 ? _rob_unsafe_T_4 : rob_unsafe_2;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_245 = _GEN_154 ? _rob_unsafe_T_4 : rob_unsafe_3;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_246 = _GEN_156 ? _rob_unsafe_T_4 : rob_unsafe_4;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_247 = _GEN_158 ? _rob_unsafe_T_4 : rob_unsafe_5;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_248 = _GEN_160 ? _rob_unsafe_T_4 : rob_unsafe_6;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_249 = _GEN_162 ? _rob_unsafe_T_4 : rob_unsafe_7;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_250 = _GEN_164 ? _rob_unsafe_T_4 : rob_unsafe_8;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_251 = _GEN_166 ? _rob_unsafe_T_4 : rob_unsafe_9;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_252 = _GEN_168 ? _rob_unsafe_T_4 : rob_unsafe_10;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_253 = _GEN_170 ? _rob_unsafe_T_4 : rob_unsafe_11;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_254 = _GEN_172 ? _rob_unsafe_T_4 : rob_unsafe_12;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_255 = _GEN_174 ? _rob_unsafe_T_4 : rob_unsafe_13;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_256 = _GEN_176 ? _rob_unsafe_T_4 : rob_unsafe_14;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_257 = _GEN_178 ? _rob_unsafe_T_4 : rob_unsafe_15;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_258 = _GEN_180 ? _rob_unsafe_T_4 : rob_unsafe_16;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_259 = _GEN_182 ? _rob_unsafe_T_4 : rob_unsafe_17;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_260 = _GEN_184 ? _rob_unsafe_T_4 : rob_unsafe_18;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_261 = _GEN_186 ? _rob_unsafe_T_4 : rob_unsafe_19;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_262 = _GEN_188 ? _rob_unsafe_T_4 : rob_unsafe_20;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_263 = _GEN_190 ? _rob_unsafe_T_4 : rob_unsafe_21;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_264 = _GEN_192 ? _rob_unsafe_T_4 : rob_unsafe_22;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_265 = _GEN_194 ? _rob_unsafe_T_4 : rob_unsafe_23;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_266 = _GEN_196 ? _rob_unsafe_T_4 : rob_unsafe_24;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_267 = _GEN_198 ? _rob_unsafe_T_4 : rob_unsafe_25;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_268 = _GEN_200 ? _rob_unsafe_T_4 : rob_unsafe_26;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_269 = _GEN_202 ? _rob_unsafe_T_4 : rob_unsafe_27;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_270 = _GEN_204 ? _rob_unsafe_T_4 : rob_unsafe_28;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_271 = _GEN_206 ? _rob_unsafe_T_4 : rob_unsafe_29;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_272 = _GEN_208 ? _rob_unsafe_T_4 : rob_unsafe_30;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_273 = _GEN_209 ? _rob_unsafe_T_4 : rob_unsafe_31;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_339 = _GEN_1 ? ~_GEN_338 & _GEN_210 : ~_GEN_275 & _GEN_210;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_342 = _GEN_1 ? ~_GEN_341 & _GEN_211 : ~_GEN_277 & _GEN_211;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_345 = _GEN_1 ? ~_GEN_344 & _GEN_212 : ~_GEN_279 & _GEN_212;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_348 = _GEN_1 ? ~_GEN_347 & _GEN_213 : ~_GEN_281 & _GEN_213;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_351 = _GEN_1 ? ~_GEN_350 & _GEN_214 : ~_GEN_283 & _GEN_214;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_354 = _GEN_1 ? ~_GEN_353 & _GEN_215 : ~_GEN_285 & _GEN_215;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_357 = _GEN_1 ? ~_GEN_356 & _GEN_216 : ~_GEN_287 & _GEN_216;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_360 = _GEN_1 ? ~_GEN_359 & _GEN_217 : ~_GEN_289 & _GEN_217;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_363 = _GEN_1 ? ~_GEN_362 & _GEN_218 : ~_GEN_291 & _GEN_218;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_366 = _GEN_1 ? ~_GEN_365 & _GEN_219 : ~_GEN_293 & _GEN_219;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_369 = _GEN_1 ? ~_GEN_368 & _GEN_220 : ~_GEN_295 & _GEN_220;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_372 = _GEN_1 ? ~_GEN_371 & _GEN_221 : ~_GEN_297 & _GEN_221;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_375 = _GEN_1 ? ~_GEN_374 & _GEN_222 : ~_GEN_299 & _GEN_222;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_378 = _GEN_1 ? ~_GEN_377 & _GEN_223 : ~_GEN_301 & _GEN_223;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_381 = _GEN_1 ? ~_GEN_380 & _GEN_224 : ~_GEN_303 & _GEN_224;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_384 = _GEN_1 ? ~_GEN_383 & _GEN_225 : ~_GEN_305 & _GEN_225;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_387 = _GEN_1 ? ~_GEN_386 & _GEN_226 : ~_GEN_307 & _GEN_226;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_390 = _GEN_1 ? ~_GEN_389 & _GEN_227 : ~_GEN_309 & _GEN_227;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_393 = _GEN_1 ? ~_GEN_392 & _GEN_228 : ~_GEN_311 & _GEN_228;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_396 = _GEN_1 ? ~_GEN_395 & _GEN_229 : ~_GEN_313 & _GEN_229;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_399 = _GEN_1 ? ~_GEN_398 & _GEN_230 : ~_GEN_315 & _GEN_230;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_402 = _GEN_1 ? ~_GEN_401 & _GEN_231 : ~_GEN_317 & _GEN_231;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_405 = _GEN_1 ? ~_GEN_404 & _GEN_232 : ~_GEN_319 & _GEN_232;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_408 = _GEN_1 ? ~_GEN_407 & _GEN_233 : ~_GEN_321 & _GEN_233;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_411 = _GEN_1 ? ~_GEN_410 & _GEN_234 : ~_GEN_323 & _GEN_234;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_414 = _GEN_1 ? ~_GEN_413 & _GEN_235 : ~_GEN_325 & _GEN_235;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_417 = _GEN_1 ? ~_GEN_416 & _GEN_236 : ~_GEN_327 & _GEN_236;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_420 = _GEN_1 ? ~_GEN_419 & _GEN_237 : ~_GEN_329 & _GEN_237;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_423 = _GEN_1 ? ~_GEN_422 & _GEN_238 : ~_GEN_331 & _GEN_238;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_426 = _GEN_1 ? ~_GEN_425 & _GEN_239 : ~_GEN_333 & _GEN_239;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_429 = _GEN_1 ? ~_GEN_428 & _GEN_240 : ~_GEN_335 & _GEN_240;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_431 = _GEN_1 ? ~_GEN_430 & _GEN_241 : ~_GEN_336 & _GEN_241;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_432 = _GEN_1 ? ~_GEN_338 & _GEN_242 : ~_GEN_275 & _GEN_242;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_433 = _GEN_1 ? ~_GEN_341 & _GEN_243 : ~_GEN_277 & _GEN_243;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_434 = _GEN_1 ? ~_GEN_344 & _GEN_244 : ~_GEN_279 & _GEN_244;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_435 = _GEN_1 ? ~_GEN_347 & _GEN_245 : ~_GEN_281 & _GEN_245;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_436 = _GEN_1 ? ~_GEN_350 & _GEN_246 : ~_GEN_283 & _GEN_246;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_437 = _GEN_1 ? ~_GEN_353 & _GEN_247 : ~_GEN_285 & _GEN_247;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_438 = _GEN_1 ? ~_GEN_356 & _GEN_248 : ~_GEN_287 & _GEN_248;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_439 = _GEN_1 ? ~_GEN_359 & _GEN_249 : ~_GEN_289 & _GEN_249;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_440 = _GEN_1 ? ~_GEN_362 & _GEN_250 : ~_GEN_291 & _GEN_250;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_441 = _GEN_1 ? ~_GEN_365 & _GEN_251 : ~_GEN_293 & _GEN_251;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_442 = _GEN_1 ? ~_GEN_368 & _GEN_252 : ~_GEN_295 & _GEN_252;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_443 = _GEN_1 ? ~_GEN_371 & _GEN_253 : ~_GEN_297 & _GEN_253;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_444 = _GEN_1 ? ~_GEN_374 & _GEN_254 : ~_GEN_299 & _GEN_254;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_445 = _GEN_1 ? ~_GEN_377 & _GEN_255 : ~_GEN_301 & _GEN_255;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_446 = _GEN_1 ? ~_GEN_380 & _GEN_256 : ~_GEN_303 & _GEN_256;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_447 = _GEN_1 ? ~_GEN_383 & _GEN_257 : ~_GEN_305 & _GEN_257;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_448 = _GEN_1 ? ~_GEN_386 & _GEN_258 : ~_GEN_307 & _GEN_258;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_449 = _GEN_1 ? ~_GEN_389 & _GEN_259 : ~_GEN_309 & _GEN_259;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_450 = _GEN_1 ? ~_GEN_392 & _GEN_260 : ~_GEN_311 & _GEN_260;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_451 = _GEN_1 ? ~_GEN_395 & _GEN_261 : ~_GEN_313 & _GEN_261;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_452 = _GEN_1 ? ~_GEN_398 & _GEN_262 : ~_GEN_315 & _GEN_262;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_453 = _GEN_1 ? ~_GEN_401 & _GEN_263 : ~_GEN_317 & _GEN_263;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_454 = _GEN_1 ? ~_GEN_404 & _GEN_264 : ~_GEN_319 & _GEN_264;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_455 = _GEN_1 ? ~_GEN_407 & _GEN_265 : ~_GEN_321 & _GEN_265;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_456 = _GEN_1 ? ~_GEN_410 & _GEN_266 : ~_GEN_323 & _GEN_266;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_457 = _GEN_1 ? ~_GEN_413 & _GEN_267 : ~_GEN_325 & _GEN_267;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_458 = _GEN_1 ? ~_GEN_416 & _GEN_268 : ~_GEN_327 & _GEN_268;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_459 = _GEN_1 ? ~_GEN_419 & _GEN_269 : ~_GEN_329 & _GEN_269;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_460 = _GEN_1 ? ~_GEN_422 & _GEN_270 : ~_GEN_331 & _GEN_270;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_461 = _GEN_1 ? ~_GEN_425 & _GEN_271 : ~_GEN_333 & _GEN_271;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_462 = _GEN_1 ? ~_GEN_428 & _GEN_272 : ~_GEN_335 & _GEN_272;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_463 = _GEN_1 ? ~_GEN_430 & _GEN_273 : ~_GEN_336 & _GEN_273;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_529 = _GEN_3 ? ~_GEN_528 & _GEN_339 : ~_GEN_465 & _GEN_339;	// rob.scala:346:{27,69}, :347:31
    _GEN_532 = _GEN_3 ? ~_GEN_531 & _GEN_342 : ~_GEN_467 & _GEN_342;	// rob.scala:346:{27,69}, :347:31
    _GEN_535 = _GEN_3 ? ~_GEN_534 & _GEN_345 : ~_GEN_469 & _GEN_345;	// rob.scala:346:{27,69}, :347:31
    _GEN_538 = _GEN_3 ? ~_GEN_537 & _GEN_348 : ~_GEN_471 & _GEN_348;	// rob.scala:346:{27,69}, :347:31
    _GEN_541 = _GEN_3 ? ~_GEN_540 & _GEN_351 : ~_GEN_473 & _GEN_351;	// rob.scala:346:{27,69}, :347:31
    _GEN_544 = _GEN_3 ? ~_GEN_543 & _GEN_354 : ~_GEN_475 & _GEN_354;	// rob.scala:346:{27,69}, :347:31
    _GEN_547 = _GEN_3 ? ~_GEN_546 & _GEN_357 : ~_GEN_477 & _GEN_357;	// rob.scala:346:{27,69}, :347:31
    _GEN_550 = _GEN_3 ? ~_GEN_549 & _GEN_360 : ~_GEN_479 & _GEN_360;	// rob.scala:346:{27,69}, :347:31
    _GEN_553 = _GEN_3 ? ~_GEN_552 & _GEN_363 : ~_GEN_481 & _GEN_363;	// rob.scala:346:{27,69}, :347:31
    _GEN_556 = _GEN_3 ? ~_GEN_555 & _GEN_366 : ~_GEN_483 & _GEN_366;	// rob.scala:346:{27,69}, :347:31
    _GEN_559 = _GEN_3 ? ~_GEN_558 & _GEN_369 : ~_GEN_485 & _GEN_369;	// rob.scala:346:{27,69}, :347:31
    _GEN_562 = _GEN_3 ? ~_GEN_561 & _GEN_372 : ~_GEN_487 & _GEN_372;	// rob.scala:346:{27,69}, :347:31
    _GEN_565 = _GEN_3 ? ~_GEN_564 & _GEN_375 : ~_GEN_489 & _GEN_375;	// rob.scala:346:{27,69}, :347:31
    _GEN_568 = _GEN_3 ? ~_GEN_567 & _GEN_378 : ~_GEN_491 & _GEN_378;	// rob.scala:346:{27,69}, :347:31
    _GEN_571 = _GEN_3 ? ~_GEN_570 & _GEN_381 : ~_GEN_493 & _GEN_381;	// rob.scala:346:{27,69}, :347:31
    _GEN_574 = _GEN_3 ? ~_GEN_573 & _GEN_384 : ~_GEN_495 & _GEN_384;	// rob.scala:346:{27,69}, :347:31
    _GEN_577 = _GEN_3 ? ~_GEN_576 & _GEN_387 : ~_GEN_497 & _GEN_387;	// rob.scala:346:{27,69}, :347:31
    _GEN_580 = _GEN_3 ? ~_GEN_579 & _GEN_390 : ~_GEN_499 & _GEN_390;	// rob.scala:346:{27,69}, :347:31
    _GEN_583 = _GEN_3 ? ~_GEN_582 & _GEN_393 : ~_GEN_501 & _GEN_393;	// rob.scala:346:{27,69}, :347:31
    _GEN_586 = _GEN_3 ? ~_GEN_585 & _GEN_396 : ~_GEN_503 & _GEN_396;	// rob.scala:346:{27,69}, :347:31
    _GEN_589 = _GEN_3 ? ~_GEN_588 & _GEN_399 : ~_GEN_505 & _GEN_399;	// rob.scala:346:{27,69}, :347:31
    _GEN_592 = _GEN_3 ? ~_GEN_591 & _GEN_402 : ~_GEN_507 & _GEN_402;	// rob.scala:346:{27,69}, :347:31
    _GEN_595 = _GEN_3 ? ~_GEN_594 & _GEN_405 : ~_GEN_509 & _GEN_405;	// rob.scala:346:{27,69}, :347:31
    _GEN_598 = _GEN_3 ? ~_GEN_597 & _GEN_408 : ~_GEN_511 & _GEN_408;	// rob.scala:346:{27,69}, :347:31
    _GEN_601 = _GEN_3 ? ~_GEN_600 & _GEN_411 : ~_GEN_513 & _GEN_411;	// rob.scala:346:{27,69}, :347:31
    _GEN_604 = _GEN_3 ? ~_GEN_603 & _GEN_414 : ~_GEN_515 & _GEN_414;	// rob.scala:346:{27,69}, :347:31
    _GEN_607 = _GEN_3 ? ~_GEN_606 & _GEN_417 : ~_GEN_517 & _GEN_417;	// rob.scala:346:{27,69}, :347:31
    _GEN_610 = _GEN_3 ? ~_GEN_609 & _GEN_420 : ~_GEN_519 & _GEN_420;	// rob.scala:346:{27,69}, :347:31
    _GEN_613 = _GEN_3 ? ~_GEN_612 & _GEN_423 : ~_GEN_521 & _GEN_423;	// rob.scala:346:{27,69}, :347:31
    _GEN_616 = _GEN_3 ? ~_GEN_615 & _GEN_426 : ~_GEN_523 & _GEN_426;	// rob.scala:346:{27,69}, :347:31
    _GEN_619 = _GEN_3 ? ~_GEN_618 & _GEN_429 : ~_GEN_525 & _GEN_429;	// rob.scala:346:{27,69}, :347:31
    _GEN_621 = _GEN_3 ? ~_GEN_620 & _GEN_431 : ~_GEN_526 & _GEN_431;	// rob.scala:346:{27,69}, :347:31
    _GEN_622 = _GEN_3 ? ~_GEN_528 & _GEN_432 : ~_GEN_465 & _GEN_432;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_623 = _GEN_3 ? ~_GEN_531 & _GEN_433 : ~_GEN_467 & _GEN_433;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_624 = _GEN_3 ? ~_GEN_534 & _GEN_434 : ~_GEN_469 & _GEN_434;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_625 = _GEN_3 ? ~_GEN_537 & _GEN_435 : ~_GEN_471 & _GEN_435;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_626 = _GEN_3 ? ~_GEN_540 & _GEN_436 : ~_GEN_473 & _GEN_436;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_627 = _GEN_3 ? ~_GEN_543 & _GEN_437 : ~_GEN_475 & _GEN_437;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_628 = _GEN_3 ? ~_GEN_546 & _GEN_438 : ~_GEN_477 & _GEN_438;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_629 = _GEN_3 ? ~_GEN_549 & _GEN_439 : ~_GEN_479 & _GEN_439;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_630 = _GEN_3 ? ~_GEN_552 & _GEN_440 : ~_GEN_481 & _GEN_440;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_631 = _GEN_3 ? ~_GEN_555 & _GEN_441 : ~_GEN_483 & _GEN_441;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_632 = _GEN_3 ? ~_GEN_558 & _GEN_442 : ~_GEN_485 & _GEN_442;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_633 = _GEN_3 ? ~_GEN_561 & _GEN_443 : ~_GEN_487 & _GEN_443;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_634 = _GEN_3 ? ~_GEN_564 & _GEN_444 : ~_GEN_489 & _GEN_444;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_635 = _GEN_3 ? ~_GEN_567 & _GEN_445 : ~_GEN_491 & _GEN_445;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_636 = _GEN_3 ? ~_GEN_570 & _GEN_446 : ~_GEN_493 & _GEN_446;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_637 = _GEN_3 ? ~_GEN_573 & _GEN_447 : ~_GEN_495 & _GEN_447;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_638 = _GEN_3 ? ~_GEN_576 & _GEN_448 : ~_GEN_497 & _GEN_448;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_639 = _GEN_3 ? ~_GEN_579 & _GEN_449 : ~_GEN_499 & _GEN_449;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_640 = _GEN_3 ? ~_GEN_582 & _GEN_450 : ~_GEN_501 & _GEN_450;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_641 = _GEN_3 ? ~_GEN_585 & _GEN_451 : ~_GEN_503 & _GEN_451;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_642 = _GEN_3 ? ~_GEN_588 & _GEN_452 : ~_GEN_505 & _GEN_452;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_643 = _GEN_3 ? ~_GEN_591 & _GEN_453 : ~_GEN_507 & _GEN_453;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_644 = _GEN_3 ? ~_GEN_594 & _GEN_454 : ~_GEN_509 & _GEN_454;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_645 = _GEN_3 ? ~_GEN_597 & _GEN_455 : ~_GEN_511 & _GEN_455;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_646 = _GEN_3 ? ~_GEN_600 & _GEN_456 : ~_GEN_513 & _GEN_456;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_647 = _GEN_3 ? ~_GEN_603 & _GEN_457 : ~_GEN_515 & _GEN_457;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_648 = _GEN_3 ? ~_GEN_606 & _GEN_458 : ~_GEN_517 & _GEN_458;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_649 = _GEN_3 ? ~_GEN_609 & _GEN_459 : ~_GEN_519 & _GEN_459;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_650 = _GEN_3 ? ~_GEN_612 & _GEN_460 : ~_GEN_521 & _GEN_460;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_651 = _GEN_3 ? ~_GEN_615 & _GEN_461 : ~_GEN_523 & _GEN_461;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_652 = _GEN_3 ? ~_GEN_618 & _GEN_462 : ~_GEN_525 & _GEN_462;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_653 = _GEN_3 ? ~_GEN_620 & _GEN_463 : ~_GEN_526 & _GEN_463;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_719 = _GEN_5 ? ~_GEN_718 & _GEN_529 : ~_GEN_655 & _GEN_529;	// rob.scala:346:{27,69}, :347:31
    _GEN_722 = _GEN_5 ? ~_GEN_721 & _GEN_532 : ~_GEN_657 & _GEN_532;	// rob.scala:346:{27,69}, :347:31
    _GEN_725 = _GEN_5 ? ~_GEN_724 & _GEN_535 : ~_GEN_659 & _GEN_535;	// rob.scala:346:{27,69}, :347:31
    _GEN_728 = _GEN_5 ? ~_GEN_727 & _GEN_538 : ~_GEN_661 & _GEN_538;	// rob.scala:346:{27,69}, :347:31
    _GEN_731 = _GEN_5 ? ~_GEN_730 & _GEN_541 : ~_GEN_663 & _GEN_541;	// rob.scala:346:{27,69}, :347:31
    _GEN_734 = _GEN_5 ? ~_GEN_733 & _GEN_544 : ~_GEN_665 & _GEN_544;	// rob.scala:346:{27,69}, :347:31
    _GEN_737 = _GEN_5 ? ~_GEN_736 & _GEN_547 : ~_GEN_667 & _GEN_547;	// rob.scala:346:{27,69}, :347:31
    _GEN_740 = _GEN_5 ? ~_GEN_739 & _GEN_550 : ~_GEN_669 & _GEN_550;	// rob.scala:346:{27,69}, :347:31
    _GEN_743 = _GEN_5 ? ~_GEN_742 & _GEN_553 : ~_GEN_671 & _GEN_553;	// rob.scala:346:{27,69}, :347:31
    _GEN_746 = _GEN_5 ? ~_GEN_745 & _GEN_556 : ~_GEN_673 & _GEN_556;	// rob.scala:346:{27,69}, :347:31
    _GEN_749 = _GEN_5 ? ~_GEN_748 & _GEN_559 : ~_GEN_675 & _GEN_559;	// rob.scala:346:{27,69}, :347:31
    _GEN_752 = _GEN_5 ? ~_GEN_751 & _GEN_562 : ~_GEN_677 & _GEN_562;	// rob.scala:346:{27,69}, :347:31
    _GEN_755 = _GEN_5 ? ~_GEN_754 & _GEN_565 : ~_GEN_679 & _GEN_565;	// rob.scala:346:{27,69}, :347:31
    _GEN_758 = _GEN_5 ? ~_GEN_757 & _GEN_568 : ~_GEN_681 & _GEN_568;	// rob.scala:346:{27,69}, :347:31
    _GEN_761 = _GEN_5 ? ~_GEN_760 & _GEN_571 : ~_GEN_683 & _GEN_571;	// rob.scala:346:{27,69}, :347:31
    _GEN_764 = _GEN_5 ? ~_GEN_763 & _GEN_574 : ~_GEN_685 & _GEN_574;	// rob.scala:346:{27,69}, :347:31
    _GEN_767 = _GEN_5 ? ~_GEN_766 & _GEN_577 : ~_GEN_687 & _GEN_577;	// rob.scala:346:{27,69}, :347:31
    _GEN_770 = _GEN_5 ? ~_GEN_769 & _GEN_580 : ~_GEN_689 & _GEN_580;	// rob.scala:346:{27,69}, :347:31
    _GEN_773 = _GEN_5 ? ~_GEN_772 & _GEN_583 : ~_GEN_691 & _GEN_583;	// rob.scala:346:{27,69}, :347:31
    _GEN_776 = _GEN_5 ? ~_GEN_775 & _GEN_586 : ~_GEN_693 & _GEN_586;	// rob.scala:346:{27,69}, :347:31
    _GEN_779 = _GEN_5 ? ~_GEN_778 & _GEN_589 : ~_GEN_695 & _GEN_589;	// rob.scala:346:{27,69}, :347:31
    _GEN_782 = _GEN_5 ? ~_GEN_781 & _GEN_592 : ~_GEN_697 & _GEN_592;	// rob.scala:346:{27,69}, :347:31
    _GEN_785 = _GEN_5 ? ~_GEN_784 & _GEN_595 : ~_GEN_699 & _GEN_595;	// rob.scala:346:{27,69}, :347:31
    _GEN_788 = _GEN_5 ? ~_GEN_787 & _GEN_598 : ~_GEN_701 & _GEN_598;	// rob.scala:346:{27,69}, :347:31
    _GEN_791 = _GEN_5 ? ~_GEN_790 & _GEN_601 : ~_GEN_703 & _GEN_601;	// rob.scala:346:{27,69}, :347:31
    _GEN_794 = _GEN_5 ? ~_GEN_793 & _GEN_604 : ~_GEN_705 & _GEN_604;	// rob.scala:346:{27,69}, :347:31
    _GEN_797 = _GEN_5 ? ~_GEN_796 & _GEN_607 : ~_GEN_707 & _GEN_607;	// rob.scala:346:{27,69}, :347:31
    _GEN_800 = _GEN_5 ? ~_GEN_799 & _GEN_610 : ~_GEN_709 & _GEN_610;	// rob.scala:346:{27,69}, :347:31
    _GEN_803 = _GEN_5 ? ~_GEN_802 & _GEN_613 : ~_GEN_711 & _GEN_613;	// rob.scala:346:{27,69}, :347:31
    _GEN_806 = _GEN_5 ? ~_GEN_805 & _GEN_616 : ~_GEN_713 & _GEN_616;	// rob.scala:346:{27,69}, :347:31
    _GEN_809 = _GEN_5 ? ~_GEN_808 & _GEN_619 : ~_GEN_715 & _GEN_619;	// rob.scala:346:{27,69}, :347:31
    _GEN_811 = _GEN_5 ? ~_GEN_810 & _GEN_621 : ~_GEN_716 & _GEN_621;	// rob.scala:346:{27,69}, :347:31
    _GEN_812 = _GEN_5 ? ~_GEN_718 & _GEN_622 : ~_GEN_655 & _GEN_622;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_813 = _GEN_5 ? ~_GEN_721 & _GEN_623 : ~_GEN_657 & _GEN_623;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_814 = _GEN_5 ? ~_GEN_724 & _GEN_624 : ~_GEN_659 & _GEN_624;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_815 = _GEN_5 ? ~_GEN_727 & _GEN_625 : ~_GEN_661 & _GEN_625;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_816 = _GEN_5 ? ~_GEN_730 & _GEN_626 : ~_GEN_663 & _GEN_626;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_817 = _GEN_5 ? ~_GEN_733 & _GEN_627 : ~_GEN_665 & _GEN_627;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_818 = _GEN_5 ? ~_GEN_736 & _GEN_628 : ~_GEN_667 & _GEN_628;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_819 = _GEN_5 ? ~_GEN_739 & _GEN_629 : ~_GEN_669 & _GEN_629;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_820 = _GEN_5 ? ~_GEN_742 & _GEN_630 : ~_GEN_671 & _GEN_630;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_821 = _GEN_5 ? ~_GEN_745 & _GEN_631 : ~_GEN_673 & _GEN_631;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_822 = _GEN_5 ? ~_GEN_748 & _GEN_632 : ~_GEN_675 & _GEN_632;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_823 = _GEN_5 ? ~_GEN_751 & _GEN_633 : ~_GEN_677 & _GEN_633;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_824 = _GEN_5 ? ~_GEN_754 & _GEN_634 : ~_GEN_679 & _GEN_634;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_825 = _GEN_5 ? ~_GEN_757 & _GEN_635 : ~_GEN_681 & _GEN_635;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_826 = _GEN_5 ? ~_GEN_760 & _GEN_636 : ~_GEN_683 & _GEN_636;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_827 = _GEN_5 ? ~_GEN_763 & _GEN_637 : ~_GEN_685 & _GEN_637;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_828 = _GEN_5 ? ~_GEN_766 & _GEN_638 : ~_GEN_687 & _GEN_638;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_829 = _GEN_5 ? ~_GEN_769 & _GEN_639 : ~_GEN_689 & _GEN_639;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_830 = _GEN_5 ? ~_GEN_772 & _GEN_640 : ~_GEN_691 & _GEN_640;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_831 = _GEN_5 ? ~_GEN_775 & _GEN_641 : ~_GEN_693 & _GEN_641;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_832 = _GEN_5 ? ~_GEN_778 & _GEN_642 : ~_GEN_695 & _GEN_642;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_833 = _GEN_5 ? ~_GEN_781 & _GEN_643 : ~_GEN_697 & _GEN_643;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_834 = _GEN_5 ? ~_GEN_784 & _GEN_644 : ~_GEN_699 & _GEN_644;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_835 = _GEN_5 ? ~_GEN_787 & _GEN_645 : ~_GEN_701 & _GEN_645;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_836 = _GEN_5 ? ~_GEN_790 & _GEN_646 : ~_GEN_703 & _GEN_646;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_837 = _GEN_5 ? ~_GEN_793 & _GEN_647 : ~_GEN_705 & _GEN_647;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_838 = _GEN_5 ? ~_GEN_796 & _GEN_648 : ~_GEN_707 & _GEN_648;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_839 = _GEN_5 ? ~_GEN_799 & _GEN_649 : ~_GEN_709 & _GEN_649;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_840 = _GEN_5 ? ~_GEN_802 & _GEN_650 : ~_GEN_711 & _GEN_650;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_841 = _GEN_5 ? ~_GEN_805 & _GEN_651 : ~_GEN_713 & _GEN_651;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_842 = _GEN_5 ? ~_GEN_808 & _GEN_652 : ~_GEN_715 & _GEN_652;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_843 = _GEN_5 ? ~_GEN_810 & _GEN_653 : ~_GEN_716 & _GEN_653;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_909 = _GEN_7 ? ~_GEN_908 & _GEN_719 : ~_GEN_845 & _GEN_719;	// rob.scala:346:{27,69}, :347:31
    _GEN_912 = _GEN_7 ? ~_GEN_911 & _GEN_722 : ~_GEN_847 & _GEN_722;	// rob.scala:346:{27,69}, :347:31
    _GEN_915 = _GEN_7 ? ~_GEN_914 & _GEN_725 : ~_GEN_849 & _GEN_725;	// rob.scala:346:{27,69}, :347:31
    _GEN_918 = _GEN_7 ? ~_GEN_917 & _GEN_728 : ~_GEN_851 & _GEN_728;	// rob.scala:346:{27,69}, :347:31
    _GEN_921 = _GEN_7 ? ~_GEN_920 & _GEN_731 : ~_GEN_853 & _GEN_731;	// rob.scala:346:{27,69}, :347:31
    _GEN_924 = _GEN_7 ? ~_GEN_923 & _GEN_734 : ~_GEN_855 & _GEN_734;	// rob.scala:346:{27,69}, :347:31
    _GEN_927 = _GEN_7 ? ~_GEN_926 & _GEN_737 : ~_GEN_857 & _GEN_737;	// rob.scala:346:{27,69}, :347:31
    _GEN_930 = _GEN_7 ? ~_GEN_929 & _GEN_740 : ~_GEN_859 & _GEN_740;	// rob.scala:346:{27,69}, :347:31
    _GEN_933 = _GEN_7 ? ~_GEN_932 & _GEN_743 : ~_GEN_861 & _GEN_743;	// rob.scala:346:{27,69}, :347:31
    _GEN_936 = _GEN_7 ? ~_GEN_935 & _GEN_746 : ~_GEN_863 & _GEN_746;	// rob.scala:346:{27,69}, :347:31
    _GEN_939 = _GEN_7 ? ~_GEN_938 & _GEN_749 : ~_GEN_865 & _GEN_749;	// rob.scala:346:{27,69}, :347:31
    _GEN_942 = _GEN_7 ? ~_GEN_941 & _GEN_752 : ~_GEN_867 & _GEN_752;	// rob.scala:346:{27,69}, :347:31
    _GEN_945 = _GEN_7 ? ~_GEN_944 & _GEN_755 : ~_GEN_869 & _GEN_755;	// rob.scala:346:{27,69}, :347:31
    _GEN_948 = _GEN_7 ? ~_GEN_947 & _GEN_758 : ~_GEN_871 & _GEN_758;	// rob.scala:346:{27,69}, :347:31
    _GEN_951 = _GEN_7 ? ~_GEN_950 & _GEN_761 : ~_GEN_873 & _GEN_761;	// rob.scala:346:{27,69}, :347:31
    _GEN_954 = _GEN_7 ? ~_GEN_953 & _GEN_764 : ~_GEN_875 & _GEN_764;	// rob.scala:346:{27,69}, :347:31
    _GEN_957 = _GEN_7 ? ~_GEN_956 & _GEN_767 : ~_GEN_877 & _GEN_767;	// rob.scala:346:{27,69}, :347:31
    _GEN_960 = _GEN_7 ? ~_GEN_959 & _GEN_770 : ~_GEN_879 & _GEN_770;	// rob.scala:346:{27,69}, :347:31
    _GEN_963 = _GEN_7 ? ~_GEN_962 & _GEN_773 : ~_GEN_881 & _GEN_773;	// rob.scala:346:{27,69}, :347:31
    _GEN_966 = _GEN_7 ? ~_GEN_965 & _GEN_776 : ~_GEN_883 & _GEN_776;	// rob.scala:346:{27,69}, :347:31
    _GEN_969 = _GEN_7 ? ~_GEN_968 & _GEN_779 : ~_GEN_885 & _GEN_779;	// rob.scala:346:{27,69}, :347:31
    _GEN_972 = _GEN_7 ? ~_GEN_971 & _GEN_782 : ~_GEN_887 & _GEN_782;	// rob.scala:346:{27,69}, :347:31
    _GEN_975 = _GEN_7 ? ~_GEN_974 & _GEN_785 : ~_GEN_889 & _GEN_785;	// rob.scala:346:{27,69}, :347:31
    _GEN_978 = _GEN_7 ? ~_GEN_977 & _GEN_788 : ~_GEN_891 & _GEN_788;	// rob.scala:346:{27,69}, :347:31
    _GEN_981 = _GEN_7 ? ~_GEN_980 & _GEN_791 : ~_GEN_893 & _GEN_791;	// rob.scala:346:{27,69}, :347:31
    _GEN_984 = _GEN_7 ? ~_GEN_983 & _GEN_794 : ~_GEN_895 & _GEN_794;	// rob.scala:346:{27,69}, :347:31
    _GEN_987 = _GEN_7 ? ~_GEN_986 & _GEN_797 : ~_GEN_897 & _GEN_797;	// rob.scala:346:{27,69}, :347:31
    _GEN_990 = _GEN_7 ? ~_GEN_989 & _GEN_800 : ~_GEN_899 & _GEN_800;	// rob.scala:346:{27,69}, :347:31
    _GEN_993 = _GEN_7 ? ~_GEN_992 & _GEN_803 : ~_GEN_901 & _GEN_803;	// rob.scala:346:{27,69}, :347:31
    _GEN_996 = _GEN_7 ? ~_GEN_995 & _GEN_806 : ~_GEN_903 & _GEN_806;	// rob.scala:346:{27,69}, :347:31
    _GEN_999 = _GEN_7 ? ~_GEN_998 & _GEN_809 : ~_GEN_905 & _GEN_809;	// rob.scala:346:{27,69}, :347:31
    _GEN_1001 = _GEN_7 ? ~_GEN_1000 & _GEN_811 : ~_GEN_906 & _GEN_811;	// rob.scala:346:{27,69}, :347:31
    _GEN_1002 = _GEN_7 ? ~_GEN_908 & _GEN_812 : ~_GEN_845 & _GEN_812;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1003 = _GEN_7 ? ~_GEN_911 & _GEN_813 : ~_GEN_847 & _GEN_813;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1004 = _GEN_7 ? ~_GEN_914 & _GEN_814 : ~_GEN_849 & _GEN_814;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1005 = _GEN_7 ? ~_GEN_917 & _GEN_815 : ~_GEN_851 & _GEN_815;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1006 = _GEN_7 ? ~_GEN_920 & _GEN_816 : ~_GEN_853 & _GEN_816;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1007 = _GEN_7 ? ~_GEN_923 & _GEN_817 : ~_GEN_855 & _GEN_817;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1008 = _GEN_7 ? ~_GEN_926 & _GEN_818 : ~_GEN_857 & _GEN_818;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1009 = _GEN_7 ? ~_GEN_929 & _GEN_819 : ~_GEN_859 & _GEN_819;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1010 = _GEN_7 ? ~_GEN_932 & _GEN_820 : ~_GEN_861 & _GEN_820;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1011 = _GEN_7 ? ~_GEN_935 & _GEN_821 : ~_GEN_863 & _GEN_821;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1012 = _GEN_7 ? ~_GEN_938 & _GEN_822 : ~_GEN_865 & _GEN_822;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1013 = _GEN_7 ? ~_GEN_941 & _GEN_823 : ~_GEN_867 & _GEN_823;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1014 = _GEN_7 ? ~_GEN_944 & _GEN_824 : ~_GEN_869 & _GEN_824;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1015 = _GEN_7 ? ~_GEN_947 & _GEN_825 : ~_GEN_871 & _GEN_825;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1016 = _GEN_7 ? ~_GEN_950 & _GEN_826 : ~_GEN_873 & _GEN_826;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1017 = _GEN_7 ? ~_GEN_953 & _GEN_827 : ~_GEN_875 & _GEN_827;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1018 = _GEN_7 ? ~_GEN_956 & _GEN_828 : ~_GEN_877 & _GEN_828;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1019 = _GEN_7 ? ~_GEN_959 & _GEN_829 : ~_GEN_879 & _GEN_829;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1020 = _GEN_7 ? ~_GEN_962 & _GEN_830 : ~_GEN_881 & _GEN_830;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1021 = _GEN_7 ? ~_GEN_965 & _GEN_831 : ~_GEN_883 & _GEN_831;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1022 = _GEN_7 ? ~_GEN_968 & _GEN_832 : ~_GEN_885 & _GEN_832;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1023 = _GEN_7 ? ~_GEN_971 & _GEN_833 : ~_GEN_887 & _GEN_833;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1024 = _GEN_7 ? ~_GEN_974 & _GEN_834 : ~_GEN_889 & _GEN_834;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1025 = _GEN_7 ? ~_GEN_977 & _GEN_835 : ~_GEN_891 & _GEN_835;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1026 = _GEN_7 ? ~_GEN_980 & _GEN_836 : ~_GEN_893 & _GEN_836;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1027 = _GEN_7 ? ~_GEN_983 & _GEN_837 : ~_GEN_895 & _GEN_837;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1028 = _GEN_7 ? ~_GEN_986 & _GEN_838 : ~_GEN_897 & _GEN_838;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1029 = _GEN_7 ? ~_GEN_989 & _GEN_839 : ~_GEN_899 & _GEN_839;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1030 = _GEN_7 ? ~_GEN_992 & _GEN_840 : ~_GEN_901 & _GEN_840;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1031 = _GEN_7 ? ~_GEN_995 & _GEN_841 : ~_GEN_903 & _GEN_841;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1032 = _GEN_7 ? ~_GEN_998 & _GEN_842 : ~_GEN_905 & _GEN_842;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1033 = _GEN_7 ? ~_GEN_1000 & _GEN_843 : ~_GEN_906 & _GEN_843;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1099 = _GEN_9 ? ~_GEN_1098 & _GEN_909 : ~_GEN_1035 & _GEN_909;	// rob.scala:346:{27,69}, :347:31
    _GEN_1102 = _GEN_9 ? ~_GEN_1101 & _GEN_912 : ~_GEN_1037 & _GEN_912;	// rob.scala:346:{27,69}, :347:31
    _GEN_1105 = _GEN_9 ? ~_GEN_1104 & _GEN_915 : ~_GEN_1039 & _GEN_915;	// rob.scala:346:{27,69}, :347:31
    _GEN_1108 = _GEN_9 ? ~_GEN_1107 & _GEN_918 : ~_GEN_1041 & _GEN_918;	// rob.scala:346:{27,69}, :347:31
    _GEN_1111 = _GEN_9 ? ~_GEN_1110 & _GEN_921 : ~_GEN_1043 & _GEN_921;	// rob.scala:346:{27,69}, :347:31
    _GEN_1114 = _GEN_9 ? ~_GEN_1113 & _GEN_924 : ~_GEN_1045 & _GEN_924;	// rob.scala:346:{27,69}, :347:31
    _GEN_1117 = _GEN_9 ? ~_GEN_1116 & _GEN_927 : ~_GEN_1047 & _GEN_927;	// rob.scala:346:{27,69}, :347:31
    _GEN_1120 = _GEN_9 ? ~_GEN_1119 & _GEN_930 : ~_GEN_1049 & _GEN_930;	// rob.scala:346:{27,69}, :347:31
    _GEN_1123 = _GEN_9 ? ~_GEN_1122 & _GEN_933 : ~_GEN_1051 & _GEN_933;	// rob.scala:346:{27,69}, :347:31
    _GEN_1126 = _GEN_9 ? ~_GEN_1125 & _GEN_936 : ~_GEN_1053 & _GEN_936;	// rob.scala:346:{27,69}, :347:31
    _GEN_1129 = _GEN_9 ? ~_GEN_1128 & _GEN_939 : ~_GEN_1055 & _GEN_939;	// rob.scala:346:{27,69}, :347:31
    _GEN_1132 = _GEN_9 ? ~_GEN_1131 & _GEN_942 : ~_GEN_1057 & _GEN_942;	// rob.scala:346:{27,69}, :347:31
    _GEN_1135 = _GEN_9 ? ~_GEN_1134 & _GEN_945 : ~_GEN_1059 & _GEN_945;	// rob.scala:346:{27,69}, :347:31
    _GEN_1138 = _GEN_9 ? ~_GEN_1137 & _GEN_948 : ~_GEN_1061 & _GEN_948;	// rob.scala:346:{27,69}, :347:31
    _GEN_1141 = _GEN_9 ? ~_GEN_1140 & _GEN_951 : ~_GEN_1063 & _GEN_951;	// rob.scala:346:{27,69}, :347:31
    _GEN_1144 = _GEN_9 ? ~_GEN_1143 & _GEN_954 : ~_GEN_1065 & _GEN_954;	// rob.scala:346:{27,69}, :347:31
    _GEN_1147 = _GEN_9 ? ~_GEN_1146 & _GEN_957 : ~_GEN_1067 & _GEN_957;	// rob.scala:346:{27,69}, :347:31
    _GEN_1150 = _GEN_9 ? ~_GEN_1149 & _GEN_960 : ~_GEN_1069 & _GEN_960;	// rob.scala:346:{27,69}, :347:31
    _GEN_1153 = _GEN_9 ? ~_GEN_1152 & _GEN_963 : ~_GEN_1071 & _GEN_963;	// rob.scala:346:{27,69}, :347:31
    _GEN_1156 = _GEN_9 ? ~_GEN_1155 & _GEN_966 : ~_GEN_1073 & _GEN_966;	// rob.scala:346:{27,69}, :347:31
    _GEN_1159 = _GEN_9 ? ~_GEN_1158 & _GEN_969 : ~_GEN_1075 & _GEN_969;	// rob.scala:346:{27,69}, :347:31
    _GEN_1162 = _GEN_9 ? ~_GEN_1161 & _GEN_972 : ~_GEN_1077 & _GEN_972;	// rob.scala:346:{27,69}, :347:31
    _GEN_1165 = _GEN_9 ? ~_GEN_1164 & _GEN_975 : ~_GEN_1079 & _GEN_975;	// rob.scala:346:{27,69}, :347:31
    _GEN_1168 = _GEN_9 ? ~_GEN_1167 & _GEN_978 : ~_GEN_1081 & _GEN_978;	// rob.scala:346:{27,69}, :347:31
    _GEN_1171 = _GEN_9 ? ~_GEN_1170 & _GEN_981 : ~_GEN_1083 & _GEN_981;	// rob.scala:346:{27,69}, :347:31
    _GEN_1174 = _GEN_9 ? ~_GEN_1173 & _GEN_984 : ~_GEN_1085 & _GEN_984;	// rob.scala:346:{27,69}, :347:31
    _GEN_1177 = _GEN_9 ? ~_GEN_1176 & _GEN_987 : ~_GEN_1087 & _GEN_987;	// rob.scala:346:{27,69}, :347:31
    _GEN_1180 = _GEN_9 ? ~_GEN_1179 & _GEN_990 : ~_GEN_1089 & _GEN_990;	// rob.scala:346:{27,69}, :347:31
    _GEN_1183 = _GEN_9 ? ~_GEN_1182 & _GEN_993 : ~_GEN_1091 & _GEN_993;	// rob.scala:346:{27,69}, :347:31
    _GEN_1186 = _GEN_9 ? ~_GEN_1185 & _GEN_996 : ~_GEN_1093 & _GEN_996;	// rob.scala:346:{27,69}, :347:31
    _GEN_1189 = _GEN_9 ? ~_GEN_1188 & _GEN_999 : ~_GEN_1095 & _GEN_999;	// rob.scala:346:{27,69}, :347:31
    _GEN_1191 = _GEN_9 ? ~_GEN_1190 & _GEN_1001 : ~_GEN_1096 & _GEN_1001;	// rob.scala:346:{27,69}, :347:31
    _GEN_1192 = _GEN_9 ? ~_GEN_1098 & _GEN_1002 : ~_GEN_1035 & _GEN_1002;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1193 = _GEN_9 ? ~_GEN_1101 & _GEN_1003 : ~_GEN_1037 & _GEN_1003;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1194 = _GEN_9 ? ~_GEN_1104 & _GEN_1004 : ~_GEN_1039 & _GEN_1004;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1195 = _GEN_9 ? ~_GEN_1107 & _GEN_1005 : ~_GEN_1041 & _GEN_1005;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1196 = _GEN_9 ? ~_GEN_1110 & _GEN_1006 : ~_GEN_1043 & _GEN_1006;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1197 = _GEN_9 ? ~_GEN_1113 & _GEN_1007 : ~_GEN_1045 & _GEN_1007;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1198 = _GEN_9 ? ~_GEN_1116 & _GEN_1008 : ~_GEN_1047 & _GEN_1008;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1199 = _GEN_9 ? ~_GEN_1119 & _GEN_1009 : ~_GEN_1049 & _GEN_1009;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1200 = _GEN_9 ? ~_GEN_1122 & _GEN_1010 : ~_GEN_1051 & _GEN_1010;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1201 = _GEN_9 ? ~_GEN_1125 & _GEN_1011 : ~_GEN_1053 & _GEN_1011;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1202 = _GEN_9 ? ~_GEN_1128 & _GEN_1012 : ~_GEN_1055 & _GEN_1012;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1203 = _GEN_9 ? ~_GEN_1131 & _GEN_1013 : ~_GEN_1057 & _GEN_1013;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1204 = _GEN_9 ? ~_GEN_1134 & _GEN_1014 : ~_GEN_1059 & _GEN_1014;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1205 = _GEN_9 ? ~_GEN_1137 & _GEN_1015 : ~_GEN_1061 & _GEN_1015;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1206 = _GEN_9 ? ~_GEN_1140 & _GEN_1016 : ~_GEN_1063 & _GEN_1016;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1207 = _GEN_9 ? ~_GEN_1143 & _GEN_1017 : ~_GEN_1065 & _GEN_1017;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1208 = _GEN_9 ? ~_GEN_1146 & _GEN_1018 : ~_GEN_1067 & _GEN_1018;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1209 = _GEN_9 ? ~_GEN_1149 & _GEN_1019 : ~_GEN_1069 & _GEN_1019;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1210 = _GEN_9 ? ~_GEN_1152 & _GEN_1020 : ~_GEN_1071 & _GEN_1020;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1211 = _GEN_9 ? ~_GEN_1155 & _GEN_1021 : ~_GEN_1073 & _GEN_1021;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1212 = _GEN_9 ? ~_GEN_1158 & _GEN_1022 : ~_GEN_1075 & _GEN_1022;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1213 = _GEN_9 ? ~_GEN_1161 & _GEN_1023 : ~_GEN_1077 & _GEN_1023;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1214 = _GEN_9 ? ~_GEN_1164 & _GEN_1024 : ~_GEN_1079 & _GEN_1024;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1215 = _GEN_9 ? ~_GEN_1167 & _GEN_1025 : ~_GEN_1081 & _GEN_1025;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1216 = _GEN_9 ? ~_GEN_1170 & _GEN_1026 : ~_GEN_1083 & _GEN_1026;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1217 = _GEN_9 ? ~_GEN_1173 & _GEN_1027 : ~_GEN_1085 & _GEN_1027;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1218 = _GEN_9 ? ~_GEN_1176 & _GEN_1028 : ~_GEN_1087 & _GEN_1028;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1219 = _GEN_9 ? ~_GEN_1179 & _GEN_1029 : ~_GEN_1089 & _GEN_1029;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1220 = _GEN_9 ? ~_GEN_1182 & _GEN_1030 : ~_GEN_1091 & _GEN_1030;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1221 = _GEN_9 ? ~_GEN_1185 & _GEN_1031 : ~_GEN_1093 & _GEN_1031;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1222 = _GEN_9 ? ~_GEN_1188 & _GEN_1032 : ~_GEN_1095 & _GEN_1032;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1223 = _GEN_9 ? ~_GEN_1190 & _GEN_1033 : ~_GEN_1096 & _GEN_1033;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1445 = rbk_row & _GEN_1444;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1447 = rbk_row & _GEN_1446;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1449 = rbk_row & _GEN_1448;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1451 = rbk_row & _GEN_1450;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1453 = rbk_row & _GEN_1452;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1455 = rbk_row & _GEN_1454;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1457 = rbk_row & _GEN_1456;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1459 = rbk_row & _GEN_1458;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1461 = rbk_row & _GEN_1460;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1463 = rbk_row & _GEN_1462;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1465 = rbk_row & _GEN_1464;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1467 = rbk_row & _GEN_1466;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1469 = rbk_row & _GEN_1468;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1471 = rbk_row & _GEN_1470;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1473 = rbk_row & _GEN_1472;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1475 = rbk_row & _GEN_1474;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1477 = rbk_row & _GEN_1476;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1479 = rbk_row & _GEN_1478;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1481 = rbk_row & _GEN_1480;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1483 = rbk_row & _GEN_1482;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1485 = rbk_row & _GEN_1484;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1487 = rbk_row & _GEN_1486;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1489 = rbk_row & _GEN_1488;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1491 = rbk_row & _GEN_1490;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1493 = rbk_row & _GEN_1492;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1495 = rbk_row & _GEN_1494;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1497 = rbk_row & _GEN_1496;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1499 = rbk_row & _GEN_1498;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1501 = rbk_row & _GEN_1500;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1503 = rbk_row & _GEN_1502;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1505 = rbk_row & _GEN_1504;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1506 = rbk_row & (&com_idx);	// rob.scala:236:20, :323:29, :425:44, :433:20, :434:30
    _GEN_1507 = io_brupdate_b1_mispredict_mask & rob_uop_0_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1508 = io_brupdate_b1_mispredict_mask & rob_uop_1_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1509 = io_brupdate_b1_mispredict_mask & rob_uop_2_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1510 = io_brupdate_b1_mispredict_mask & rob_uop_3_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1511 = io_brupdate_b1_mispredict_mask & rob_uop_4_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1512 = io_brupdate_b1_mispredict_mask & rob_uop_5_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1513 = io_brupdate_b1_mispredict_mask & rob_uop_6_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1514 = io_brupdate_b1_mispredict_mask & rob_uop_7_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1515 = io_brupdate_b1_mispredict_mask & rob_uop_8_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1516 = io_brupdate_b1_mispredict_mask & rob_uop_9_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1517 = io_brupdate_b1_mispredict_mask & rob_uop_10_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1518 = io_brupdate_b1_mispredict_mask & rob_uop_11_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1519 = io_brupdate_b1_mispredict_mask & rob_uop_12_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1520 = io_brupdate_b1_mispredict_mask & rob_uop_13_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1521 = io_brupdate_b1_mispredict_mask & rob_uop_14_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1522 = io_brupdate_b1_mispredict_mask & rob_uop_15_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1523 = io_brupdate_b1_mispredict_mask & rob_uop_16_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1524 = io_brupdate_b1_mispredict_mask & rob_uop_17_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1525 = io_brupdate_b1_mispredict_mask & rob_uop_18_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1526 = io_brupdate_b1_mispredict_mask & rob_uop_19_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1527 = io_brupdate_b1_mispredict_mask & rob_uop_20_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1528 = io_brupdate_b1_mispredict_mask & rob_uop_21_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1529 = io_brupdate_b1_mispredict_mask & rob_uop_22_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1530 = io_brupdate_b1_mispredict_mask & rob_uop_23_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1531 = io_brupdate_b1_mispredict_mask & rob_uop_24_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1532 = io_brupdate_b1_mispredict_mask & rob_uop_25_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1533 = io_brupdate_b1_mispredict_mask & rob_uop_26_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1534 = io_brupdate_b1_mispredict_mask & rob_uop_27_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1535 = io_brupdate_b1_mispredict_mask & rob_uop_28_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1536 = io_brupdate_b1_mispredict_mask & rob_uop_29_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1537 = io_brupdate_b1_mispredict_mask & rob_uop_30_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1538 = io_brupdate_b1_mispredict_mask & rob_uop_31_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1539 = io_enq_valids_1 & _GEN_147;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1540 = io_enq_valids_1 & _GEN_149;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1541 = io_enq_valids_1 & _GEN_151;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1542 = io_enq_valids_1 & _GEN_153;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1543 = io_enq_valids_1 & _GEN_155;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1544 = io_enq_valids_1 & _GEN_157;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1545 = io_enq_valids_1 & _GEN_159;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1546 = io_enq_valids_1 & _GEN_161;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1547 = io_enq_valids_1 & _GEN_163;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1548 = io_enq_valids_1 & _GEN_165;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1549 = io_enq_valids_1 & _GEN_167;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1550 = io_enq_valids_1 & _GEN_169;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1551 = io_enq_valids_1 & _GEN_171;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1552 = io_enq_valids_1 & _GEN_173;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1553 = io_enq_valids_1 & _GEN_175;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1554 = io_enq_valids_1 & _GEN_177;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1555 = io_enq_valids_1 & _GEN_179;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1556 = io_enq_valids_1 & _GEN_181;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1557 = io_enq_valids_1 & _GEN_183;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1558 = io_enq_valids_1 & _GEN_185;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1559 = io_enq_valids_1 & _GEN_187;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1560 = io_enq_valids_1 & _GEN_189;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1561 = io_enq_valids_1 & _GEN_191;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1562 = io_enq_valids_1 & _GEN_193;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1563 = io_enq_valids_1 & _GEN_195;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1564 = io_enq_valids_1 & _GEN_197;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1565 = io_enq_valids_1 & _GEN_199;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1566 = io_enq_valids_1 & _GEN_201;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1567 = io_enq_valids_1 & _GEN_203;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1568 = io_enq_valids_1 & _GEN_205;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1569 = io_enq_valids_1 & _GEN_207;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1570 = io_enq_valids_1 & (&rob_tail);	// rob.scala:228:29, :307:32, :323:29, :324:31
    _GEN_1571 = _GEN_1539 ? ~_rob_bsy_T_2 : rob_bsy_1_0;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1572 = _GEN_1540 ? ~_rob_bsy_T_2 : rob_bsy_1_1;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1573 = _GEN_1541 ? ~_rob_bsy_T_2 : rob_bsy_1_2;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1574 = _GEN_1542 ? ~_rob_bsy_T_2 : rob_bsy_1_3;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1575 = _GEN_1543 ? ~_rob_bsy_T_2 : rob_bsy_1_4;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1576 = _GEN_1544 ? ~_rob_bsy_T_2 : rob_bsy_1_5;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1577 = _GEN_1545 ? ~_rob_bsy_T_2 : rob_bsy_1_6;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1578 = _GEN_1546 ? ~_rob_bsy_T_2 : rob_bsy_1_7;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1579 = _GEN_1547 ? ~_rob_bsy_T_2 : rob_bsy_1_8;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1580 = _GEN_1548 ? ~_rob_bsy_T_2 : rob_bsy_1_9;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1581 = _GEN_1549 ? ~_rob_bsy_T_2 : rob_bsy_1_10;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1582 = _GEN_1550 ? ~_rob_bsy_T_2 : rob_bsy_1_11;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1583 = _GEN_1551 ? ~_rob_bsy_T_2 : rob_bsy_1_12;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1584 = _GEN_1552 ? ~_rob_bsy_T_2 : rob_bsy_1_13;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1585 = _GEN_1553 ? ~_rob_bsy_T_2 : rob_bsy_1_14;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1586 = _GEN_1554 ? ~_rob_bsy_T_2 : rob_bsy_1_15;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1587 = _GEN_1555 ? ~_rob_bsy_T_2 : rob_bsy_1_16;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1588 = _GEN_1556 ? ~_rob_bsy_T_2 : rob_bsy_1_17;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1589 = _GEN_1557 ? ~_rob_bsy_T_2 : rob_bsy_1_18;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1590 = _GEN_1558 ? ~_rob_bsy_T_2 : rob_bsy_1_19;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1591 = _GEN_1559 ? ~_rob_bsy_T_2 : rob_bsy_1_20;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1592 = _GEN_1560 ? ~_rob_bsy_T_2 : rob_bsy_1_21;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1593 = _GEN_1561 ? ~_rob_bsy_T_2 : rob_bsy_1_22;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1594 = _GEN_1562 ? ~_rob_bsy_T_2 : rob_bsy_1_23;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1595 = _GEN_1563 ? ~_rob_bsy_T_2 : rob_bsy_1_24;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1596 = _GEN_1564 ? ~_rob_bsy_T_2 : rob_bsy_1_25;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1597 = _GEN_1565 ? ~_rob_bsy_T_2 : rob_bsy_1_26;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1598 = _GEN_1566 ? ~_rob_bsy_T_2 : rob_bsy_1_27;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1599 = _GEN_1567 ? ~_rob_bsy_T_2 : rob_bsy_1_28;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1600 = _GEN_1568 ? ~_rob_bsy_T_2 : rob_bsy_1_29;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1601 = _GEN_1569 ? ~_rob_bsy_T_2 : rob_bsy_1_30;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1602 = _GEN_1570 ? ~_rob_bsy_T_2 : rob_bsy_1_31;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1603 = _GEN_1539 ? _rob_unsafe_T_9 : rob_unsafe_1_0;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1604 = _GEN_1540 ? _rob_unsafe_T_9 : rob_unsafe_1_1;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1605 = _GEN_1541 ? _rob_unsafe_T_9 : rob_unsafe_1_2;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1606 = _GEN_1542 ? _rob_unsafe_T_9 : rob_unsafe_1_3;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1607 = _GEN_1543 ? _rob_unsafe_T_9 : rob_unsafe_1_4;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1608 = _GEN_1544 ? _rob_unsafe_T_9 : rob_unsafe_1_5;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1609 = _GEN_1545 ? _rob_unsafe_T_9 : rob_unsafe_1_6;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1610 = _GEN_1546 ? _rob_unsafe_T_9 : rob_unsafe_1_7;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1611 = _GEN_1547 ? _rob_unsafe_T_9 : rob_unsafe_1_8;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1612 = _GEN_1548 ? _rob_unsafe_T_9 : rob_unsafe_1_9;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1613 = _GEN_1549 ? _rob_unsafe_T_9 : rob_unsafe_1_10;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1614 = _GEN_1550 ? _rob_unsafe_T_9 : rob_unsafe_1_11;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1615 = _GEN_1551 ? _rob_unsafe_T_9 : rob_unsafe_1_12;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1616 = _GEN_1552 ? _rob_unsafe_T_9 : rob_unsafe_1_13;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1617 = _GEN_1553 ? _rob_unsafe_T_9 : rob_unsafe_1_14;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1618 = _GEN_1554 ? _rob_unsafe_T_9 : rob_unsafe_1_15;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1619 = _GEN_1555 ? _rob_unsafe_T_9 : rob_unsafe_1_16;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1620 = _GEN_1556 ? _rob_unsafe_T_9 : rob_unsafe_1_17;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1621 = _GEN_1557 ? _rob_unsafe_T_9 : rob_unsafe_1_18;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1622 = _GEN_1558 ? _rob_unsafe_T_9 : rob_unsafe_1_19;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1623 = _GEN_1559 ? _rob_unsafe_T_9 : rob_unsafe_1_20;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1624 = _GEN_1560 ? _rob_unsafe_T_9 : rob_unsafe_1_21;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1625 = _GEN_1561 ? _rob_unsafe_T_9 : rob_unsafe_1_22;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1626 = _GEN_1562 ? _rob_unsafe_T_9 : rob_unsafe_1_23;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1627 = _GEN_1563 ? _rob_unsafe_T_9 : rob_unsafe_1_24;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1628 = _GEN_1564 ? _rob_unsafe_T_9 : rob_unsafe_1_25;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1629 = _GEN_1565 ? _rob_unsafe_T_9 : rob_unsafe_1_26;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1630 = _GEN_1566 ? _rob_unsafe_T_9 : rob_unsafe_1_27;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1631 = _GEN_1567 ? _rob_unsafe_T_9 : rob_unsafe_1_28;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1632 = _GEN_1568 ? _rob_unsafe_T_9 : rob_unsafe_1_29;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1633 = _GEN_1569 ? _rob_unsafe_T_9 : rob_unsafe_1_30;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1634 = _GEN_1570 ? _rob_unsafe_T_9 : rob_unsafe_1_31;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1668 = _GEN_36 ? ~_GEN_1667 & _GEN_1571 : ~_GEN_1635 & _GEN_1571;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1670 = _GEN_36 ? ~_GEN_1669 & _GEN_1572 : ~_GEN_1636 & _GEN_1572;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1672 = _GEN_36 ? ~_GEN_1671 & _GEN_1573 : ~_GEN_1637 & _GEN_1573;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1674 = _GEN_36 ? ~_GEN_1673 & _GEN_1574 : ~_GEN_1638 & _GEN_1574;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1676 = _GEN_36 ? ~_GEN_1675 & _GEN_1575 : ~_GEN_1639 & _GEN_1575;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1678 = _GEN_36 ? ~_GEN_1677 & _GEN_1576 : ~_GEN_1640 & _GEN_1576;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1680 = _GEN_36 ? ~_GEN_1679 & _GEN_1577 : ~_GEN_1641 & _GEN_1577;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1682 = _GEN_36 ? ~_GEN_1681 & _GEN_1578 : ~_GEN_1642 & _GEN_1578;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1684 = _GEN_36 ? ~_GEN_1683 & _GEN_1579 : ~_GEN_1643 & _GEN_1579;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1686 = _GEN_36 ? ~_GEN_1685 & _GEN_1580 : ~_GEN_1644 & _GEN_1580;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1688 = _GEN_36 ? ~_GEN_1687 & _GEN_1581 : ~_GEN_1645 & _GEN_1581;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1690 = _GEN_36 ? ~_GEN_1689 & _GEN_1582 : ~_GEN_1646 & _GEN_1582;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1692 = _GEN_36 ? ~_GEN_1691 & _GEN_1583 : ~_GEN_1647 & _GEN_1583;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1694 = _GEN_36 ? ~_GEN_1693 & _GEN_1584 : ~_GEN_1648 & _GEN_1584;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1696 = _GEN_36 ? ~_GEN_1695 & _GEN_1585 : ~_GEN_1649 & _GEN_1585;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1698 = _GEN_36 ? ~_GEN_1697 & _GEN_1586 : ~_GEN_1650 & _GEN_1586;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1700 = _GEN_36 ? ~_GEN_1699 & _GEN_1587 : ~_GEN_1651 & _GEN_1587;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1702 = _GEN_36 ? ~_GEN_1701 & _GEN_1588 : ~_GEN_1652 & _GEN_1588;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1704 = _GEN_36 ? ~_GEN_1703 & _GEN_1589 : ~_GEN_1653 & _GEN_1589;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1706 = _GEN_36 ? ~_GEN_1705 & _GEN_1590 : ~_GEN_1654 & _GEN_1590;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1708 = _GEN_36 ? ~_GEN_1707 & _GEN_1591 : ~_GEN_1655 & _GEN_1591;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1710 = _GEN_36 ? ~_GEN_1709 & _GEN_1592 : ~_GEN_1656 & _GEN_1592;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1712 = _GEN_36 ? ~_GEN_1711 & _GEN_1593 : ~_GEN_1657 & _GEN_1593;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1714 = _GEN_36 ? ~_GEN_1713 & _GEN_1594 : ~_GEN_1658 & _GEN_1594;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1716 = _GEN_36 ? ~_GEN_1715 & _GEN_1595 : ~_GEN_1659 & _GEN_1595;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1718 = _GEN_36 ? ~_GEN_1717 & _GEN_1596 : ~_GEN_1660 & _GEN_1596;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1720 = _GEN_36 ? ~_GEN_1719 & _GEN_1597 : ~_GEN_1661 & _GEN_1597;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1722 = _GEN_36 ? ~_GEN_1721 & _GEN_1598 : ~_GEN_1662 & _GEN_1598;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1724 = _GEN_36 ? ~_GEN_1723 & _GEN_1599 : ~_GEN_1663 & _GEN_1599;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1726 = _GEN_36 ? ~_GEN_1725 & _GEN_1600 : ~_GEN_1664 & _GEN_1600;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1728 = _GEN_36 ? ~_GEN_1727 & _GEN_1601 : ~_GEN_1665 & _GEN_1601;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1730 = _GEN_36 ? ~_GEN_1729 & _GEN_1602 : ~_GEN_1666 & _GEN_1602;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1731 = _GEN_36 ? ~_GEN_1667 & _GEN_1603 : ~_GEN_1635 & _GEN_1603;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1732 = _GEN_36 ? ~_GEN_1669 & _GEN_1604 : ~_GEN_1636 & _GEN_1604;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1733 = _GEN_36 ? ~_GEN_1671 & _GEN_1605 : ~_GEN_1637 & _GEN_1605;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1734 = _GEN_36 ? ~_GEN_1673 & _GEN_1606 : ~_GEN_1638 & _GEN_1606;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1735 = _GEN_36 ? ~_GEN_1675 & _GEN_1607 : ~_GEN_1639 & _GEN_1607;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1736 = _GEN_36 ? ~_GEN_1677 & _GEN_1608 : ~_GEN_1640 & _GEN_1608;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1737 = _GEN_36 ? ~_GEN_1679 & _GEN_1609 : ~_GEN_1641 & _GEN_1609;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1738 = _GEN_36 ? ~_GEN_1681 & _GEN_1610 : ~_GEN_1642 & _GEN_1610;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1739 = _GEN_36 ? ~_GEN_1683 & _GEN_1611 : ~_GEN_1643 & _GEN_1611;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1740 = _GEN_36 ? ~_GEN_1685 & _GEN_1612 : ~_GEN_1644 & _GEN_1612;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1741 = _GEN_36 ? ~_GEN_1687 & _GEN_1613 : ~_GEN_1645 & _GEN_1613;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1742 = _GEN_36 ? ~_GEN_1689 & _GEN_1614 : ~_GEN_1646 & _GEN_1614;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1743 = _GEN_36 ? ~_GEN_1691 & _GEN_1615 : ~_GEN_1647 & _GEN_1615;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1744 = _GEN_36 ? ~_GEN_1693 & _GEN_1616 : ~_GEN_1648 & _GEN_1616;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1745 = _GEN_36 ? ~_GEN_1695 & _GEN_1617 : ~_GEN_1649 & _GEN_1617;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1746 = _GEN_36 ? ~_GEN_1697 & _GEN_1618 : ~_GEN_1650 & _GEN_1618;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1747 = _GEN_36 ? ~_GEN_1699 & _GEN_1619 : ~_GEN_1651 & _GEN_1619;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1748 = _GEN_36 ? ~_GEN_1701 & _GEN_1620 : ~_GEN_1652 & _GEN_1620;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1749 = _GEN_36 ? ~_GEN_1703 & _GEN_1621 : ~_GEN_1653 & _GEN_1621;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1750 = _GEN_36 ? ~_GEN_1705 & _GEN_1622 : ~_GEN_1654 & _GEN_1622;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1751 = _GEN_36 ? ~_GEN_1707 & _GEN_1623 : ~_GEN_1655 & _GEN_1623;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1752 = _GEN_36 ? ~_GEN_1709 & _GEN_1624 : ~_GEN_1656 & _GEN_1624;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1753 = _GEN_36 ? ~_GEN_1711 & _GEN_1625 : ~_GEN_1657 & _GEN_1625;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1754 = _GEN_36 ? ~_GEN_1713 & _GEN_1626 : ~_GEN_1658 & _GEN_1626;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1755 = _GEN_36 ? ~_GEN_1715 & _GEN_1627 : ~_GEN_1659 & _GEN_1627;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1756 = _GEN_36 ? ~_GEN_1717 & _GEN_1628 : ~_GEN_1660 & _GEN_1628;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1757 = _GEN_36 ? ~_GEN_1719 & _GEN_1629 : ~_GEN_1661 & _GEN_1629;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1758 = _GEN_36 ? ~_GEN_1721 & _GEN_1630 : ~_GEN_1662 & _GEN_1630;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1759 = _GEN_36 ? ~_GEN_1723 & _GEN_1631 : ~_GEN_1663 & _GEN_1631;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1760 = _GEN_36 ? ~_GEN_1725 & _GEN_1632 : ~_GEN_1664 & _GEN_1632;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1761 = _GEN_36 ? ~_GEN_1727 & _GEN_1633 : ~_GEN_1665 & _GEN_1633;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1762 = _GEN_36 ? ~_GEN_1729 & _GEN_1634 : ~_GEN_1666 & _GEN_1634;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1796 = _GEN_38 ? ~_GEN_1795 & _GEN_1668 : ~_GEN_1763 & _GEN_1668;	// rob.scala:346:{27,69}, :347:31
    _GEN_1798 = _GEN_38 ? ~_GEN_1797 & _GEN_1670 : ~_GEN_1764 & _GEN_1670;	// rob.scala:346:{27,69}, :347:31
    _GEN_1800 = _GEN_38 ? ~_GEN_1799 & _GEN_1672 : ~_GEN_1765 & _GEN_1672;	// rob.scala:346:{27,69}, :347:31
    _GEN_1802 = _GEN_38 ? ~_GEN_1801 & _GEN_1674 : ~_GEN_1766 & _GEN_1674;	// rob.scala:346:{27,69}, :347:31
    _GEN_1804 = _GEN_38 ? ~_GEN_1803 & _GEN_1676 : ~_GEN_1767 & _GEN_1676;	// rob.scala:346:{27,69}, :347:31
    _GEN_1806 = _GEN_38 ? ~_GEN_1805 & _GEN_1678 : ~_GEN_1768 & _GEN_1678;	// rob.scala:346:{27,69}, :347:31
    _GEN_1808 = _GEN_38 ? ~_GEN_1807 & _GEN_1680 : ~_GEN_1769 & _GEN_1680;	// rob.scala:346:{27,69}, :347:31
    _GEN_1810 = _GEN_38 ? ~_GEN_1809 & _GEN_1682 : ~_GEN_1770 & _GEN_1682;	// rob.scala:346:{27,69}, :347:31
    _GEN_1812 = _GEN_38 ? ~_GEN_1811 & _GEN_1684 : ~_GEN_1771 & _GEN_1684;	// rob.scala:346:{27,69}, :347:31
    _GEN_1814 = _GEN_38 ? ~_GEN_1813 & _GEN_1686 : ~_GEN_1772 & _GEN_1686;	// rob.scala:346:{27,69}, :347:31
    _GEN_1816 = _GEN_38 ? ~_GEN_1815 & _GEN_1688 : ~_GEN_1773 & _GEN_1688;	// rob.scala:346:{27,69}, :347:31
    _GEN_1818 = _GEN_38 ? ~_GEN_1817 & _GEN_1690 : ~_GEN_1774 & _GEN_1690;	// rob.scala:346:{27,69}, :347:31
    _GEN_1820 = _GEN_38 ? ~_GEN_1819 & _GEN_1692 : ~_GEN_1775 & _GEN_1692;	// rob.scala:346:{27,69}, :347:31
    _GEN_1822 = _GEN_38 ? ~_GEN_1821 & _GEN_1694 : ~_GEN_1776 & _GEN_1694;	// rob.scala:346:{27,69}, :347:31
    _GEN_1824 = _GEN_38 ? ~_GEN_1823 & _GEN_1696 : ~_GEN_1777 & _GEN_1696;	// rob.scala:346:{27,69}, :347:31
    _GEN_1826 = _GEN_38 ? ~_GEN_1825 & _GEN_1698 : ~_GEN_1778 & _GEN_1698;	// rob.scala:346:{27,69}, :347:31
    _GEN_1828 = _GEN_38 ? ~_GEN_1827 & _GEN_1700 : ~_GEN_1779 & _GEN_1700;	// rob.scala:346:{27,69}, :347:31
    _GEN_1830 = _GEN_38 ? ~_GEN_1829 & _GEN_1702 : ~_GEN_1780 & _GEN_1702;	// rob.scala:346:{27,69}, :347:31
    _GEN_1832 = _GEN_38 ? ~_GEN_1831 & _GEN_1704 : ~_GEN_1781 & _GEN_1704;	// rob.scala:346:{27,69}, :347:31
    _GEN_1834 = _GEN_38 ? ~_GEN_1833 & _GEN_1706 : ~_GEN_1782 & _GEN_1706;	// rob.scala:346:{27,69}, :347:31
    _GEN_1836 = _GEN_38 ? ~_GEN_1835 & _GEN_1708 : ~_GEN_1783 & _GEN_1708;	// rob.scala:346:{27,69}, :347:31
    _GEN_1838 = _GEN_38 ? ~_GEN_1837 & _GEN_1710 : ~_GEN_1784 & _GEN_1710;	// rob.scala:346:{27,69}, :347:31
    _GEN_1840 = _GEN_38 ? ~_GEN_1839 & _GEN_1712 : ~_GEN_1785 & _GEN_1712;	// rob.scala:346:{27,69}, :347:31
    _GEN_1842 = _GEN_38 ? ~_GEN_1841 & _GEN_1714 : ~_GEN_1786 & _GEN_1714;	// rob.scala:346:{27,69}, :347:31
    _GEN_1844 = _GEN_38 ? ~_GEN_1843 & _GEN_1716 : ~_GEN_1787 & _GEN_1716;	// rob.scala:346:{27,69}, :347:31
    _GEN_1846 = _GEN_38 ? ~_GEN_1845 & _GEN_1718 : ~_GEN_1788 & _GEN_1718;	// rob.scala:346:{27,69}, :347:31
    _GEN_1848 = _GEN_38 ? ~_GEN_1847 & _GEN_1720 : ~_GEN_1789 & _GEN_1720;	// rob.scala:346:{27,69}, :347:31
    _GEN_1850 = _GEN_38 ? ~_GEN_1849 & _GEN_1722 : ~_GEN_1790 & _GEN_1722;	// rob.scala:346:{27,69}, :347:31
    _GEN_1852 = _GEN_38 ? ~_GEN_1851 & _GEN_1724 : ~_GEN_1791 & _GEN_1724;	// rob.scala:346:{27,69}, :347:31
    _GEN_1854 = _GEN_38 ? ~_GEN_1853 & _GEN_1726 : ~_GEN_1792 & _GEN_1726;	// rob.scala:346:{27,69}, :347:31
    _GEN_1856 = _GEN_38 ? ~_GEN_1855 & _GEN_1728 : ~_GEN_1793 & _GEN_1728;	// rob.scala:346:{27,69}, :347:31
    _GEN_1858 = _GEN_38 ? ~_GEN_1857 & _GEN_1730 : ~_GEN_1794 & _GEN_1730;	// rob.scala:346:{27,69}, :347:31
    _GEN_1859 = _GEN_38 ? ~_GEN_1795 & _GEN_1731 : ~_GEN_1763 & _GEN_1731;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1860 = _GEN_38 ? ~_GEN_1797 & _GEN_1732 : ~_GEN_1764 & _GEN_1732;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1861 = _GEN_38 ? ~_GEN_1799 & _GEN_1733 : ~_GEN_1765 & _GEN_1733;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1862 = _GEN_38 ? ~_GEN_1801 & _GEN_1734 : ~_GEN_1766 & _GEN_1734;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1863 = _GEN_38 ? ~_GEN_1803 & _GEN_1735 : ~_GEN_1767 & _GEN_1735;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1864 = _GEN_38 ? ~_GEN_1805 & _GEN_1736 : ~_GEN_1768 & _GEN_1736;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1865 = _GEN_38 ? ~_GEN_1807 & _GEN_1737 : ~_GEN_1769 & _GEN_1737;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1866 = _GEN_38 ? ~_GEN_1809 & _GEN_1738 : ~_GEN_1770 & _GEN_1738;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1867 = _GEN_38 ? ~_GEN_1811 & _GEN_1739 : ~_GEN_1771 & _GEN_1739;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1868 = _GEN_38 ? ~_GEN_1813 & _GEN_1740 : ~_GEN_1772 & _GEN_1740;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1869 = _GEN_38 ? ~_GEN_1815 & _GEN_1741 : ~_GEN_1773 & _GEN_1741;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1870 = _GEN_38 ? ~_GEN_1817 & _GEN_1742 : ~_GEN_1774 & _GEN_1742;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1871 = _GEN_38 ? ~_GEN_1819 & _GEN_1743 : ~_GEN_1775 & _GEN_1743;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1872 = _GEN_38 ? ~_GEN_1821 & _GEN_1744 : ~_GEN_1776 & _GEN_1744;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1873 = _GEN_38 ? ~_GEN_1823 & _GEN_1745 : ~_GEN_1777 & _GEN_1745;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1874 = _GEN_38 ? ~_GEN_1825 & _GEN_1746 : ~_GEN_1778 & _GEN_1746;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1875 = _GEN_38 ? ~_GEN_1827 & _GEN_1747 : ~_GEN_1779 & _GEN_1747;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1876 = _GEN_38 ? ~_GEN_1829 & _GEN_1748 : ~_GEN_1780 & _GEN_1748;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1877 = _GEN_38 ? ~_GEN_1831 & _GEN_1749 : ~_GEN_1781 & _GEN_1749;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1878 = _GEN_38 ? ~_GEN_1833 & _GEN_1750 : ~_GEN_1782 & _GEN_1750;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1879 = _GEN_38 ? ~_GEN_1835 & _GEN_1751 : ~_GEN_1783 & _GEN_1751;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1880 = _GEN_38 ? ~_GEN_1837 & _GEN_1752 : ~_GEN_1784 & _GEN_1752;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1881 = _GEN_38 ? ~_GEN_1839 & _GEN_1753 : ~_GEN_1785 & _GEN_1753;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1882 = _GEN_38 ? ~_GEN_1841 & _GEN_1754 : ~_GEN_1786 & _GEN_1754;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1883 = _GEN_38 ? ~_GEN_1843 & _GEN_1755 : ~_GEN_1787 & _GEN_1755;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1884 = _GEN_38 ? ~_GEN_1845 & _GEN_1756 : ~_GEN_1788 & _GEN_1756;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1885 = _GEN_38 ? ~_GEN_1847 & _GEN_1757 : ~_GEN_1789 & _GEN_1757;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1886 = _GEN_38 ? ~_GEN_1849 & _GEN_1758 : ~_GEN_1790 & _GEN_1758;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1887 = _GEN_38 ? ~_GEN_1851 & _GEN_1759 : ~_GEN_1791 & _GEN_1759;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1888 = _GEN_38 ? ~_GEN_1853 & _GEN_1760 : ~_GEN_1792 & _GEN_1760;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1889 = _GEN_38 ? ~_GEN_1855 & _GEN_1761 : ~_GEN_1793 & _GEN_1761;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1890 = _GEN_38 ? ~_GEN_1857 & _GEN_1762 : ~_GEN_1794 & _GEN_1762;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1924 = _GEN_40 ? ~_GEN_1923 & _GEN_1796 : ~_GEN_1891 & _GEN_1796;	// rob.scala:346:{27,69}, :347:31
    _GEN_1926 = _GEN_40 ? ~_GEN_1925 & _GEN_1798 : ~_GEN_1892 & _GEN_1798;	// rob.scala:346:{27,69}, :347:31
    _GEN_1928 = _GEN_40 ? ~_GEN_1927 & _GEN_1800 : ~_GEN_1893 & _GEN_1800;	// rob.scala:346:{27,69}, :347:31
    _GEN_1930 = _GEN_40 ? ~_GEN_1929 & _GEN_1802 : ~_GEN_1894 & _GEN_1802;	// rob.scala:346:{27,69}, :347:31
    _GEN_1932 = _GEN_40 ? ~_GEN_1931 & _GEN_1804 : ~_GEN_1895 & _GEN_1804;	// rob.scala:346:{27,69}, :347:31
    _GEN_1934 = _GEN_40 ? ~_GEN_1933 & _GEN_1806 : ~_GEN_1896 & _GEN_1806;	// rob.scala:346:{27,69}, :347:31
    _GEN_1936 = _GEN_40 ? ~_GEN_1935 & _GEN_1808 : ~_GEN_1897 & _GEN_1808;	// rob.scala:346:{27,69}, :347:31
    _GEN_1938 = _GEN_40 ? ~_GEN_1937 & _GEN_1810 : ~_GEN_1898 & _GEN_1810;	// rob.scala:346:{27,69}, :347:31
    _GEN_1940 = _GEN_40 ? ~_GEN_1939 & _GEN_1812 : ~_GEN_1899 & _GEN_1812;	// rob.scala:346:{27,69}, :347:31
    _GEN_1942 = _GEN_40 ? ~_GEN_1941 & _GEN_1814 : ~_GEN_1900 & _GEN_1814;	// rob.scala:346:{27,69}, :347:31
    _GEN_1944 = _GEN_40 ? ~_GEN_1943 & _GEN_1816 : ~_GEN_1901 & _GEN_1816;	// rob.scala:346:{27,69}, :347:31
    _GEN_1946 = _GEN_40 ? ~_GEN_1945 & _GEN_1818 : ~_GEN_1902 & _GEN_1818;	// rob.scala:346:{27,69}, :347:31
    _GEN_1948 = _GEN_40 ? ~_GEN_1947 & _GEN_1820 : ~_GEN_1903 & _GEN_1820;	// rob.scala:346:{27,69}, :347:31
    _GEN_1950 = _GEN_40 ? ~_GEN_1949 & _GEN_1822 : ~_GEN_1904 & _GEN_1822;	// rob.scala:346:{27,69}, :347:31
    _GEN_1952 = _GEN_40 ? ~_GEN_1951 & _GEN_1824 : ~_GEN_1905 & _GEN_1824;	// rob.scala:346:{27,69}, :347:31
    _GEN_1954 = _GEN_40 ? ~_GEN_1953 & _GEN_1826 : ~_GEN_1906 & _GEN_1826;	// rob.scala:346:{27,69}, :347:31
    _GEN_1956 = _GEN_40 ? ~_GEN_1955 & _GEN_1828 : ~_GEN_1907 & _GEN_1828;	// rob.scala:346:{27,69}, :347:31
    _GEN_1958 = _GEN_40 ? ~_GEN_1957 & _GEN_1830 : ~_GEN_1908 & _GEN_1830;	// rob.scala:346:{27,69}, :347:31
    _GEN_1960 = _GEN_40 ? ~_GEN_1959 & _GEN_1832 : ~_GEN_1909 & _GEN_1832;	// rob.scala:346:{27,69}, :347:31
    _GEN_1962 = _GEN_40 ? ~_GEN_1961 & _GEN_1834 : ~_GEN_1910 & _GEN_1834;	// rob.scala:346:{27,69}, :347:31
    _GEN_1964 = _GEN_40 ? ~_GEN_1963 & _GEN_1836 : ~_GEN_1911 & _GEN_1836;	// rob.scala:346:{27,69}, :347:31
    _GEN_1966 = _GEN_40 ? ~_GEN_1965 & _GEN_1838 : ~_GEN_1912 & _GEN_1838;	// rob.scala:346:{27,69}, :347:31
    _GEN_1968 = _GEN_40 ? ~_GEN_1967 & _GEN_1840 : ~_GEN_1913 & _GEN_1840;	// rob.scala:346:{27,69}, :347:31
    _GEN_1970 = _GEN_40 ? ~_GEN_1969 & _GEN_1842 : ~_GEN_1914 & _GEN_1842;	// rob.scala:346:{27,69}, :347:31
    _GEN_1972 = _GEN_40 ? ~_GEN_1971 & _GEN_1844 : ~_GEN_1915 & _GEN_1844;	// rob.scala:346:{27,69}, :347:31
    _GEN_1974 = _GEN_40 ? ~_GEN_1973 & _GEN_1846 : ~_GEN_1916 & _GEN_1846;	// rob.scala:346:{27,69}, :347:31
    _GEN_1976 = _GEN_40 ? ~_GEN_1975 & _GEN_1848 : ~_GEN_1917 & _GEN_1848;	// rob.scala:346:{27,69}, :347:31
    _GEN_1978 = _GEN_40 ? ~_GEN_1977 & _GEN_1850 : ~_GEN_1918 & _GEN_1850;	// rob.scala:346:{27,69}, :347:31
    _GEN_1980 = _GEN_40 ? ~_GEN_1979 & _GEN_1852 : ~_GEN_1919 & _GEN_1852;	// rob.scala:346:{27,69}, :347:31
    _GEN_1982 = _GEN_40 ? ~_GEN_1981 & _GEN_1854 : ~_GEN_1920 & _GEN_1854;	// rob.scala:346:{27,69}, :347:31
    _GEN_1984 = _GEN_40 ? ~_GEN_1983 & _GEN_1856 : ~_GEN_1921 & _GEN_1856;	// rob.scala:346:{27,69}, :347:31
    _GEN_1986 = _GEN_40 ? ~_GEN_1985 & _GEN_1858 : ~_GEN_1922 & _GEN_1858;	// rob.scala:346:{27,69}, :347:31
    _GEN_1987 = _GEN_40 ? ~_GEN_1923 & _GEN_1859 : ~_GEN_1891 & _GEN_1859;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1988 = _GEN_40 ? ~_GEN_1925 & _GEN_1860 : ~_GEN_1892 & _GEN_1860;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1989 = _GEN_40 ? ~_GEN_1927 & _GEN_1861 : ~_GEN_1893 & _GEN_1861;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1990 = _GEN_40 ? ~_GEN_1929 & _GEN_1862 : ~_GEN_1894 & _GEN_1862;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1991 = _GEN_40 ? ~_GEN_1931 & _GEN_1863 : ~_GEN_1895 & _GEN_1863;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1992 = _GEN_40 ? ~_GEN_1933 & _GEN_1864 : ~_GEN_1896 & _GEN_1864;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1993 = _GEN_40 ? ~_GEN_1935 & _GEN_1865 : ~_GEN_1897 & _GEN_1865;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1994 = _GEN_40 ? ~_GEN_1937 & _GEN_1866 : ~_GEN_1898 & _GEN_1866;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1995 = _GEN_40 ? ~_GEN_1939 & _GEN_1867 : ~_GEN_1899 & _GEN_1867;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1996 = _GEN_40 ? ~_GEN_1941 & _GEN_1868 : ~_GEN_1900 & _GEN_1868;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1997 = _GEN_40 ? ~_GEN_1943 & _GEN_1869 : ~_GEN_1901 & _GEN_1869;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1998 = _GEN_40 ? ~_GEN_1945 & _GEN_1870 : ~_GEN_1902 & _GEN_1870;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1999 = _GEN_40 ? ~_GEN_1947 & _GEN_1871 : ~_GEN_1903 & _GEN_1871;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2000 = _GEN_40 ? ~_GEN_1949 & _GEN_1872 : ~_GEN_1904 & _GEN_1872;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2001 = _GEN_40 ? ~_GEN_1951 & _GEN_1873 : ~_GEN_1905 & _GEN_1873;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2002 = _GEN_40 ? ~_GEN_1953 & _GEN_1874 : ~_GEN_1906 & _GEN_1874;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2003 = _GEN_40 ? ~_GEN_1955 & _GEN_1875 : ~_GEN_1907 & _GEN_1875;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2004 = _GEN_40 ? ~_GEN_1957 & _GEN_1876 : ~_GEN_1908 & _GEN_1876;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2005 = _GEN_40 ? ~_GEN_1959 & _GEN_1877 : ~_GEN_1909 & _GEN_1877;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2006 = _GEN_40 ? ~_GEN_1961 & _GEN_1878 : ~_GEN_1910 & _GEN_1878;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2007 = _GEN_40 ? ~_GEN_1963 & _GEN_1879 : ~_GEN_1911 & _GEN_1879;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2008 = _GEN_40 ? ~_GEN_1965 & _GEN_1880 : ~_GEN_1912 & _GEN_1880;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2009 = _GEN_40 ? ~_GEN_1967 & _GEN_1881 : ~_GEN_1913 & _GEN_1881;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2010 = _GEN_40 ? ~_GEN_1969 & _GEN_1882 : ~_GEN_1914 & _GEN_1882;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2011 = _GEN_40 ? ~_GEN_1971 & _GEN_1883 : ~_GEN_1915 & _GEN_1883;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2012 = _GEN_40 ? ~_GEN_1973 & _GEN_1884 : ~_GEN_1916 & _GEN_1884;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2013 = _GEN_40 ? ~_GEN_1975 & _GEN_1885 : ~_GEN_1917 & _GEN_1885;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2014 = _GEN_40 ? ~_GEN_1977 & _GEN_1886 : ~_GEN_1918 & _GEN_1886;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2015 = _GEN_40 ? ~_GEN_1979 & _GEN_1887 : ~_GEN_1919 & _GEN_1887;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2016 = _GEN_40 ? ~_GEN_1981 & _GEN_1888 : ~_GEN_1920 & _GEN_1888;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2017 = _GEN_40 ? ~_GEN_1983 & _GEN_1889 : ~_GEN_1921 & _GEN_1889;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2018 = _GEN_40 ? ~_GEN_1985 & _GEN_1890 : ~_GEN_1922 & _GEN_1890;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2052 = _GEN_42 ? ~_GEN_2051 & _GEN_1924 : ~_GEN_2019 & _GEN_1924;	// rob.scala:346:{27,69}, :347:31
    _GEN_2054 = _GEN_42 ? ~_GEN_2053 & _GEN_1926 : ~_GEN_2020 & _GEN_1926;	// rob.scala:346:{27,69}, :347:31
    _GEN_2056 = _GEN_42 ? ~_GEN_2055 & _GEN_1928 : ~_GEN_2021 & _GEN_1928;	// rob.scala:346:{27,69}, :347:31
    _GEN_2058 = _GEN_42 ? ~_GEN_2057 & _GEN_1930 : ~_GEN_2022 & _GEN_1930;	// rob.scala:346:{27,69}, :347:31
    _GEN_2060 = _GEN_42 ? ~_GEN_2059 & _GEN_1932 : ~_GEN_2023 & _GEN_1932;	// rob.scala:346:{27,69}, :347:31
    _GEN_2062 = _GEN_42 ? ~_GEN_2061 & _GEN_1934 : ~_GEN_2024 & _GEN_1934;	// rob.scala:346:{27,69}, :347:31
    _GEN_2064 = _GEN_42 ? ~_GEN_2063 & _GEN_1936 : ~_GEN_2025 & _GEN_1936;	// rob.scala:346:{27,69}, :347:31
    _GEN_2066 = _GEN_42 ? ~_GEN_2065 & _GEN_1938 : ~_GEN_2026 & _GEN_1938;	// rob.scala:346:{27,69}, :347:31
    _GEN_2068 = _GEN_42 ? ~_GEN_2067 & _GEN_1940 : ~_GEN_2027 & _GEN_1940;	// rob.scala:346:{27,69}, :347:31
    _GEN_2070 = _GEN_42 ? ~_GEN_2069 & _GEN_1942 : ~_GEN_2028 & _GEN_1942;	// rob.scala:346:{27,69}, :347:31
    _GEN_2072 = _GEN_42 ? ~_GEN_2071 & _GEN_1944 : ~_GEN_2029 & _GEN_1944;	// rob.scala:346:{27,69}, :347:31
    _GEN_2074 = _GEN_42 ? ~_GEN_2073 & _GEN_1946 : ~_GEN_2030 & _GEN_1946;	// rob.scala:346:{27,69}, :347:31
    _GEN_2076 = _GEN_42 ? ~_GEN_2075 & _GEN_1948 : ~_GEN_2031 & _GEN_1948;	// rob.scala:346:{27,69}, :347:31
    _GEN_2078 = _GEN_42 ? ~_GEN_2077 & _GEN_1950 : ~_GEN_2032 & _GEN_1950;	// rob.scala:346:{27,69}, :347:31
    _GEN_2080 = _GEN_42 ? ~_GEN_2079 & _GEN_1952 : ~_GEN_2033 & _GEN_1952;	// rob.scala:346:{27,69}, :347:31
    _GEN_2082 = _GEN_42 ? ~_GEN_2081 & _GEN_1954 : ~_GEN_2034 & _GEN_1954;	// rob.scala:346:{27,69}, :347:31
    _GEN_2084 = _GEN_42 ? ~_GEN_2083 & _GEN_1956 : ~_GEN_2035 & _GEN_1956;	// rob.scala:346:{27,69}, :347:31
    _GEN_2086 = _GEN_42 ? ~_GEN_2085 & _GEN_1958 : ~_GEN_2036 & _GEN_1958;	// rob.scala:346:{27,69}, :347:31
    _GEN_2088 = _GEN_42 ? ~_GEN_2087 & _GEN_1960 : ~_GEN_2037 & _GEN_1960;	// rob.scala:346:{27,69}, :347:31
    _GEN_2090 = _GEN_42 ? ~_GEN_2089 & _GEN_1962 : ~_GEN_2038 & _GEN_1962;	// rob.scala:346:{27,69}, :347:31
    _GEN_2092 = _GEN_42 ? ~_GEN_2091 & _GEN_1964 : ~_GEN_2039 & _GEN_1964;	// rob.scala:346:{27,69}, :347:31
    _GEN_2094 = _GEN_42 ? ~_GEN_2093 & _GEN_1966 : ~_GEN_2040 & _GEN_1966;	// rob.scala:346:{27,69}, :347:31
    _GEN_2096 = _GEN_42 ? ~_GEN_2095 & _GEN_1968 : ~_GEN_2041 & _GEN_1968;	// rob.scala:346:{27,69}, :347:31
    _GEN_2098 = _GEN_42 ? ~_GEN_2097 & _GEN_1970 : ~_GEN_2042 & _GEN_1970;	// rob.scala:346:{27,69}, :347:31
    _GEN_2100 = _GEN_42 ? ~_GEN_2099 & _GEN_1972 : ~_GEN_2043 & _GEN_1972;	// rob.scala:346:{27,69}, :347:31
    _GEN_2102 = _GEN_42 ? ~_GEN_2101 & _GEN_1974 : ~_GEN_2044 & _GEN_1974;	// rob.scala:346:{27,69}, :347:31
    _GEN_2104 = _GEN_42 ? ~_GEN_2103 & _GEN_1976 : ~_GEN_2045 & _GEN_1976;	// rob.scala:346:{27,69}, :347:31
    _GEN_2106 = _GEN_42 ? ~_GEN_2105 & _GEN_1978 : ~_GEN_2046 & _GEN_1978;	// rob.scala:346:{27,69}, :347:31
    _GEN_2108 = _GEN_42 ? ~_GEN_2107 & _GEN_1980 : ~_GEN_2047 & _GEN_1980;	// rob.scala:346:{27,69}, :347:31
    _GEN_2110 = _GEN_42 ? ~_GEN_2109 & _GEN_1982 : ~_GEN_2048 & _GEN_1982;	// rob.scala:346:{27,69}, :347:31
    _GEN_2112 = _GEN_42 ? ~_GEN_2111 & _GEN_1984 : ~_GEN_2049 & _GEN_1984;	// rob.scala:346:{27,69}, :347:31
    _GEN_2114 = _GEN_42 ? ~_GEN_2113 & _GEN_1986 : ~_GEN_2050 & _GEN_1986;	// rob.scala:346:{27,69}, :347:31
    _GEN_2115 = _GEN_42 ? ~_GEN_2051 & _GEN_1987 : ~_GEN_2019 & _GEN_1987;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2116 = _GEN_42 ? ~_GEN_2053 & _GEN_1988 : ~_GEN_2020 & _GEN_1988;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2117 = _GEN_42 ? ~_GEN_2055 & _GEN_1989 : ~_GEN_2021 & _GEN_1989;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2118 = _GEN_42 ? ~_GEN_2057 & _GEN_1990 : ~_GEN_2022 & _GEN_1990;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2119 = _GEN_42 ? ~_GEN_2059 & _GEN_1991 : ~_GEN_2023 & _GEN_1991;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2120 = _GEN_42 ? ~_GEN_2061 & _GEN_1992 : ~_GEN_2024 & _GEN_1992;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2121 = _GEN_42 ? ~_GEN_2063 & _GEN_1993 : ~_GEN_2025 & _GEN_1993;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2122 = _GEN_42 ? ~_GEN_2065 & _GEN_1994 : ~_GEN_2026 & _GEN_1994;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2123 = _GEN_42 ? ~_GEN_2067 & _GEN_1995 : ~_GEN_2027 & _GEN_1995;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2124 = _GEN_42 ? ~_GEN_2069 & _GEN_1996 : ~_GEN_2028 & _GEN_1996;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2125 = _GEN_42 ? ~_GEN_2071 & _GEN_1997 : ~_GEN_2029 & _GEN_1997;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2126 = _GEN_42 ? ~_GEN_2073 & _GEN_1998 : ~_GEN_2030 & _GEN_1998;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2127 = _GEN_42 ? ~_GEN_2075 & _GEN_1999 : ~_GEN_2031 & _GEN_1999;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2128 = _GEN_42 ? ~_GEN_2077 & _GEN_2000 : ~_GEN_2032 & _GEN_2000;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2129 = _GEN_42 ? ~_GEN_2079 & _GEN_2001 : ~_GEN_2033 & _GEN_2001;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2130 = _GEN_42 ? ~_GEN_2081 & _GEN_2002 : ~_GEN_2034 & _GEN_2002;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2131 = _GEN_42 ? ~_GEN_2083 & _GEN_2003 : ~_GEN_2035 & _GEN_2003;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2132 = _GEN_42 ? ~_GEN_2085 & _GEN_2004 : ~_GEN_2036 & _GEN_2004;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2133 = _GEN_42 ? ~_GEN_2087 & _GEN_2005 : ~_GEN_2037 & _GEN_2005;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2134 = _GEN_42 ? ~_GEN_2089 & _GEN_2006 : ~_GEN_2038 & _GEN_2006;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2135 = _GEN_42 ? ~_GEN_2091 & _GEN_2007 : ~_GEN_2039 & _GEN_2007;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2136 = _GEN_42 ? ~_GEN_2093 & _GEN_2008 : ~_GEN_2040 & _GEN_2008;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2137 = _GEN_42 ? ~_GEN_2095 & _GEN_2009 : ~_GEN_2041 & _GEN_2009;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2138 = _GEN_42 ? ~_GEN_2097 & _GEN_2010 : ~_GEN_2042 & _GEN_2010;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2139 = _GEN_42 ? ~_GEN_2099 & _GEN_2011 : ~_GEN_2043 & _GEN_2011;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2140 = _GEN_42 ? ~_GEN_2101 & _GEN_2012 : ~_GEN_2044 & _GEN_2012;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2141 = _GEN_42 ? ~_GEN_2103 & _GEN_2013 : ~_GEN_2045 & _GEN_2013;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2142 = _GEN_42 ? ~_GEN_2105 & _GEN_2014 : ~_GEN_2046 & _GEN_2014;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2143 = _GEN_42 ? ~_GEN_2107 & _GEN_2015 : ~_GEN_2047 & _GEN_2015;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2144 = _GEN_42 ? ~_GEN_2109 & _GEN_2016 : ~_GEN_2048 & _GEN_2016;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2145 = _GEN_42 ? ~_GEN_2111 & _GEN_2017 : ~_GEN_2049 & _GEN_2017;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2146 = _GEN_42 ? ~_GEN_2113 & _GEN_2018 : ~_GEN_2050 & _GEN_2018;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2180 = _GEN_44 ? ~_GEN_2179 & _GEN_2052 : ~_GEN_2147 & _GEN_2052;	// rob.scala:346:{27,69}, :347:31
    _GEN_2182 = _GEN_44 ? ~_GEN_2181 & _GEN_2054 : ~_GEN_2148 & _GEN_2054;	// rob.scala:346:{27,69}, :347:31
    _GEN_2184 = _GEN_44 ? ~_GEN_2183 & _GEN_2056 : ~_GEN_2149 & _GEN_2056;	// rob.scala:346:{27,69}, :347:31
    _GEN_2186 = _GEN_44 ? ~_GEN_2185 & _GEN_2058 : ~_GEN_2150 & _GEN_2058;	// rob.scala:346:{27,69}, :347:31
    _GEN_2188 = _GEN_44 ? ~_GEN_2187 & _GEN_2060 : ~_GEN_2151 & _GEN_2060;	// rob.scala:346:{27,69}, :347:31
    _GEN_2190 = _GEN_44 ? ~_GEN_2189 & _GEN_2062 : ~_GEN_2152 & _GEN_2062;	// rob.scala:346:{27,69}, :347:31
    _GEN_2192 = _GEN_44 ? ~_GEN_2191 & _GEN_2064 : ~_GEN_2153 & _GEN_2064;	// rob.scala:346:{27,69}, :347:31
    _GEN_2194 = _GEN_44 ? ~_GEN_2193 & _GEN_2066 : ~_GEN_2154 & _GEN_2066;	// rob.scala:346:{27,69}, :347:31
    _GEN_2196 = _GEN_44 ? ~_GEN_2195 & _GEN_2068 : ~_GEN_2155 & _GEN_2068;	// rob.scala:346:{27,69}, :347:31
    _GEN_2198 = _GEN_44 ? ~_GEN_2197 & _GEN_2070 : ~_GEN_2156 & _GEN_2070;	// rob.scala:346:{27,69}, :347:31
    _GEN_2200 = _GEN_44 ? ~_GEN_2199 & _GEN_2072 : ~_GEN_2157 & _GEN_2072;	// rob.scala:346:{27,69}, :347:31
    _GEN_2202 = _GEN_44 ? ~_GEN_2201 & _GEN_2074 : ~_GEN_2158 & _GEN_2074;	// rob.scala:346:{27,69}, :347:31
    _GEN_2204 = _GEN_44 ? ~_GEN_2203 & _GEN_2076 : ~_GEN_2159 & _GEN_2076;	// rob.scala:346:{27,69}, :347:31
    _GEN_2206 = _GEN_44 ? ~_GEN_2205 & _GEN_2078 : ~_GEN_2160 & _GEN_2078;	// rob.scala:346:{27,69}, :347:31
    _GEN_2208 = _GEN_44 ? ~_GEN_2207 & _GEN_2080 : ~_GEN_2161 & _GEN_2080;	// rob.scala:346:{27,69}, :347:31
    _GEN_2210 = _GEN_44 ? ~_GEN_2209 & _GEN_2082 : ~_GEN_2162 & _GEN_2082;	// rob.scala:346:{27,69}, :347:31
    _GEN_2212 = _GEN_44 ? ~_GEN_2211 & _GEN_2084 : ~_GEN_2163 & _GEN_2084;	// rob.scala:346:{27,69}, :347:31
    _GEN_2214 = _GEN_44 ? ~_GEN_2213 & _GEN_2086 : ~_GEN_2164 & _GEN_2086;	// rob.scala:346:{27,69}, :347:31
    _GEN_2216 = _GEN_44 ? ~_GEN_2215 & _GEN_2088 : ~_GEN_2165 & _GEN_2088;	// rob.scala:346:{27,69}, :347:31
    _GEN_2218 = _GEN_44 ? ~_GEN_2217 & _GEN_2090 : ~_GEN_2166 & _GEN_2090;	// rob.scala:346:{27,69}, :347:31
    _GEN_2220 = _GEN_44 ? ~_GEN_2219 & _GEN_2092 : ~_GEN_2167 & _GEN_2092;	// rob.scala:346:{27,69}, :347:31
    _GEN_2222 = _GEN_44 ? ~_GEN_2221 & _GEN_2094 : ~_GEN_2168 & _GEN_2094;	// rob.scala:346:{27,69}, :347:31
    _GEN_2224 = _GEN_44 ? ~_GEN_2223 & _GEN_2096 : ~_GEN_2169 & _GEN_2096;	// rob.scala:346:{27,69}, :347:31
    _GEN_2226 = _GEN_44 ? ~_GEN_2225 & _GEN_2098 : ~_GEN_2170 & _GEN_2098;	// rob.scala:346:{27,69}, :347:31
    _GEN_2228 = _GEN_44 ? ~_GEN_2227 & _GEN_2100 : ~_GEN_2171 & _GEN_2100;	// rob.scala:346:{27,69}, :347:31
    _GEN_2230 = _GEN_44 ? ~_GEN_2229 & _GEN_2102 : ~_GEN_2172 & _GEN_2102;	// rob.scala:346:{27,69}, :347:31
    _GEN_2232 = _GEN_44 ? ~_GEN_2231 & _GEN_2104 : ~_GEN_2173 & _GEN_2104;	// rob.scala:346:{27,69}, :347:31
    _GEN_2234 = _GEN_44 ? ~_GEN_2233 & _GEN_2106 : ~_GEN_2174 & _GEN_2106;	// rob.scala:346:{27,69}, :347:31
    _GEN_2236 = _GEN_44 ? ~_GEN_2235 & _GEN_2108 : ~_GEN_2175 & _GEN_2108;	// rob.scala:346:{27,69}, :347:31
    _GEN_2238 = _GEN_44 ? ~_GEN_2237 & _GEN_2110 : ~_GEN_2176 & _GEN_2110;	// rob.scala:346:{27,69}, :347:31
    _GEN_2240 = _GEN_44 ? ~_GEN_2239 & _GEN_2112 : ~_GEN_2177 & _GEN_2112;	// rob.scala:346:{27,69}, :347:31
    _GEN_2242 = _GEN_44 ? ~_GEN_2241 & _GEN_2114 : ~_GEN_2178 & _GEN_2114;	// rob.scala:346:{27,69}, :347:31
    _GEN_2243 = _GEN_44 ? ~_GEN_2179 & _GEN_2115 : ~_GEN_2147 & _GEN_2115;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2244 = _GEN_44 ? ~_GEN_2181 & _GEN_2116 : ~_GEN_2148 & _GEN_2116;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2245 = _GEN_44 ? ~_GEN_2183 & _GEN_2117 : ~_GEN_2149 & _GEN_2117;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2246 = _GEN_44 ? ~_GEN_2185 & _GEN_2118 : ~_GEN_2150 & _GEN_2118;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2247 = _GEN_44 ? ~_GEN_2187 & _GEN_2119 : ~_GEN_2151 & _GEN_2119;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2248 = _GEN_44 ? ~_GEN_2189 & _GEN_2120 : ~_GEN_2152 & _GEN_2120;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2249 = _GEN_44 ? ~_GEN_2191 & _GEN_2121 : ~_GEN_2153 & _GEN_2121;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2250 = _GEN_44 ? ~_GEN_2193 & _GEN_2122 : ~_GEN_2154 & _GEN_2122;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2251 = _GEN_44 ? ~_GEN_2195 & _GEN_2123 : ~_GEN_2155 & _GEN_2123;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2252 = _GEN_44 ? ~_GEN_2197 & _GEN_2124 : ~_GEN_2156 & _GEN_2124;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2253 = _GEN_44 ? ~_GEN_2199 & _GEN_2125 : ~_GEN_2157 & _GEN_2125;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2254 = _GEN_44 ? ~_GEN_2201 & _GEN_2126 : ~_GEN_2158 & _GEN_2126;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2255 = _GEN_44 ? ~_GEN_2203 & _GEN_2127 : ~_GEN_2159 & _GEN_2127;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2256 = _GEN_44 ? ~_GEN_2205 & _GEN_2128 : ~_GEN_2160 & _GEN_2128;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2257 = _GEN_44 ? ~_GEN_2207 & _GEN_2129 : ~_GEN_2161 & _GEN_2129;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2258 = _GEN_44 ? ~_GEN_2209 & _GEN_2130 : ~_GEN_2162 & _GEN_2130;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2259 = _GEN_44 ? ~_GEN_2211 & _GEN_2131 : ~_GEN_2163 & _GEN_2131;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2260 = _GEN_44 ? ~_GEN_2213 & _GEN_2132 : ~_GEN_2164 & _GEN_2132;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2261 = _GEN_44 ? ~_GEN_2215 & _GEN_2133 : ~_GEN_2165 & _GEN_2133;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2262 = _GEN_44 ? ~_GEN_2217 & _GEN_2134 : ~_GEN_2166 & _GEN_2134;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2263 = _GEN_44 ? ~_GEN_2219 & _GEN_2135 : ~_GEN_2167 & _GEN_2135;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2264 = _GEN_44 ? ~_GEN_2221 & _GEN_2136 : ~_GEN_2168 & _GEN_2136;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2265 = _GEN_44 ? ~_GEN_2223 & _GEN_2137 : ~_GEN_2169 & _GEN_2137;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2266 = _GEN_44 ? ~_GEN_2225 & _GEN_2138 : ~_GEN_2170 & _GEN_2138;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2267 = _GEN_44 ? ~_GEN_2227 & _GEN_2139 : ~_GEN_2171 & _GEN_2139;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2268 = _GEN_44 ? ~_GEN_2229 & _GEN_2140 : ~_GEN_2172 & _GEN_2140;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2269 = _GEN_44 ? ~_GEN_2231 & _GEN_2141 : ~_GEN_2173 & _GEN_2141;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2270 = _GEN_44 ? ~_GEN_2233 & _GEN_2142 : ~_GEN_2174 & _GEN_2142;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2271 = _GEN_44 ? ~_GEN_2235 & _GEN_2143 : ~_GEN_2175 & _GEN_2143;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2272 = _GEN_44 ? ~_GEN_2237 & _GEN_2144 : ~_GEN_2176 & _GEN_2144;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2273 = _GEN_44 ? ~_GEN_2239 & _GEN_2145 : ~_GEN_2177 & _GEN_2145;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2274 = _GEN_44 ? ~_GEN_2241 & _GEN_2146 : ~_GEN_2178 & _GEN_2146;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2371 = rbk_row_1 & _GEN_1444;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2372 = rbk_row_1 & _GEN_1446;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2373 = rbk_row_1 & _GEN_1448;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2374 = rbk_row_1 & _GEN_1450;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2375 = rbk_row_1 & _GEN_1452;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2376 = rbk_row_1 & _GEN_1454;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2377 = rbk_row_1 & _GEN_1456;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2378 = rbk_row_1 & _GEN_1458;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2379 = rbk_row_1 & _GEN_1460;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2380 = rbk_row_1 & _GEN_1462;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2381 = rbk_row_1 & _GEN_1464;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2382 = rbk_row_1 & _GEN_1466;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2383 = rbk_row_1 & _GEN_1468;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2384 = rbk_row_1 & _GEN_1470;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2385 = rbk_row_1 & _GEN_1472;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2386 = rbk_row_1 & _GEN_1474;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2387 = rbk_row_1 & _GEN_1476;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2388 = rbk_row_1 & _GEN_1478;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2389 = rbk_row_1 & _GEN_1480;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2390 = rbk_row_1 & _GEN_1482;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2391 = rbk_row_1 & _GEN_1484;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2392 = rbk_row_1 & _GEN_1486;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2393 = rbk_row_1 & _GEN_1488;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2394 = rbk_row_1 & _GEN_1490;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2395 = rbk_row_1 & _GEN_1492;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2396 = rbk_row_1 & _GEN_1494;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2397 = rbk_row_1 & _GEN_1496;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2398 = rbk_row_1 & _GEN_1498;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2399 = rbk_row_1 & _GEN_1500;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2400 = rbk_row_1 & _GEN_1502;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2401 = rbk_row_1 & _GEN_1504;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2402 = rbk_row_1 & (&com_idx);	// rob.scala:236:20, :323:29, :425:44, :433:20, :434:30
    _GEN_2403 = io_brupdate_b1_mispredict_mask & rob_uop_1_0_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2404 = io_brupdate_b1_mispredict_mask & rob_uop_1_1_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2405 = io_brupdate_b1_mispredict_mask & rob_uop_1_2_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2406 = io_brupdate_b1_mispredict_mask & rob_uop_1_3_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2407 = io_brupdate_b1_mispredict_mask & rob_uop_1_4_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2408 = io_brupdate_b1_mispredict_mask & rob_uop_1_5_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2409 = io_brupdate_b1_mispredict_mask & rob_uop_1_6_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2410 = io_brupdate_b1_mispredict_mask & rob_uop_1_7_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2411 = io_brupdate_b1_mispredict_mask & rob_uop_1_8_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2412 = io_brupdate_b1_mispredict_mask & rob_uop_1_9_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2413 = io_brupdate_b1_mispredict_mask & rob_uop_1_10_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2414 = io_brupdate_b1_mispredict_mask & rob_uop_1_11_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2415 = io_brupdate_b1_mispredict_mask & rob_uop_1_12_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2416 = io_brupdate_b1_mispredict_mask & rob_uop_1_13_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2417 = io_brupdate_b1_mispredict_mask & rob_uop_1_14_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2418 = io_brupdate_b1_mispredict_mask & rob_uop_1_15_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2419 = io_brupdate_b1_mispredict_mask & rob_uop_1_16_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2420 = io_brupdate_b1_mispredict_mask & rob_uop_1_17_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2421 = io_brupdate_b1_mispredict_mask & rob_uop_1_18_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2422 = io_brupdate_b1_mispredict_mask & rob_uop_1_19_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2423 = io_brupdate_b1_mispredict_mask & rob_uop_1_20_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2424 = io_brupdate_b1_mispredict_mask & rob_uop_1_21_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2425 = io_brupdate_b1_mispredict_mask & rob_uop_1_22_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2426 = io_brupdate_b1_mispredict_mask & rob_uop_1_23_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2427 = io_brupdate_b1_mispredict_mask & rob_uop_1_24_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2428 = io_brupdate_b1_mispredict_mask & rob_uop_1_25_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2429 = io_brupdate_b1_mispredict_mask & rob_uop_1_26_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2430 = io_brupdate_b1_mispredict_mask & rob_uop_1_27_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2431 = io_brupdate_b1_mispredict_mask & rob_uop_1_28_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2432 = io_brupdate_b1_mispredict_mask & rob_uop_1_29_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2433 = io_brupdate_b1_mispredict_mask & rob_uop_1_30_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2434 = io_brupdate_b1_mispredict_mask & rob_uop_1_31_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2435 = io_enq_valids_2 & _GEN_147;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2436 = io_enq_valids_2 & _GEN_149;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2437 = io_enq_valids_2 & _GEN_151;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2438 = io_enq_valids_2 & _GEN_153;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2439 = io_enq_valids_2 & _GEN_155;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2440 = io_enq_valids_2 & _GEN_157;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2441 = io_enq_valids_2 & _GEN_159;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2442 = io_enq_valids_2 & _GEN_161;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2443 = io_enq_valids_2 & _GEN_163;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2444 = io_enq_valids_2 & _GEN_165;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2445 = io_enq_valids_2 & _GEN_167;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2446 = io_enq_valids_2 & _GEN_169;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2447 = io_enq_valids_2 & _GEN_171;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2448 = io_enq_valids_2 & _GEN_173;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2449 = io_enq_valids_2 & _GEN_175;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2450 = io_enq_valids_2 & _GEN_177;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2451 = io_enq_valids_2 & _GEN_179;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2452 = io_enq_valids_2 & _GEN_181;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2453 = io_enq_valids_2 & _GEN_183;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2454 = io_enq_valids_2 & _GEN_185;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2455 = io_enq_valids_2 & _GEN_187;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2456 = io_enq_valids_2 & _GEN_189;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2457 = io_enq_valids_2 & _GEN_191;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2458 = io_enq_valids_2 & _GEN_193;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2459 = io_enq_valids_2 & _GEN_195;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2460 = io_enq_valids_2 & _GEN_197;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2461 = io_enq_valids_2 & _GEN_199;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2462 = io_enq_valids_2 & _GEN_201;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2463 = io_enq_valids_2 & _GEN_203;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2464 = io_enq_valids_2 & _GEN_205;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2465 = io_enq_valids_2 & _GEN_207;	// rob.scala:307:32, :323:29, :324:31
    _GEN_2466 = io_enq_valids_2 & (&rob_tail);	// rob.scala:228:29, :307:32, :323:29, :324:31
    _GEN_2467 = _GEN_2435 ? ~_rob_bsy_T_4 : rob_bsy_2_0;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2468 = _GEN_2436 ? ~_rob_bsy_T_4 : rob_bsy_2_1;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2469 = _GEN_2437 ? ~_rob_bsy_T_4 : rob_bsy_2_2;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2470 = _GEN_2438 ? ~_rob_bsy_T_4 : rob_bsy_2_3;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2471 = _GEN_2439 ? ~_rob_bsy_T_4 : rob_bsy_2_4;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2472 = _GEN_2440 ? ~_rob_bsy_T_4 : rob_bsy_2_5;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2473 = _GEN_2441 ? ~_rob_bsy_T_4 : rob_bsy_2_6;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2474 = _GEN_2442 ? ~_rob_bsy_T_4 : rob_bsy_2_7;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2475 = _GEN_2443 ? ~_rob_bsy_T_4 : rob_bsy_2_8;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2476 = _GEN_2444 ? ~_rob_bsy_T_4 : rob_bsy_2_9;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2477 = _GEN_2445 ? ~_rob_bsy_T_4 : rob_bsy_2_10;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2478 = _GEN_2446 ? ~_rob_bsy_T_4 : rob_bsy_2_11;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2479 = _GEN_2447 ? ~_rob_bsy_T_4 : rob_bsy_2_12;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2480 = _GEN_2448 ? ~_rob_bsy_T_4 : rob_bsy_2_13;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2481 = _GEN_2449 ? ~_rob_bsy_T_4 : rob_bsy_2_14;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2482 = _GEN_2450 ? ~_rob_bsy_T_4 : rob_bsy_2_15;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2483 = _GEN_2451 ? ~_rob_bsy_T_4 : rob_bsy_2_16;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2484 = _GEN_2452 ? ~_rob_bsy_T_4 : rob_bsy_2_17;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2485 = _GEN_2453 ? ~_rob_bsy_T_4 : rob_bsy_2_18;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2486 = _GEN_2454 ? ~_rob_bsy_T_4 : rob_bsy_2_19;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2487 = _GEN_2455 ? ~_rob_bsy_T_4 : rob_bsy_2_20;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2488 = _GEN_2456 ? ~_rob_bsy_T_4 : rob_bsy_2_21;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2489 = _GEN_2457 ? ~_rob_bsy_T_4 : rob_bsy_2_22;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2490 = _GEN_2458 ? ~_rob_bsy_T_4 : rob_bsy_2_23;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2491 = _GEN_2459 ? ~_rob_bsy_T_4 : rob_bsy_2_24;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2492 = _GEN_2460 ? ~_rob_bsy_T_4 : rob_bsy_2_25;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2493 = _GEN_2461 ? ~_rob_bsy_T_4 : rob_bsy_2_26;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2494 = _GEN_2462 ? ~_rob_bsy_T_4 : rob_bsy_2_27;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2495 = _GEN_2463 ? ~_rob_bsy_T_4 : rob_bsy_2_28;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2496 = _GEN_2464 ? ~_rob_bsy_T_4 : rob_bsy_2_29;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2497 = _GEN_2465 ? ~_rob_bsy_T_4 : rob_bsy_2_30;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2498 = _GEN_2466 ? ~_rob_bsy_T_4 : rob_bsy_2_31;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_2499 = _GEN_2435 ? _rob_unsafe_T_14 : rob_unsafe_2_0;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2500 = _GEN_2436 ? _rob_unsafe_T_14 : rob_unsafe_2_1;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2501 = _GEN_2437 ? _rob_unsafe_T_14 : rob_unsafe_2_2;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2502 = _GEN_2438 ? _rob_unsafe_T_14 : rob_unsafe_2_3;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2503 = _GEN_2439 ? _rob_unsafe_T_14 : rob_unsafe_2_4;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2504 = _GEN_2440 ? _rob_unsafe_T_14 : rob_unsafe_2_5;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2505 = _GEN_2441 ? _rob_unsafe_T_14 : rob_unsafe_2_6;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2506 = _GEN_2442 ? _rob_unsafe_T_14 : rob_unsafe_2_7;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2507 = _GEN_2443 ? _rob_unsafe_T_14 : rob_unsafe_2_8;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2508 = _GEN_2444 ? _rob_unsafe_T_14 : rob_unsafe_2_9;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2509 = _GEN_2445 ? _rob_unsafe_T_14 : rob_unsafe_2_10;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2510 = _GEN_2446 ? _rob_unsafe_T_14 : rob_unsafe_2_11;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2511 = _GEN_2447 ? _rob_unsafe_T_14 : rob_unsafe_2_12;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2512 = _GEN_2448 ? _rob_unsafe_T_14 : rob_unsafe_2_13;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2513 = _GEN_2449 ? _rob_unsafe_T_14 : rob_unsafe_2_14;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2514 = _GEN_2450 ? _rob_unsafe_T_14 : rob_unsafe_2_15;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2515 = _GEN_2451 ? _rob_unsafe_T_14 : rob_unsafe_2_16;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2516 = _GEN_2452 ? _rob_unsafe_T_14 : rob_unsafe_2_17;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2517 = _GEN_2453 ? _rob_unsafe_T_14 : rob_unsafe_2_18;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2518 = _GEN_2454 ? _rob_unsafe_T_14 : rob_unsafe_2_19;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2519 = _GEN_2455 ? _rob_unsafe_T_14 : rob_unsafe_2_20;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2520 = _GEN_2456 ? _rob_unsafe_T_14 : rob_unsafe_2_21;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2521 = _GEN_2457 ? _rob_unsafe_T_14 : rob_unsafe_2_22;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2522 = _GEN_2458 ? _rob_unsafe_T_14 : rob_unsafe_2_23;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2523 = _GEN_2459 ? _rob_unsafe_T_14 : rob_unsafe_2_24;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2524 = _GEN_2460 ? _rob_unsafe_T_14 : rob_unsafe_2_25;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2525 = _GEN_2461 ? _rob_unsafe_T_14 : rob_unsafe_2_26;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2526 = _GEN_2462 ? _rob_unsafe_T_14 : rob_unsafe_2_27;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2527 = _GEN_2463 ? _rob_unsafe_T_14 : rob_unsafe_2_28;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2528 = _GEN_2464 ? _rob_unsafe_T_14 : rob_unsafe_2_29;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2529 = _GEN_2465 ? _rob_unsafe_T_14 : rob_unsafe_2_30;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2530 = _GEN_2466 ? _rob_unsafe_T_14 : rob_unsafe_2_31;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_2564 = _GEN_71 ? ~_GEN_2563 & _GEN_2467 : ~_GEN_2531 & _GEN_2467;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2566 = _GEN_71 ? ~_GEN_2565 & _GEN_2468 : ~_GEN_2532 & _GEN_2468;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2568 = _GEN_71 ? ~_GEN_2567 & _GEN_2469 : ~_GEN_2533 & _GEN_2469;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2570 = _GEN_71 ? ~_GEN_2569 & _GEN_2470 : ~_GEN_2534 & _GEN_2470;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2572 = _GEN_71 ? ~_GEN_2571 & _GEN_2471 : ~_GEN_2535 & _GEN_2471;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2574 = _GEN_71 ? ~_GEN_2573 & _GEN_2472 : ~_GEN_2536 & _GEN_2472;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2576 = _GEN_71 ? ~_GEN_2575 & _GEN_2473 : ~_GEN_2537 & _GEN_2473;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2578 = _GEN_71 ? ~_GEN_2577 & _GEN_2474 : ~_GEN_2538 & _GEN_2474;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2580 = _GEN_71 ? ~_GEN_2579 & _GEN_2475 : ~_GEN_2539 & _GEN_2475;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2582 = _GEN_71 ? ~_GEN_2581 & _GEN_2476 : ~_GEN_2540 & _GEN_2476;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2584 = _GEN_71 ? ~_GEN_2583 & _GEN_2477 : ~_GEN_2541 & _GEN_2477;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2586 = _GEN_71 ? ~_GEN_2585 & _GEN_2478 : ~_GEN_2542 & _GEN_2478;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2588 = _GEN_71 ? ~_GEN_2587 & _GEN_2479 : ~_GEN_2543 & _GEN_2479;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2590 = _GEN_71 ? ~_GEN_2589 & _GEN_2480 : ~_GEN_2544 & _GEN_2480;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2592 = _GEN_71 ? ~_GEN_2591 & _GEN_2481 : ~_GEN_2545 & _GEN_2481;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2594 = _GEN_71 ? ~_GEN_2593 & _GEN_2482 : ~_GEN_2546 & _GEN_2482;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2596 = _GEN_71 ? ~_GEN_2595 & _GEN_2483 : ~_GEN_2547 & _GEN_2483;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2598 = _GEN_71 ? ~_GEN_2597 & _GEN_2484 : ~_GEN_2548 & _GEN_2484;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2600 = _GEN_71 ? ~_GEN_2599 & _GEN_2485 : ~_GEN_2549 & _GEN_2485;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2602 = _GEN_71 ? ~_GEN_2601 & _GEN_2486 : ~_GEN_2550 & _GEN_2486;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2604 = _GEN_71 ? ~_GEN_2603 & _GEN_2487 : ~_GEN_2551 & _GEN_2487;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2606 = _GEN_71 ? ~_GEN_2605 & _GEN_2488 : ~_GEN_2552 & _GEN_2488;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2608 = _GEN_71 ? ~_GEN_2607 & _GEN_2489 : ~_GEN_2553 & _GEN_2489;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2610 = _GEN_71 ? ~_GEN_2609 & _GEN_2490 : ~_GEN_2554 & _GEN_2490;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2612 = _GEN_71 ? ~_GEN_2611 & _GEN_2491 : ~_GEN_2555 & _GEN_2491;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2614 = _GEN_71 ? ~_GEN_2613 & _GEN_2492 : ~_GEN_2556 & _GEN_2492;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2616 = _GEN_71 ? ~_GEN_2615 & _GEN_2493 : ~_GEN_2557 & _GEN_2493;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2618 = _GEN_71 ? ~_GEN_2617 & _GEN_2494 : ~_GEN_2558 & _GEN_2494;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2620 = _GEN_71 ? ~_GEN_2619 & _GEN_2495 : ~_GEN_2559 & _GEN_2495;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2622 = _GEN_71 ? ~_GEN_2621 & _GEN_2496 : ~_GEN_2560 & _GEN_2496;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2624 = _GEN_71 ? ~_GEN_2623 & _GEN_2497 : ~_GEN_2561 & _GEN_2497;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2626 = _GEN_71 ? ~_GEN_2625 & _GEN_2498 : ~_GEN_2562 & _GEN_2498;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_2627 = _GEN_71 ? ~_GEN_2563 & _GEN_2499 : ~_GEN_2531 & _GEN_2499;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2628 = _GEN_71 ? ~_GEN_2565 & _GEN_2500 : ~_GEN_2532 & _GEN_2500;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2629 = _GEN_71 ? ~_GEN_2567 & _GEN_2501 : ~_GEN_2533 & _GEN_2501;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2630 = _GEN_71 ? ~_GEN_2569 & _GEN_2502 : ~_GEN_2534 & _GEN_2502;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2631 = _GEN_71 ? ~_GEN_2571 & _GEN_2503 : ~_GEN_2535 & _GEN_2503;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2632 = _GEN_71 ? ~_GEN_2573 & _GEN_2504 : ~_GEN_2536 & _GEN_2504;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2633 = _GEN_71 ? ~_GEN_2575 & _GEN_2505 : ~_GEN_2537 & _GEN_2505;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2634 = _GEN_71 ? ~_GEN_2577 & _GEN_2506 : ~_GEN_2538 & _GEN_2506;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2635 = _GEN_71 ? ~_GEN_2579 & _GEN_2507 : ~_GEN_2539 & _GEN_2507;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2636 = _GEN_71 ? ~_GEN_2581 & _GEN_2508 : ~_GEN_2540 & _GEN_2508;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2637 = _GEN_71 ? ~_GEN_2583 & _GEN_2509 : ~_GEN_2541 & _GEN_2509;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2638 = _GEN_71 ? ~_GEN_2585 & _GEN_2510 : ~_GEN_2542 & _GEN_2510;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2639 = _GEN_71 ? ~_GEN_2587 & _GEN_2511 : ~_GEN_2543 & _GEN_2511;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2640 = _GEN_71 ? ~_GEN_2589 & _GEN_2512 : ~_GEN_2544 & _GEN_2512;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2641 = _GEN_71 ? ~_GEN_2591 & _GEN_2513 : ~_GEN_2545 & _GEN_2513;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2642 = _GEN_71 ? ~_GEN_2593 & _GEN_2514 : ~_GEN_2546 & _GEN_2514;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2643 = _GEN_71 ? ~_GEN_2595 & _GEN_2515 : ~_GEN_2547 & _GEN_2515;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2644 = _GEN_71 ? ~_GEN_2597 & _GEN_2516 : ~_GEN_2548 & _GEN_2516;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2645 = _GEN_71 ? ~_GEN_2599 & _GEN_2517 : ~_GEN_2549 & _GEN_2517;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2646 = _GEN_71 ? ~_GEN_2601 & _GEN_2518 : ~_GEN_2550 & _GEN_2518;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2647 = _GEN_71 ? ~_GEN_2603 & _GEN_2519 : ~_GEN_2551 & _GEN_2519;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2648 = _GEN_71 ? ~_GEN_2605 & _GEN_2520 : ~_GEN_2552 & _GEN_2520;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2649 = _GEN_71 ? ~_GEN_2607 & _GEN_2521 : ~_GEN_2553 & _GEN_2521;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2650 = _GEN_71 ? ~_GEN_2609 & _GEN_2522 : ~_GEN_2554 & _GEN_2522;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2651 = _GEN_71 ? ~_GEN_2611 & _GEN_2523 : ~_GEN_2555 & _GEN_2523;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2652 = _GEN_71 ? ~_GEN_2613 & _GEN_2524 : ~_GEN_2556 & _GEN_2524;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2653 = _GEN_71 ? ~_GEN_2615 & _GEN_2525 : ~_GEN_2557 & _GEN_2525;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2654 = _GEN_71 ? ~_GEN_2617 & _GEN_2526 : ~_GEN_2558 & _GEN_2526;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2655 = _GEN_71 ? ~_GEN_2619 & _GEN_2527 : ~_GEN_2559 & _GEN_2527;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2656 = _GEN_71 ? ~_GEN_2621 & _GEN_2528 : ~_GEN_2560 & _GEN_2528;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2657 = _GEN_71 ? ~_GEN_2623 & _GEN_2529 : ~_GEN_2561 & _GEN_2529;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2658 = _GEN_71 ? ~_GEN_2625 & _GEN_2530 : ~_GEN_2562 & _GEN_2530;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_2692 = _GEN_73 ? ~_GEN_2691 & _GEN_2564 : ~_GEN_2659 & _GEN_2564;	// rob.scala:346:{27,69}, :347:31
    _GEN_2694 = _GEN_73 ? ~_GEN_2693 & _GEN_2566 : ~_GEN_2660 & _GEN_2566;	// rob.scala:346:{27,69}, :347:31
    _GEN_2696 = _GEN_73 ? ~_GEN_2695 & _GEN_2568 : ~_GEN_2661 & _GEN_2568;	// rob.scala:346:{27,69}, :347:31
    _GEN_2698 = _GEN_73 ? ~_GEN_2697 & _GEN_2570 : ~_GEN_2662 & _GEN_2570;	// rob.scala:346:{27,69}, :347:31
    _GEN_2700 = _GEN_73 ? ~_GEN_2699 & _GEN_2572 : ~_GEN_2663 & _GEN_2572;	// rob.scala:346:{27,69}, :347:31
    _GEN_2702 = _GEN_73 ? ~_GEN_2701 & _GEN_2574 : ~_GEN_2664 & _GEN_2574;	// rob.scala:346:{27,69}, :347:31
    _GEN_2704 = _GEN_73 ? ~_GEN_2703 & _GEN_2576 : ~_GEN_2665 & _GEN_2576;	// rob.scala:346:{27,69}, :347:31
    _GEN_2706 = _GEN_73 ? ~_GEN_2705 & _GEN_2578 : ~_GEN_2666 & _GEN_2578;	// rob.scala:346:{27,69}, :347:31
    _GEN_2708 = _GEN_73 ? ~_GEN_2707 & _GEN_2580 : ~_GEN_2667 & _GEN_2580;	// rob.scala:346:{27,69}, :347:31
    _GEN_2710 = _GEN_73 ? ~_GEN_2709 & _GEN_2582 : ~_GEN_2668 & _GEN_2582;	// rob.scala:346:{27,69}, :347:31
    _GEN_2712 = _GEN_73 ? ~_GEN_2711 & _GEN_2584 : ~_GEN_2669 & _GEN_2584;	// rob.scala:346:{27,69}, :347:31
    _GEN_2714 = _GEN_73 ? ~_GEN_2713 & _GEN_2586 : ~_GEN_2670 & _GEN_2586;	// rob.scala:346:{27,69}, :347:31
    _GEN_2716 = _GEN_73 ? ~_GEN_2715 & _GEN_2588 : ~_GEN_2671 & _GEN_2588;	// rob.scala:346:{27,69}, :347:31
    _GEN_2718 = _GEN_73 ? ~_GEN_2717 & _GEN_2590 : ~_GEN_2672 & _GEN_2590;	// rob.scala:346:{27,69}, :347:31
    _GEN_2720 = _GEN_73 ? ~_GEN_2719 & _GEN_2592 : ~_GEN_2673 & _GEN_2592;	// rob.scala:346:{27,69}, :347:31
    _GEN_2722 = _GEN_73 ? ~_GEN_2721 & _GEN_2594 : ~_GEN_2674 & _GEN_2594;	// rob.scala:346:{27,69}, :347:31
    _GEN_2724 = _GEN_73 ? ~_GEN_2723 & _GEN_2596 : ~_GEN_2675 & _GEN_2596;	// rob.scala:346:{27,69}, :347:31
    _GEN_2726 = _GEN_73 ? ~_GEN_2725 & _GEN_2598 : ~_GEN_2676 & _GEN_2598;	// rob.scala:346:{27,69}, :347:31
    _GEN_2728 = _GEN_73 ? ~_GEN_2727 & _GEN_2600 : ~_GEN_2677 & _GEN_2600;	// rob.scala:346:{27,69}, :347:31
    _GEN_2730 = _GEN_73 ? ~_GEN_2729 & _GEN_2602 : ~_GEN_2678 & _GEN_2602;	// rob.scala:346:{27,69}, :347:31
    _GEN_2732 = _GEN_73 ? ~_GEN_2731 & _GEN_2604 : ~_GEN_2679 & _GEN_2604;	// rob.scala:346:{27,69}, :347:31
    _GEN_2734 = _GEN_73 ? ~_GEN_2733 & _GEN_2606 : ~_GEN_2680 & _GEN_2606;	// rob.scala:346:{27,69}, :347:31
    _GEN_2736 = _GEN_73 ? ~_GEN_2735 & _GEN_2608 : ~_GEN_2681 & _GEN_2608;	// rob.scala:346:{27,69}, :347:31
    _GEN_2738 = _GEN_73 ? ~_GEN_2737 & _GEN_2610 : ~_GEN_2682 & _GEN_2610;	// rob.scala:346:{27,69}, :347:31
    _GEN_2740 = _GEN_73 ? ~_GEN_2739 & _GEN_2612 : ~_GEN_2683 & _GEN_2612;	// rob.scala:346:{27,69}, :347:31
    _GEN_2742 = _GEN_73 ? ~_GEN_2741 & _GEN_2614 : ~_GEN_2684 & _GEN_2614;	// rob.scala:346:{27,69}, :347:31
    _GEN_2744 = _GEN_73 ? ~_GEN_2743 & _GEN_2616 : ~_GEN_2685 & _GEN_2616;	// rob.scala:346:{27,69}, :347:31
    _GEN_2746 = _GEN_73 ? ~_GEN_2745 & _GEN_2618 : ~_GEN_2686 & _GEN_2618;	// rob.scala:346:{27,69}, :347:31
    _GEN_2748 = _GEN_73 ? ~_GEN_2747 & _GEN_2620 : ~_GEN_2687 & _GEN_2620;	// rob.scala:346:{27,69}, :347:31
    _GEN_2750 = _GEN_73 ? ~_GEN_2749 & _GEN_2622 : ~_GEN_2688 & _GEN_2622;	// rob.scala:346:{27,69}, :347:31
    _GEN_2752 = _GEN_73 ? ~_GEN_2751 & _GEN_2624 : ~_GEN_2689 & _GEN_2624;	// rob.scala:346:{27,69}, :347:31
    _GEN_2754 = _GEN_73 ? ~_GEN_2753 & _GEN_2626 : ~_GEN_2690 & _GEN_2626;	// rob.scala:346:{27,69}, :347:31
    _GEN_2755 = _GEN_73 ? ~_GEN_2691 & _GEN_2627 : ~_GEN_2659 & _GEN_2627;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2756 = _GEN_73 ? ~_GEN_2693 & _GEN_2628 : ~_GEN_2660 & _GEN_2628;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2757 = _GEN_73 ? ~_GEN_2695 & _GEN_2629 : ~_GEN_2661 & _GEN_2629;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2758 = _GEN_73 ? ~_GEN_2697 & _GEN_2630 : ~_GEN_2662 & _GEN_2630;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2759 = _GEN_73 ? ~_GEN_2699 & _GEN_2631 : ~_GEN_2663 & _GEN_2631;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2760 = _GEN_73 ? ~_GEN_2701 & _GEN_2632 : ~_GEN_2664 & _GEN_2632;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2761 = _GEN_73 ? ~_GEN_2703 & _GEN_2633 : ~_GEN_2665 & _GEN_2633;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2762 = _GEN_73 ? ~_GEN_2705 & _GEN_2634 : ~_GEN_2666 & _GEN_2634;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2763 = _GEN_73 ? ~_GEN_2707 & _GEN_2635 : ~_GEN_2667 & _GEN_2635;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2764 = _GEN_73 ? ~_GEN_2709 & _GEN_2636 : ~_GEN_2668 & _GEN_2636;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2765 = _GEN_73 ? ~_GEN_2711 & _GEN_2637 : ~_GEN_2669 & _GEN_2637;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2766 = _GEN_73 ? ~_GEN_2713 & _GEN_2638 : ~_GEN_2670 & _GEN_2638;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2767 = _GEN_73 ? ~_GEN_2715 & _GEN_2639 : ~_GEN_2671 & _GEN_2639;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2768 = _GEN_73 ? ~_GEN_2717 & _GEN_2640 : ~_GEN_2672 & _GEN_2640;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2769 = _GEN_73 ? ~_GEN_2719 & _GEN_2641 : ~_GEN_2673 & _GEN_2641;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2770 = _GEN_73 ? ~_GEN_2721 & _GEN_2642 : ~_GEN_2674 & _GEN_2642;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2771 = _GEN_73 ? ~_GEN_2723 & _GEN_2643 : ~_GEN_2675 & _GEN_2643;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2772 = _GEN_73 ? ~_GEN_2725 & _GEN_2644 : ~_GEN_2676 & _GEN_2644;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2773 = _GEN_73 ? ~_GEN_2727 & _GEN_2645 : ~_GEN_2677 & _GEN_2645;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2774 = _GEN_73 ? ~_GEN_2729 & _GEN_2646 : ~_GEN_2678 & _GEN_2646;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2775 = _GEN_73 ? ~_GEN_2731 & _GEN_2647 : ~_GEN_2679 & _GEN_2647;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2776 = _GEN_73 ? ~_GEN_2733 & _GEN_2648 : ~_GEN_2680 & _GEN_2648;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2777 = _GEN_73 ? ~_GEN_2735 & _GEN_2649 : ~_GEN_2681 & _GEN_2649;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2778 = _GEN_73 ? ~_GEN_2737 & _GEN_2650 : ~_GEN_2682 & _GEN_2650;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2779 = _GEN_73 ? ~_GEN_2739 & _GEN_2651 : ~_GEN_2683 & _GEN_2651;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2780 = _GEN_73 ? ~_GEN_2741 & _GEN_2652 : ~_GEN_2684 & _GEN_2652;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2781 = _GEN_73 ? ~_GEN_2743 & _GEN_2653 : ~_GEN_2685 & _GEN_2653;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2782 = _GEN_73 ? ~_GEN_2745 & _GEN_2654 : ~_GEN_2686 & _GEN_2654;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2783 = _GEN_73 ? ~_GEN_2747 & _GEN_2655 : ~_GEN_2687 & _GEN_2655;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2784 = _GEN_73 ? ~_GEN_2749 & _GEN_2656 : ~_GEN_2688 & _GEN_2656;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2785 = _GEN_73 ? ~_GEN_2751 & _GEN_2657 : ~_GEN_2689 & _GEN_2657;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2786 = _GEN_73 ? ~_GEN_2753 & _GEN_2658 : ~_GEN_2690 & _GEN_2658;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2820 = _GEN_75 ? ~_GEN_2819 & _GEN_2692 : ~_GEN_2787 & _GEN_2692;	// rob.scala:346:{27,69}, :347:31
    _GEN_2822 = _GEN_75 ? ~_GEN_2821 & _GEN_2694 : ~_GEN_2788 & _GEN_2694;	// rob.scala:346:{27,69}, :347:31
    _GEN_2824 = _GEN_75 ? ~_GEN_2823 & _GEN_2696 : ~_GEN_2789 & _GEN_2696;	// rob.scala:346:{27,69}, :347:31
    _GEN_2826 = _GEN_75 ? ~_GEN_2825 & _GEN_2698 : ~_GEN_2790 & _GEN_2698;	// rob.scala:346:{27,69}, :347:31
    _GEN_2828 = _GEN_75 ? ~_GEN_2827 & _GEN_2700 : ~_GEN_2791 & _GEN_2700;	// rob.scala:346:{27,69}, :347:31
    _GEN_2830 = _GEN_75 ? ~_GEN_2829 & _GEN_2702 : ~_GEN_2792 & _GEN_2702;	// rob.scala:346:{27,69}, :347:31
    _GEN_2832 = _GEN_75 ? ~_GEN_2831 & _GEN_2704 : ~_GEN_2793 & _GEN_2704;	// rob.scala:346:{27,69}, :347:31
    _GEN_2834 = _GEN_75 ? ~_GEN_2833 & _GEN_2706 : ~_GEN_2794 & _GEN_2706;	// rob.scala:346:{27,69}, :347:31
    _GEN_2836 = _GEN_75 ? ~_GEN_2835 & _GEN_2708 : ~_GEN_2795 & _GEN_2708;	// rob.scala:346:{27,69}, :347:31
    _GEN_2838 = _GEN_75 ? ~_GEN_2837 & _GEN_2710 : ~_GEN_2796 & _GEN_2710;	// rob.scala:346:{27,69}, :347:31
    _GEN_2840 = _GEN_75 ? ~_GEN_2839 & _GEN_2712 : ~_GEN_2797 & _GEN_2712;	// rob.scala:346:{27,69}, :347:31
    _GEN_2842 = _GEN_75 ? ~_GEN_2841 & _GEN_2714 : ~_GEN_2798 & _GEN_2714;	// rob.scala:346:{27,69}, :347:31
    _GEN_2844 = _GEN_75 ? ~_GEN_2843 & _GEN_2716 : ~_GEN_2799 & _GEN_2716;	// rob.scala:346:{27,69}, :347:31
    _GEN_2846 = _GEN_75 ? ~_GEN_2845 & _GEN_2718 : ~_GEN_2800 & _GEN_2718;	// rob.scala:346:{27,69}, :347:31
    _GEN_2848 = _GEN_75 ? ~_GEN_2847 & _GEN_2720 : ~_GEN_2801 & _GEN_2720;	// rob.scala:346:{27,69}, :347:31
    _GEN_2850 = _GEN_75 ? ~_GEN_2849 & _GEN_2722 : ~_GEN_2802 & _GEN_2722;	// rob.scala:346:{27,69}, :347:31
    _GEN_2852 = _GEN_75 ? ~_GEN_2851 & _GEN_2724 : ~_GEN_2803 & _GEN_2724;	// rob.scala:346:{27,69}, :347:31
    _GEN_2854 = _GEN_75 ? ~_GEN_2853 & _GEN_2726 : ~_GEN_2804 & _GEN_2726;	// rob.scala:346:{27,69}, :347:31
    _GEN_2856 = _GEN_75 ? ~_GEN_2855 & _GEN_2728 : ~_GEN_2805 & _GEN_2728;	// rob.scala:346:{27,69}, :347:31
    _GEN_2858 = _GEN_75 ? ~_GEN_2857 & _GEN_2730 : ~_GEN_2806 & _GEN_2730;	// rob.scala:346:{27,69}, :347:31
    _GEN_2860 = _GEN_75 ? ~_GEN_2859 & _GEN_2732 : ~_GEN_2807 & _GEN_2732;	// rob.scala:346:{27,69}, :347:31
    _GEN_2862 = _GEN_75 ? ~_GEN_2861 & _GEN_2734 : ~_GEN_2808 & _GEN_2734;	// rob.scala:346:{27,69}, :347:31
    _GEN_2864 = _GEN_75 ? ~_GEN_2863 & _GEN_2736 : ~_GEN_2809 & _GEN_2736;	// rob.scala:346:{27,69}, :347:31
    _GEN_2866 = _GEN_75 ? ~_GEN_2865 & _GEN_2738 : ~_GEN_2810 & _GEN_2738;	// rob.scala:346:{27,69}, :347:31
    _GEN_2868 = _GEN_75 ? ~_GEN_2867 & _GEN_2740 : ~_GEN_2811 & _GEN_2740;	// rob.scala:346:{27,69}, :347:31
    _GEN_2870 = _GEN_75 ? ~_GEN_2869 & _GEN_2742 : ~_GEN_2812 & _GEN_2742;	// rob.scala:346:{27,69}, :347:31
    _GEN_2872 = _GEN_75 ? ~_GEN_2871 & _GEN_2744 : ~_GEN_2813 & _GEN_2744;	// rob.scala:346:{27,69}, :347:31
    _GEN_2874 = _GEN_75 ? ~_GEN_2873 & _GEN_2746 : ~_GEN_2814 & _GEN_2746;	// rob.scala:346:{27,69}, :347:31
    _GEN_2876 = _GEN_75 ? ~_GEN_2875 & _GEN_2748 : ~_GEN_2815 & _GEN_2748;	// rob.scala:346:{27,69}, :347:31
    _GEN_2878 = _GEN_75 ? ~_GEN_2877 & _GEN_2750 : ~_GEN_2816 & _GEN_2750;	// rob.scala:346:{27,69}, :347:31
    _GEN_2880 = _GEN_75 ? ~_GEN_2879 & _GEN_2752 : ~_GEN_2817 & _GEN_2752;	// rob.scala:346:{27,69}, :347:31
    _GEN_2882 = _GEN_75 ? ~_GEN_2881 & _GEN_2754 : ~_GEN_2818 & _GEN_2754;	// rob.scala:346:{27,69}, :347:31
    _GEN_2883 = _GEN_75 ? ~_GEN_2819 & _GEN_2755 : ~_GEN_2787 & _GEN_2755;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2884 = _GEN_75 ? ~_GEN_2821 & _GEN_2756 : ~_GEN_2788 & _GEN_2756;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2885 = _GEN_75 ? ~_GEN_2823 & _GEN_2757 : ~_GEN_2789 & _GEN_2757;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2886 = _GEN_75 ? ~_GEN_2825 & _GEN_2758 : ~_GEN_2790 & _GEN_2758;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2887 = _GEN_75 ? ~_GEN_2827 & _GEN_2759 : ~_GEN_2791 & _GEN_2759;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2888 = _GEN_75 ? ~_GEN_2829 & _GEN_2760 : ~_GEN_2792 & _GEN_2760;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2889 = _GEN_75 ? ~_GEN_2831 & _GEN_2761 : ~_GEN_2793 & _GEN_2761;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2890 = _GEN_75 ? ~_GEN_2833 & _GEN_2762 : ~_GEN_2794 & _GEN_2762;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2891 = _GEN_75 ? ~_GEN_2835 & _GEN_2763 : ~_GEN_2795 & _GEN_2763;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2892 = _GEN_75 ? ~_GEN_2837 & _GEN_2764 : ~_GEN_2796 & _GEN_2764;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2893 = _GEN_75 ? ~_GEN_2839 & _GEN_2765 : ~_GEN_2797 & _GEN_2765;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2894 = _GEN_75 ? ~_GEN_2841 & _GEN_2766 : ~_GEN_2798 & _GEN_2766;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2895 = _GEN_75 ? ~_GEN_2843 & _GEN_2767 : ~_GEN_2799 & _GEN_2767;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2896 = _GEN_75 ? ~_GEN_2845 & _GEN_2768 : ~_GEN_2800 & _GEN_2768;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2897 = _GEN_75 ? ~_GEN_2847 & _GEN_2769 : ~_GEN_2801 & _GEN_2769;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2898 = _GEN_75 ? ~_GEN_2849 & _GEN_2770 : ~_GEN_2802 & _GEN_2770;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2899 = _GEN_75 ? ~_GEN_2851 & _GEN_2771 : ~_GEN_2803 & _GEN_2771;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2900 = _GEN_75 ? ~_GEN_2853 & _GEN_2772 : ~_GEN_2804 & _GEN_2772;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2901 = _GEN_75 ? ~_GEN_2855 & _GEN_2773 : ~_GEN_2805 & _GEN_2773;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2902 = _GEN_75 ? ~_GEN_2857 & _GEN_2774 : ~_GEN_2806 & _GEN_2774;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2903 = _GEN_75 ? ~_GEN_2859 & _GEN_2775 : ~_GEN_2807 & _GEN_2775;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2904 = _GEN_75 ? ~_GEN_2861 & _GEN_2776 : ~_GEN_2808 & _GEN_2776;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2905 = _GEN_75 ? ~_GEN_2863 & _GEN_2777 : ~_GEN_2809 & _GEN_2777;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2906 = _GEN_75 ? ~_GEN_2865 & _GEN_2778 : ~_GEN_2810 & _GEN_2778;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2907 = _GEN_75 ? ~_GEN_2867 & _GEN_2779 : ~_GEN_2811 & _GEN_2779;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2908 = _GEN_75 ? ~_GEN_2869 & _GEN_2780 : ~_GEN_2812 & _GEN_2780;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2909 = _GEN_75 ? ~_GEN_2871 & _GEN_2781 : ~_GEN_2813 & _GEN_2781;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2910 = _GEN_75 ? ~_GEN_2873 & _GEN_2782 : ~_GEN_2814 & _GEN_2782;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2911 = _GEN_75 ? ~_GEN_2875 & _GEN_2783 : ~_GEN_2815 & _GEN_2783;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2912 = _GEN_75 ? ~_GEN_2877 & _GEN_2784 : ~_GEN_2816 & _GEN_2784;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2913 = _GEN_75 ? ~_GEN_2879 & _GEN_2785 : ~_GEN_2817 & _GEN_2785;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2914 = _GEN_75 ? ~_GEN_2881 & _GEN_2786 : ~_GEN_2818 & _GEN_2786;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2948 = _GEN_77 ? ~_GEN_2947 & _GEN_2820 : ~_GEN_2915 & _GEN_2820;	// rob.scala:346:{27,69}, :347:31
    _GEN_2950 = _GEN_77 ? ~_GEN_2949 & _GEN_2822 : ~_GEN_2916 & _GEN_2822;	// rob.scala:346:{27,69}, :347:31
    _GEN_2952 = _GEN_77 ? ~_GEN_2951 & _GEN_2824 : ~_GEN_2917 & _GEN_2824;	// rob.scala:346:{27,69}, :347:31
    _GEN_2954 = _GEN_77 ? ~_GEN_2953 & _GEN_2826 : ~_GEN_2918 & _GEN_2826;	// rob.scala:346:{27,69}, :347:31
    _GEN_2956 = _GEN_77 ? ~_GEN_2955 & _GEN_2828 : ~_GEN_2919 & _GEN_2828;	// rob.scala:346:{27,69}, :347:31
    _GEN_2958 = _GEN_77 ? ~_GEN_2957 & _GEN_2830 : ~_GEN_2920 & _GEN_2830;	// rob.scala:346:{27,69}, :347:31
    _GEN_2960 = _GEN_77 ? ~_GEN_2959 & _GEN_2832 : ~_GEN_2921 & _GEN_2832;	// rob.scala:346:{27,69}, :347:31
    _GEN_2962 = _GEN_77 ? ~_GEN_2961 & _GEN_2834 : ~_GEN_2922 & _GEN_2834;	// rob.scala:346:{27,69}, :347:31
    _GEN_2964 = _GEN_77 ? ~_GEN_2963 & _GEN_2836 : ~_GEN_2923 & _GEN_2836;	// rob.scala:346:{27,69}, :347:31
    _GEN_2966 = _GEN_77 ? ~_GEN_2965 & _GEN_2838 : ~_GEN_2924 & _GEN_2838;	// rob.scala:346:{27,69}, :347:31
    _GEN_2968 = _GEN_77 ? ~_GEN_2967 & _GEN_2840 : ~_GEN_2925 & _GEN_2840;	// rob.scala:346:{27,69}, :347:31
    _GEN_2970 = _GEN_77 ? ~_GEN_2969 & _GEN_2842 : ~_GEN_2926 & _GEN_2842;	// rob.scala:346:{27,69}, :347:31
    _GEN_2972 = _GEN_77 ? ~_GEN_2971 & _GEN_2844 : ~_GEN_2927 & _GEN_2844;	// rob.scala:346:{27,69}, :347:31
    _GEN_2974 = _GEN_77 ? ~_GEN_2973 & _GEN_2846 : ~_GEN_2928 & _GEN_2846;	// rob.scala:346:{27,69}, :347:31
    _GEN_2976 = _GEN_77 ? ~_GEN_2975 & _GEN_2848 : ~_GEN_2929 & _GEN_2848;	// rob.scala:346:{27,69}, :347:31
    _GEN_2978 = _GEN_77 ? ~_GEN_2977 & _GEN_2850 : ~_GEN_2930 & _GEN_2850;	// rob.scala:346:{27,69}, :347:31
    _GEN_2980 = _GEN_77 ? ~_GEN_2979 & _GEN_2852 : ~_GEN_2931 & _GEN_2852;	// rob.scala:346:{27,69}, :347:31
    _GEN_2982 = _GEN_77 ? ~_GEN_2981 & _GEN_2854 : ~_GEN_2932 & _GEN_2854;	// rob.scala:346:{27,69}, :347:31
    _GEN_2984 = _GEN_77 ? ~_GEN_2983 & _GEN_2856 : ~_GEN_2933 & _GEN_2856;	// rob.scala:346:{27,69}, :347:31
    _GEN_2986 = _GEN_77 ? ~_GEN_2985 & _GEN_2858 : ~_GEN_2934 & _GEN_2858;	// rob.scala:346:{27,69}, :347:31
    _GEN_2988 = _GEN_77 ? ~_GEN_2987 & _GEN_2860 : ~_GEN_2935 & _GEN_2860;	// rob.scala:346:{27,69}, :347:31
    _GEN_2990 = _GEN_77 ? ~_GEN_2989 & _GEN_2862 : ~_GEN_2936 & _GEN_2862;	// rob.scala:346:{27,69}, :347:31
    _GEN_2992 = _GEN_77 ? ~_GEN_2991 & _GEN_2864 : ~_GEN_2937 & _GEN_2864;	// rob.scala:346:{27,69}, :347:31
    _GEN_2994 = _GEN_77 ? ~_GEN_2993 & _GEN_2866 : ~_GEN_2938 & _GEN_2866;	// rob.scala:346:{27,69}, :347:31
    _GEN_2996 = _GEN_77 ? ~_GEN_2995 & _GEN_2868 : ~_GEN_2939 & _GEN_2868;	// rob.scala:346:{27,69}, :347:31
    _GEN_2998 = _GEN_77 ? ~_GEN_2997 & _GEN_2870 : ~_GEN_2940 & _GEN_2870;	// rob.scala:346:{27,69}, :347:31
    _GEN_3000 = _GEN_77 ? ~_GEN_2999 & _GEN_2872 : ~_GEN_2941 & _GEN_2872;	// rob.scala:346:{27,69}, :347:31
    _GEN_3002 = _GEN_77 ? ~_GEN_3001 & _GEN_2874 : ~_GEN_2942 & _GEN_2874;	// rob.scala:346:{27,69}, :347:31
    _GEN_3004 = _GEN_77 ? ~_GEN_3003 & _GEN_2876 : ~_GEN_2943 & _GEN_2876;	// rob.scala:346:{27,69}, :347:31
    _GEN_3006 = _GEN_77 ? ~_GEN_3005 & _GEN_2878 : ~_GEN_2944 & _GEN_2878;	// rob.scala:346:{27,69}, :347:31
    _GEN_3008 = _GEN_77 ? ~_GEN_3007 & _GEN_2880 : ~_GEN_2945 & _GEN_2880;	// rob.scala:346:{27,69}, :347:31
    _GEN_3010 = _GEN_77 ? ~_GEN_3009 & _GEN_2882 : ~_GEN_2946 & _GEN_2882;	// rob.scala:346:{27,69}, :347:31
    _GEN_3011 = _GEN_77 ? ~_GEN_2947 & _GEN_2883 : ~_GEN_2915 & _GEN_2883;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3012 = _GEN_77 ? ~_GEN_2949 & _GEN_2884 : ~_GEN_2916 & _GEN_2884;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3013 = _GEN_77 ? ~_GEN_2951 & _GEN_2885 : ~_GEN_2917 & _GEN_2885;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3014 = _GEN_77 ? ~_GEN_2953 & _GEN_2886 : ~_GEN_2918 & _GEN_2886;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3015 = _GEN_77 ? ~_GEN_2955 & _GEN_2887 : ~_GEN_2919 & _GEN_2887;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3016 = _GEN_77 ? ~_GEN_2957 & _GEN_2888 : ~_GEN_2920 & _GEN_2888;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3017 = _GEN_77 ? ~_GEN_2959 & _GEN_2889 : ~_GEN_2921 & _GEN_2889;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3018 = _GEN_77 ? ~_GEN_2961 & _GEN_2890 : ~_GEN_2922 & _GEN_2890;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3019 = _GEN_77 ? ~_GEN_2963 & _GEN_2891 : ~_GEN_2923 & _GEN_2891;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3020 = _GEN_77 ? ~_GEN_2965 & _GEN_2892 : ~_GEN_2924 & _GEN_2892;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3021 = _GEN_77 ? ~_GEN_2967 & _GEN_2893 : ~_GEN_2925 & _GEN_2893;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3022 = _GEN_77 ? ~_GEN_2969 & _GEN_2894 : ~_GEN_2926 & _GEN_2894;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3023 = _GEN_77 ? ~_GEN_2971 & _GEN_2895 : ~_GEN_2927 & _GEN_2895;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3024 = _GEN_77 ? ~_GEN_2973 & _GEN_2896 : ~_GEN_2928 & _GEN_2896;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3025 = _GEN_77 ? ~_GEN_2975 & _GEN_2897 : ~_GEN_2929 & _GEN_2897;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3026 = _GEN_77 ? ~_GEN_2977 & _GEN_2898 : ~_GEN_2930 & _GEN_2898;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3027 = _GEN_77 ? ~_GEN_2979 & _GEN_2899 : ~_GEN_2931 & _GEN_2899;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3028 = _GEN_77 ? ~_GEN_2981 & _GEN_2900 : ~_GEN_2932 & _GEN_2900;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3029 = _GEN_77 ? ~_GEN_2983 & _GEN_2901 : ~_GEN_2933 & _GEN_2901;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3030 = _GEN_77 ? ~_GEN_2985 & _GEN_2902 : ~_GEN_2934 & _GEN_2902;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3031 = _GEN_77 ? ~_GEN_2987 & _GEN_2903 : ~_GEN_2935 & _GEN_2903;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3032 = _GEN_77 ? ~_GEN_2989 & _GEN_2904 : ~_GEN_2936 & _GEN_2904;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3033 = _GEN_77 ? ~_GEN_2991 & _GEN_2905 : ~_GEN_2937 & _GEN_2905;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3034 = _GEN_77 ? ~_GEN_2993 & _GEN_2906 : ~_GEN_2938 & _GEN_2906;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3035 = _GEN_77 ? ~_GEN_2995 & _GEN_2907 : ~_GEN_2939 & _GEN_2907;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3036 = _GEN_77 ? ~_GEN_2997 & _GEN_2908 : ~_GEN_2940 & _GEN_2908;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3037 = _GEN_77 ? ~_GEN_2999 & _GEN_2909 : ~_GEN_2941 & _GEN_2909;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3038 = _GEN_77 ? ~_GEN_3001 & _GEN_2910 : ~_GEN_2942 & _GEN_2910;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3039 = _GEN_77 ? ~_GEN_3003 & _GEN_2911 : ~_GEN_2943 & _GEN_2911;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3040 = _GEN_77 ? ~_GEN_3005 & _GEN_2912 : ~_GEN_2944 & _GEN_2912;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3041 = _GEN_77 ? ~_GEN_3007 & _GEN_2913 : ~_GEN_2945 & _GEN_2913;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3042 = _GEN_77 ? ~_GEN_3009 & _GEN_2914 : ~_GEN_2946 & _GEN_2914;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3076 = _GEN_79 ? ~_GEN_3075 & _GEN_2948 : ~_GEN_3043 & _GEN_2948;	// rob.scala:346:{27,69}, :347:31
    _GEN_3078 = _GEN_79 ? ~_GEN_3077 & _GEN_2950 : ~_GEN_3044 & _GEN_2950;	// rob.scala:346:{27,69}, :347:31
    _GEN_3080 = _GEN_79 ? ~_GEN_3079 & _GEN_2952 : ~_GEN_3045 & _GEN_2952;	// rob.scala:346:{27,69}, :347:31
    _GEN_3082 = _GEN_79 ? ~_GEN_3081 & _GEN_2954 : ~_GEN_3046 & _GEN_2954;	// rob.scala:346:{27,69}, :347:31
    _GEN_3084 = _GEN_79 ? ~_GEN_3083 & _GEN_2956 : ~_GEN_3047 & _GEN_2956;	// rob.scala:346:{27,69}, :347:31
    _GEN_3086 = _GEN_79 ? ~_GEN_3085 & _GEN_2958 : ~_GEN_3048 & _GEN_2958;	// rob.scala:346:{27,69}, :347:31
    _GEN_3088 = _GEN_79 ? ~_GEN_3087 & _GEN_2960 : ~_GEN_3049 & _GEN_2960;	// rob.scala:346:{27,69}, :347:31
    _GEN_3090 = _GEN_79 ? ~_GEN_3089 & _GEN_2962 : ~_GEN_3050 & _GEN_2962;	// rob.scala:346:{27,69}, :347:31
    _GEN_3092 = _GEN_79 ? ~_GEN_3091 & _GEN_2964 : ~_GEN_3051 & _GEN_2964;	// rob.scala:346:{27,69}, :347:31
    _GEN_3094 = _GEN_79 ? ~_GEN_3093 & _GEN_2966 : ~_GEN_3052 & _GEN_2966;	// rob.scala:346:{27,69}, :347:31
    _GEN_3096 = _GEN_79 ? ~_GEN_3095 & _GEN_2968 : ~_GEN_3053 & _GEN_2968;	// rob.scala:346:{27,69}, :347:31
    _GEN_3098 = _GEN_79 ? ~_GEN_3097 & _GEN_2970 : ~_GEN_3054 & _GEN_2970;	// rob.scala:346:{27,69}, :347:31
    _GEN_3100 = _GEN_79 ? ~_GEN_3099 & _GEN_2972 : ~_GEN_3055 & _GEN_2972;	// rob.scala:346:{27,69}, :347:31
    _GEN_3102 = _GEN_79 ? ~_GEN_3101 & _GEN_2974 : ~_GEN_3056 & _GEN_2974;	// rob.scala:346:{27,69}, :347:31
    _GEN_3104 = _GEN_79 ? ~_GEN_3103 & _GEN_2976 : ~_GEN_3057 & _GEN_2976;	// rob.scala:346:{27,69}, :347:31
    _GEN_3106 = _GEN_79 ? ~_GEN_3105 & _GEN_2978 : ~_GEN_3058 & _GEN_2978;	// rob.scala:346:{27,69}, :347:31
    _GEN_3108 = _GEN_79 ? ~_GEN_3107 & _GEN_2980 : ~_GEN_3059 & _GEN_2980;	// rob.scala:346:{27,69}, :347:31
    _GEN_3110 = _GEN_79 ? ~_GEN_3109 & _GEN_2982 : ~_GEN_3060 & _GEN_2982;	// rob.scala:346:{27,69}, :347:31
    _GEN_3112 = _GEN_79 ? ~_GEN_3111 & _GEN_2984 : ~_GEN_3061 & _GEN_2984;	// rob.scala:346:{27,69}, :347:31
    _GEN_3114 = _GEN_79 ? ~_GEN_3113 & _GEN_2986 : ~_GEN_3062 & _GEN_2986;	// rob.scala:346:{27,69}, :347:31
    _GEN_3116 = _GEN_79 ? ~_GEN_3115 & _GEN_2988 : ~_GEN_3063 & _GEN_2988;	// rob.scala:346:{27,69}, :347:31
    _GEN_3118 = _GEN_79 ? ~_GEN_3117 & _GEN_2990 : ~_GEN_3064 & _GEN_2990;	// rob.scala:346:{27,69}, :347:31
    _GEN_3120 = _GEN_79 ? ~_GEN_3119 & _GEN_2992 : ~_GEN_3065 & _GEN_2992;	// rob.scala:346:{27,69}, :347:31
    _GEN_3122 = _GEN_79 ? ~_GEN_3121 & _GEN_2994 : ~_GEN_3066 & _GEN_2994;	// rob.scala:346:{27,69}, :347:31
    _GEN_3124 = _GEN_79 ? ~_GEN_3123 & _GEN_2996 : ~_GEN_3067 & _GEN_2996;	// rob.scala:346:{27,69}, :347:31
    _GEN_3126 = _GEN_79 ? ~_GEN_3125 & _GEN_2998 : ~_GEN_3068 & _GEN_2998;	// rob.scala:346:{27,69}, :347:31
    _GEN_3128 = _GEN_79 ? ~_GEN_3127 & _GEN_3000 : ~_GEN_3069 & _GEN_3000;	// rob.scala:346:{27,69}, :347:31
    _GEN_3130 = _GEN_79 ? ~_GEN_3129 & _GEN_3002 : ~_GEN_3070 & _GEN_3002;	// rob.scala:346:{27,69}, :347:31
    _GEN_3132 = _GEN_79 ? ~_GEN_3131 & _GEN_3004 : ~_GEN_3071 & _GEN_3004;	// rob.scala:346:{27,69}, :347:31
    _GEN_3134 = _GEN_79 ? ~_GEN_3133 & _GEN_3006 : ~_GEN_3072 & _GEN_3006;	// rob.scala:346:{27,69}, :347:31
    _GEN_3136 = _GEN_79 ? ~_GEN_3135 & _GEN_3008 : ~_GEN_3073 & _GEN_3008;	// rob.scala:346:{27,69}, :347:31
    _GEN_3138 = _GEN_79 ? ~_GEN_3137 & _GEN_3010 : ~_GEN_3074 & _GEN_3010;	// rob.scala:346:{27,69}, :347:31
    _GEN_3139 = _GEN_79 ? ~_GEN_3075 & _GEN_3011 : ~_GEN_3043 & _GEN_3011;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3140 = _GEN_79 ? ~_GEN_3077 & _GEN_3012 : ~_GEN_3044 & _GEN_3012;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3141 = _GEN_79 ? ~_GEN_3079 & _GEN_3013 : ~_GEN_3045 & _GEN_3013;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3142 = _GEN_79 ? ~_GEN_3081 & _GEN_3014 : ~_GEN_3046 & _GEN_3014;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3143 = _GEN_79 ? ~_GEN_3083 & _GEN_3015 : ~_GEN_3047 & _GEN_3015;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3144 = _GEN_79 ? ~_GEN_3085 & _GEN_3016 : ~_GEN_3048 & _GEN_3016;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3145 = _GEN_79 ? ~_GEN_3087 & _GEN_3017 : ~_GEN_3049 & _GEN_3017;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3146 = _GEN_79 ? ~_GEN_3089 & _GEN_3018 : ~_GEN_3050 & _GEN_3018;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3147 = _GEN_79 ? ~_GEN_3091 & _GEN_3019 : ~_GEN_3051 & _GEN_3019;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3148 = _GEN_79 ? ~_GEN_3093 & _GEN_3020 : ~_GEN_3052 & _GEN_3020;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3149 = _GEN_79 ? ~_GEN_3095 & _GEN_3021 : ~_GEN_3053 & _GEN_3021;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3150 = _GEN_79 ? ~_GEN_3097 & _GEN_3022 : ~_GEN_3054 & _GEN_3022;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3151 = _GEN_79 ? ~_GEN_3099 & _GEN_3023 : ~_GEN_3055 & _GEN_3023;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3152 = _GEN_79 ? ~_GEN_3101 & _GEN_3024 : ~_GEN_3056 & _GEN_3024;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3153 = _GEN_79 ? ~_GEN_3103 & _GEN_3025 : ~_GEN_3057 & _GEN_3025;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3154 = _GEN_79 ? ~_GEN_3105 & _GEN_3026 : ~_GEN_3058 & _GEN_3026;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3155 = _GEN_79 ? ~_GEN_3107 & _GEN_3027 : ~_GEN_3059 & _GEN_3027;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3156 = _GEN_79 ? ~_GEN_3109 & _GEN_3028 : ~_GEN_3060 & _GEN_3028;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3157 = _GEN_79 ? ~_GEN_3111 & _GEN_3029 : ~_GEN_3061 & _GEN_3029;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3158 = _GEN_79 ? ~_GEN_3113 & _GEN_3030 : ~_GEN_3062 & _GEN_3030;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3159 = _GEN_79 ? ~_GEN_3115 & _GEN_3031 : ~_GEN_3063 & _GEN_3031;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3160 = _GEN_79 ? ~_GEN_3117 & _GEN_3032 : ~_GEN_3064 & _GEN_3032;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3161 = _GEN_79 ? ~_GEN_3119 & _GEN_3033 : ~_GEN_3065 & _GEN_3033;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3162 = _GEN_79 ? ~_GEN_3121 & _GEN_3034 : ~_GEN_3066 & _GEN_3034;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3163 = _GEN_79 ? ~_GEN_3123 & _GEN_3035 : ~_GEN_3067 & _GEN_3035;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3164 = _GEN_79 ? ~_GEN_3125 & _GEN_3036 : ~_GEN_3068 & _GEN_3036;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3165 = _GEN_79 ? ~_GEN_3127 & _GEN_3037 : ~_GEN_3069 & _GEN_3037;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3166 = _GEN_79 ? ~_GEN_3129 & _GEN_3038 : ~_GEN_3070 & _GEN_3038;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3167 = _GEN_79 ? ~_GEN_3131 & _GEN_3039 : ~_GEN_3071 & _GEN_3039;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3168 = _GEN_79 ? ~_GEN_3133 & _GEN_3040 : ~_GEN_3072 & _GEN_3040;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3169 = _GEN_79 ? ~_GEN_3135 & _GEN_3041 : ~_GEN_3073 & _GEN_3041;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3170 = _GEN_79 ? ~_GEN_3137 & _GEN_3042 : ~_GEN_3074 & _GEN_3042;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3267 = rbk_row_2 & _GEN_1444;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3268 = rbk_row_2 & _GEN_1446;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3269 = rbk_row_2 & _GEN_1448;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3270 = rbk_row_2 & _GEN_1450;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3271 = rbk_row_2 & _GEN_1452;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3272 = rbk_row_2 & _GEN_1454;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3273 = rbk_row_2 & _GEN_1456;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3274 = rbk_row_2 & _GEN_1458;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3275 = rbk_row_2 & _GEN_1460;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3276 = rbk_row_2 & _GEN_1462;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3277 = rbk_row_2 & _GEN_1464;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3278 = rbk_row_2 & _GEN_1466;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3279 = rbk_row_2 & _GEN_1468;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3280 = rbk_row_2 & _GEN_1470;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3281 = rbk_row_2 & _GEN_1472;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3282 = rbk_row_2 & _GEN_1474;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3283 = rbk_row_2 & _GEN_1476;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3284 = rbk_row_2 & _GEN_1478;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3285 = rbk_row_2 & _GEN_1480;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3286 = rbk_row_2 & _GEN_1482;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3287 = rbk_row_2 & _GEN_1484;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3288 = rbk_row_2 & _GEN_1486;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3289 = rbk_row_2 & _GEN_1488;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3290 = rbk_row_2 & _GEN_1490;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3291 = rbk_row_2 & _GEN_1492;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3292 = rbk_row_2 & _GEN_1494;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3293 = rbk_row_2 & _GEN_1496;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3294 = rbk_row_2 & _GEN_1498;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3295 = rbk_row_2 & _GEN_1500;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3296 = rbk_row_2 & _GEN_1502;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3297 = rbk_row_2 & _GEN_1504;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_3298 = rbk_row_2 & (&com_idx);	// rob.scala:236:20, :323:29, :425:44, :433:20, :434:30
    _GEN_3299 = io_brupdate_b1_mispredict_mask & rob_uop_2_0_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3300 = io_brupdate_b1_mispredict_mask & rob_uop_2_1_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3301 = io_brupdate_b1_mispredict_mask & rob_uop_2_2_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3302 = io_brupdate_b1_mispredict_mask & rob_uop_2_3_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3303 = io_brupdate_b1_mispredict_mask & rob_uop_2_4_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3304 = io_brupdate_b1_mispredict_mask & rob_uop_2_5_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3305 = io_brupdate_b1_mispredict_mask & rob_uop_2_6_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3306 = io_brupdate_b1_mispredict_mask & rob_uop_2_7_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3307 = io_brupdate_b1_mispredict_mask & rob_uop_2_8_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3308 = io_brupdate_b1_mispredict_mask & rob_uop_2_9_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3309 = io_brupdate_b1_mispredict_mask & rob_uop_2_10_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3310 = io_brupdate_b1_mispredict_mask & rob_uop_2_11_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3311 = io_brupdate_b1_mispredict_mask & rob_uop_2_12_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3312 = io_brupdate_b1_mispredict_mask & rob_uop_2_13_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3313 = io_brupdate_b1_mispredict_mask & rob_uop_2_14_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3314 = io_brupdate_b1_mispredict_mask & rob_uop_2_15_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3315 = io_brupdate_b1_mispredict_mask & rob_uop_2_16_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3316 = io_brupdate_b1_mispredict_mask & rob_uop_2_17_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3317 = io_brupdate_b1_mispredict_mask & rob_uop_2_18_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3318 = io_brupdate_b1_mispredict_mask & rob_uop_2_19_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3319 = io_brupdate_b1_mispredict_mask & rob_uop_2_20_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3320 = io_brupdate_b1_mispredict_mask & rob_uop_2_21_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3321 = io_brupdate_b1_mispredict_mask & rob_uop_2_22_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3322 = io_brupdate_b1_mispredict_mask & rob_uop_2_23_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3323 = io_brupdate_b1_mispredict_mask & rob_uop_2_24_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3324 = io_brupdate_b1_mispredict_mask & rob_uop_2_25_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3325 = io_brupdate_b1_mispredict_mask & rob_uop_2_26_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3326 = io_brupdate_b1_mispredict_mask & rob_uop_2_27_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3327 = io_brupdate_b1_mispredict_mask & rob_uop_2_28_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3328 = io_brupdate_b1_mispredict_mask & rob_uop_2_29_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3329 = io_brupdate_b1_mispredict_mask & rob_uop_2_30_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3330 = io_brupdate_b1_mispredict_mask & rob_uop_2_31_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_3331 = io_enq_valids_3 & _GEN_147;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3332 = io_enq_valids_3 & _GEN_149;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3333 = io_enq_valids_3 & _GEN_151;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3334 = io_enq_valids_3 & _GEN_153;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3335 = io_enq_valids_3 & _GEN_155;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3336 = io_enq_valids_3 & _GEN_157;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3337 = io_enq_valids_3 & _GEN_159;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3338 = io_enq_valids_3 & _GEN_161;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3339 = io_enq_valids_3 & _GEN_163;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3340 = io_enq_valids_3 & _GEN_165;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3341 = io_enq_valids_3 & _GEN_167;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3342 = io_enq_valids_3 & _GEN_169;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3343 = io_enq_valids_3 & _GEN_171;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3344 = io_enq_valids_3 & _GEN_173;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3345 = io_enq_valids_3 & _GEN_175;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3346 = io_enq_valids_3 & _GEN_177;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3347 = io_enq_valids_3 & _GEN_179;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3348 = io_enq_valids_3 & _GEN_181;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3349 = io_enq_valids_3 & _GEN_183;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3350 = io_enq_valids_3 & _GEN_185;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3351 = io_enq_valids_3 & _GEN_187;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3352 = io_enq_valids_3 & _GEN_189;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3353 = io_enq_valids_3 & _GEN_191;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3354 = io_enq_valids_3 & _GEN_193;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3355 = io_enq_valids_3 & _GEN_195;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3356 = io_enq_valids_3 & _GEN_197;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3357 = io_enq_valids_3 & _GEN_199;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3358 = io_enq_valids_3 & _GEN_201;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3359 = io_enq_valids_3 & _GEN_203;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3360 = io_enq_valids_3 & _GEN_205;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3361 = io_enq_valids_3 & _GEN_207;	// rob.scala:307:32, :323:29, :324:31
    _GEN_3362 = io_enq_valids_3 & (&rob_tail);	// rob.scala:228:29, :307:32, :323:29, :324:31
    _GEN_3363 = _GEN_3331 ? ~_rob_bsy_T_6 : rob_bsy_3_0;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3364 = _GEN_3332 ? ~_rob_bsy_T_6 : rob_bsy_3_1;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3365 = _GEN_3333 ? ~_rob_bsy_T_6 : rob_bsy_3_2;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3366 = _GEN_3334 ? ~_rob_bsy_T_6 : rob_bsy_3_3;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3367 = _GEN_3335 ? ~_rob_bsy_T_6 : rob_bsy_3_4;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3368 = _GEN_3336 ? ~_rob_bsy_T_6 : rob_bsy_3_5;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3369 = _GEN_3337 ? ~_rob_bsy_T_6 : rob_bsy_3_6;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3370 = _GEN_3338 ? ~_rob_bsy_T_6 : rob_bsy_3_7;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3371 = _GEN_3339 ? ~_rob_bsy_T_6 : rob_bsy_3_8;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3372 = _GEN_3340 ? ~_rob_bsy_T_6 : rob_bsy_3_9;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3373 = _GEN_3341 ? ~_rob_bsy_T_6 : rob_bsy_3_10;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3374 = _GEN_3342 ? ~_rob_bsy_T_6 : rob_bsy_3_11;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3375 = _GEN_3343 ? ~_rob_bsy_T_6 : rob_bsy_3_12;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3376 = _GEN_3344 ? ~_rob_bsy_T_6 : rob_bsy_3_13;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3377 = _GEN_3345 ? ~_rob_bsy_T_6 : rob_bsy_3_14;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3378 = _GEN_3346 ? ~_rob_bsy_T_6 : rob_bsy_3_15;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3379 = _GEN_3347 ? ~_rob_bsy_T_6 : rob_bsy_3_16;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3380 = _GEN_3348 ? ~_rob_bsy_T_6 : rob_bsy_3_17;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3381 = _GEN_3349 ? ~_rob_bsy_T_6 : rob_bsy_3_18;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3382 = _GEN_3350 ? ~_rob_bsy_T_6 : rob_bsy_3_19;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3383 = _GEN_3351 ? ~_rob_bsy_T_6 : rob_bsy_3_20;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3384 = _GEN_3352 ? ~_rob_bsy_T_6 : rob_bsy_3_21;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3385 = _GEN_3353 ? ~_rob_bsy_T_6 : rob_bsy_3_22;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3386 = _GEN_3354 ? ~_rob_bsy_T_6 : rob_bsy_3_23;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3387 = _GEN_3355 ? ~_rob_bsy_T_6 : rob_bsy_3_24;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3388 = _GEN_3356 ? ~_rob_bsy_T_6 : rob_bsy_3_25;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3389 = _GEN_3357 ? ~_rob_bsy_T_6 : rob_bsy_3_26;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3390 = _GEN_3358 ? ~_rob_bsy_T_6 : rob_bsy_3_27;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3391 = _GEN_3359 ? ~_rob_bsy_T_6 : rob_bsy_3_28;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3392 = _GEN_3360 ? ~_rob_bsy_T_6 : rob_bsy_3_29;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3393 = _GEN_3361 ? ~_rob_bsy_T_6 : rob_bsy_3_30;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3394 = _GEN_3362 ? ~_rob_bsy_T_6 : rob_bsy_3_31;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_3395 = _GEN_3331 ? _rob_unsafe_T_19 : rob_unsafe_3_0;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3396 = _GEN_3332 ? _rob_unsafe_T_19 : rob_unsafe_3_1;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3397 = _GEN_3333 ? _rob_unsafe_T_19 : rob_unsafe_3_2;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3398 = _GEN_3334 ? _rob_unsafe_T_19 : rob_unsafe_3_3;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3399 = _GEN_3335 ? _rob_unsafe_T_19 : rob_unsafe_3_4;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3400 = _GEN_3336 ? _rob_unsafe_T_19 : rob_unsafe_3_5;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3401 = _GEN_3337 ? _rob_unsafe_T_19 : rob_unsafe_3_6;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3402 = _GEN_3338 ? _rob_unsafe_T_19 : rob_unsafe_3_7;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3403 = _GEN_3339 ? _rob_unsafe_T_19 : rob_unsafe_3_8;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3404 = _GEN_3340 ? _rob_unsafe_T_19 : rob_unsafe_3_9;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3405 = _GEN_3341 ? _rob_unsafe_T_19 : rob_unsafe_3_10;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3406 = _GEN_3342 ? _rob_unsafe_T_19 : rob_unsafe_3_11;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3407 = _GEN_3343 ? _rob_unsafe_T_19 : rob_unsafe_3_12;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3408 = _GEN_3344 ? _rob_unsafe_T_19 : rob_unsafe_3_13;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3409 = _GEN_3345 ? _rob_unsafe_T_19 : rob_unsafe_3_14;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3410 = _GEN_3346 ? _rob_unsafe_T_19 : rob_unsafe_3_15;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3411 = _GEN_3347 ? _rob_unsafe_T_19 : rob_unsafe_3_16;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3412 = _GEN_3348 ? _rob_unsafe_T_19 : rob_unsafe_3_17;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3413 = _GEN_3349 ? _rob_unsafe_T_19 : rob_unsafe_3_18;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3414 = _GEN_3350 ? _rob_unsafe_T_19 : rob_unsafe_3_19;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3415 = _GEN_3351 ? _rob_unsafe_T_19 : rob_unsafe_3_20;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3416 = _GEN_3352 ? _rob_unsafe_T_19 : rob_unsafe_3_21;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3417 = _GEN_3353 ? _rob_unsafe_T_19 : rob_unsafe_3_22;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3418 = _GEN_3354 ? _rob_unsafe_T_19 : rob_unsafe_3_23;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3419 = _GEN_3355 ? _rob_unsafe_T_19 : rob_unsafe_3_24;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3420 = _GEN_3356 ? _rob_unsafe_T_19 : rob_unsafe_3_25;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3421 = _GEN_3357 ? _rob_unsafe_T_19 : rob_unsafe_3_26;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3422 = _GEN_3358 ? _rob_unsafe_T_19 : rob_unsafe_3_27;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3423 = _GEN_3359 ? _rob_unsafe_T_19 : rob_unsafe_3_28;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3424 = _GEN_3360 ? _rob_unsafe_T_19 : rob_unsafe_3_29;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3425 = _GEN_3361 ? _rob_unsafe_T_19 : rob_unsafe_3_30;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3426 = _GEN_3362 ? _rob_unsafe_T_19 : rob_unsafe_3_31;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_3460 = _GEN_106 ? ~_GEN_3459 & _GEN_3363 : ~_GEN_3427 & _GEN_3363;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3462 = _GEN_106 ? ~_GEN_3461 & _GEN_3364 : ~_GEN_3428 & _GEN_3364;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3464 = _GEN_106 ? ~_GEN_3463 & _GEN_3365 : ~_GEN_3429 & _GEN_3365;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3466 = _GEN_106 ? ~_GEN_3465 & _GEN_3366 : ~_GEN_3430 & _GEN_3366;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3468 = _GEN_106 ? ~_GEN_3467 & _GEN_3367 : ~_GEN_3431 & _GEN_3367;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3470 = _GEN_106 ? ~_GEN_3469 & _GEN_3368 : ~_GEN_3432 & _GEN_3368;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3472 = _GEN_106 ? ~_GEN_3471 & _GEN_3369 : ~_GEN_3433 & _GEN_3369;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3474 = _GEN_106 ? ~_GEN_3473 & _GEN_3370 : ~_GEN_3434 & _GEN_3370;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3476 = _GEN_106 ? ~_GEN_3475 & _GEN_3371 : ~_GEN_3435 & _GEN_3371;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3478 = _GEN_106 ? ~_GEN_3477 & _GEN_3372 : ~_GEN_3436 & _GEN_3372;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3480 = _GEN_106 ? ~_GEN_3479 & _GEN_3373 : ~_GEN_3437 & _GEN_3373;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3482 = _GEN_106 ? ~_GEN_3481 & _GEN_3374 : ~_GEN_3438 & _GEN_3374;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3484 = _GEN_106 ? ~_GEN_3483 & _GEN_3375 : ~_GEN_3439 & _GEN_3375;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3486 = _GEN_106 ? ~_GEN_3485 & _GEN_3376 : ~_GEN_3440 & _GEN_3376;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3488 = _GEN_106 ? ~_GEN_3487 & _GEN_3377 : ~_GEN_3441 & _GEN_3377;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3490 = _GEN_106 ? ~_GEN_3489 & _GEN_3378 : ~_GEN_3442 & _GEN_3378;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3492 = _GEN_106 ? ~_GEN_3491 & _GEN_3379 : ~_GEN_3443 & _GEN_3379;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3494 = _GEN_106 ? ~_GEN_3493 & _GEN_3380 : ~_GEN_3444 & _GEN_3380;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3496 = _GEN_106 ? ~_GEN_3495 & _GEN_3381 : ~_GEN_3445 & _GEN_3381;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3498 = _GEN_106 ? ~_GEN_3497 & _GEN_3382 : ~_GEN_3446 & _GEN_3382;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3500 = _GEN_106 ? ~_GEN_3499 & _GEN_3383 : ~_GEN_3447 & _GEN_3383;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3502 = _GEN_106 ? ~_GEN_3501 & _GEN_3384 : ~_GEN_3448 & _GEN_3384;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3504 = _GEN_106 ? ~_GEN_3503 & _GEN_3385 : ~_GEN_3449 & _GEN_3385;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3506 = _GEN_106 ? ~_GEN_3505 & _GEN_3386 : ~_GEN_3450 & _GEN_3386;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3508 = _GEN_106 ? ~_GEN_3507 & _GEN_3387 : ~_GEN_3451 & _GEN_3387;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3510 = _GEN_106 ? ~_GEN_3509 & _GEN_3388 : ~_GEN_3452 & _GEN_3388;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3512 = _GEN_106 ? ~_GEN_3511 & _GEN_3389 : ~_GEN_3453 & _GEN_3389;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3514 = _GEN_106 ? ~_GEN_3513 & _GEN_3390 : ~_GEN_3454 & _GEN_3390;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3516 = _GEN_106 ? ~_GEN_3515 & _GEN_3391 : ~_GEN_3455 & _GEN_3391;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3518 = _GEN_106 ? ~_GEN_3517 & _GEN_3392 : ~_GEN_3456 & _GEN_3392;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3520 = _GEN_106 ? ~_GEN_3519 & _GEN_3393 : ~_GEN_3457 & _GEN_3393;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3522 = _GEN_106 ? ~_GEN_3521 & _GEN_3394 : ~_GEN_3458 & _GEN_3394;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_3523 = _GEN_106 ? ~_GEN_3459 & _GEN_3395 : ~_GEN_3427 & _GEN_3395;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3524 = _GEN_106 ? ~_GEN_3461 & _GEN_3396 : ~_GEN_3428 & _GEN_3396;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3525 = _GEN_106 ? ~_GEN_3463 & _GEN_3397 : ~_GEN_3429 & _GEN_3397;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3526 = _GEN_106 ? ~_GEN_3465 & _GEN_3398 : ~_GEN_3430 & _GEN_3398;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3527 = _GEN_106 ? ~_GEN_3467 & _GEN_3399 : ~_GEN_3431 & _GEN_3399;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3528 = _GEN_106 ? ~_GEN_3469 & _GEN_3400 : ~_GEN_3432 & _GEN_3400;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3529 = _GEN_106 ? ~_GEN_3471 & _GEN_3401 : ~_GEN_3433 & _GEN_3401;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3530 = _GEN_106 ? ~_GEN_3473 & _GEN_3402 : ~_GEN_3434 & _GEN_3402;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3531 = _GEN_106 ? ~_GEN_3475 & _GEN_3403 : ~_GEN_3435 & _GEN_3403;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3532 = _GEN_106 ? ~_GEN_3477 & _GEN_3404 : ~_GEN_3436 & _GEN_3404;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3533 = _GEN_106 ? ~_GEN_3479 & _GEN_3405 : ~_GEN_3437 & _GEN_3405;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3534 = _GEN_106 ? ~_GEN_3481 & _GEN_3406 : ~_GEN_3438 & _GEN_3406;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3535 = _GEN_106 ? ~_GEN_3483 & _GEN_3407 : ~_GEN_3439 & _GEN_3407;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3536 = _GEN_106 ? ~_GEN_3485 & _GEN_3408 : ~_GEN_3440 & _GEN_3408;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3537 = _GEN_106 ? ~_GEN_3487 & _GEN_3409 : ~_GEN_3441 & _GEN_3409;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3538 = _GEN_106 ? ~_GEN_3489 & _GEN_3410 : ~_GEN_3442 & _GEN_3410;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3539 = _GEN_106 ? ~_GEN_3491 & _GEN_3411 : ~_GEN_3443 & _GEN_3411;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3540 = _GEN_106 ? ~_GEN_3493 & _GEN_3412 : ~_GEN_3444 & _GEN_3412;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3541 = _GEN_106 ? ~_GEN_3495 & _GEN_3413 : ~_GEN_3445 & _GEN_3413;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3542 = _GEN_106 ? ~_GEN_3497 & _GEN_3414 : ~_GEN_3446 & _GEN_3414;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3543 = _GEN_106 ? ~_GEN_3499 & _GEN_3415 : ~_GEN_3447 & _GEN_3415;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3544 = _GEN_106 ? ~_GEN_3501 & _GEN_3416 : ~_GEN_3448 & _GEN_3416;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3545 = _GEN_106 ? ~_GEN_3503 & _GEN_3417 : ~_GEN_3449 & _GEN_3417;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3546 = _GEN_106 ? ~_GEN_3505 & _GEN_3418 : ~_GEN_3450 & _GEN_3418;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3547 = _GEN_106 ? ~_GEN_3507 & _GEN_3419 : ~_GEN_3451 & _GEN_3419;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3548 = _GEN_106 ? ~_GEN_3509 & _GEN_3420 : ~_GEN_3452 & _GEN_3420;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3549 = _GEN_106 ? ~_GEN_3511 & _GEN_3421 : ~_GEN_3453 & _GEN_3421;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3550 = _GEN_106 ? ~_GEN_3513 & _GEN_3422 : ~_GEN_3454 & _GEN_3422;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3551 = _GEN_106 ? ~_GEN_3515 & _GEN_3423 : ~_GEN_3455 & _GEN_3423;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3552 = _GEN_106 ? ~_GEN_3517 & _GEN_3424 : ~_GEN_3456 & _GEN_3424;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3553 = _GEN_106 ? ~_GEN_3519 & _GEN_3425 : ~_GEN_3457 & _GEN_3425;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3554 = _GEN_106 ? ~_GEN_3521 & _GEN_3426 : ~_GEN_3458 & _GEN_3426;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_3588 = _GEN_108 ? ~_GEN_3587 & _GEN_3460 : ~_GEN_3555 & _GEN_3460;	// rob.scala:346:{27,69}, :347:31
    _GEN_3590 = _GEN_108 ? ~_GEN_3589 & _GEN_3462 : ~_GEN_3556 & _GEN_3462;	// rob.scala:346:{27,69}, :347:31
    _GEN_3592 = _GEN_108 ? ~_GEN_3591 & _GEN_3464 : ~_GEN_3557 & _GEN_3464;	// rob.scala:346:{27,69}, :347:31
    _GEN_3594 = _GEN_108 ? ~_GEN_3593 & _GEN_3466 : ~_GEN_3558 & _GEN_3466;	// rob.scala:346:{27,69}, :347:31
    _GEN_3596 = _GEN_108 ? ~_GEN_3595 & _GEN_3468 : ~_GEN_3559 & _GEN_3468;	// rob.scala:346:{27,69}, :347:31
    _GEN_3598 = _GEN_108 ? ~_GEN_3597 & _GEN_3470 : ~_GEN_3560 & _GEN_3470;	// rob.scala:346:{27,69}, :347:31
    _GEN_3600 = _GEN_108 ? ~_GEN_3599 & _GEN_3472 : ~_GEN_3561 & _GEN_3472;	// rob.scala:346:{27,69}, :347:31
    _GEN_3602 = _GEN_108 ? ~_GEN_3601 & _GEN_3474 : ~_GEN_3562 & _GEN_3474;	// rob.scala:346:{27,69}, :347:31
    _GEN_3604 = _GEN_108 ? ~_GEN_3603 & _GEN_3476 : ~_GEN_3563 & _GEN_3476;	// rob.scala:346:{27,69}, :347:31
    _GEN_3606 = _GEN_108 ? ~_GEN_3605 & _GEN_3478 : ~_GEN_3564 & _GEN_3478;	// rob.scala:346:{27,69}, :347:31
    _GEN_3608 = _GEN_108 ? ~_GEN_3607 & _GEN_3480 : ~_GEN_3565 & _GEN_3480;	// rob.scala:346:{27,69}, :347:31
    _GEN_3610 = _GEN_108 ? ~_GEN_3609 & _GEN_3482 : ~_GEN_3566 & _GEN_3482;	// rob.scala:346:{27,69}, :347:31
    _GEN_3612 = _GEN_108 ? ~_GEN_3611 & _GEN_3484 : ~_GEN_3567 & _GEN_3484;	// rob.scala:346:{27,69}, :347:31
    _GEN_3614 = _GEN_108 ? ~_GEN_3613 & _GEN_3486 : ~_GEN_3568 & _GEN_3486;	// rob.scala:346:{27,69}, :347:31
    _GEN_3616 = _GEN_108 ? ~_GEN_3615 & _GEN_3488 : ~_GEN_3569 & _GEN_3488;	// rob.scala:346:{27,69}, :347:31
    _GEN_3618 = _GEN_108 ? ~_GEN_3617 & _GEN_3490 : ~_GEN_3570 & _GEN_3490;	// rob.scala:346:{27,69}, :347:31
    _GEN_3620 = _GEN_108 ? ~_GEN_3619 & _GEN_3492 : ~_GEN_3571 & _GEN_3492;	// rob.scala:346:{27,69}, :347:31
    _GEN_3622 = _GEN_108 ? ~_GEN_3621 & _GEN_3494 : ~_GEN_3572 & _GEN_3494;	// rob.scala:346:{27,69}, :347:31
    _GEN_3624 = _GEN_108 ? ~_GEN_3623 & _GEN_3496 : ~_GEN_3573 & _GEN_3496;	// rob.scala:346:{27,69}, :347:31
    _GEN_3626 = _GEN_108 ? ~_GEN_3625 & _GEN_3498 : ~_GEN_3574 & _GEN_3498;	// rob.scala:346:{27,69}, :347:31
    _GEN_3628 = _GEN_108 ? ~_GEN_3627 & _GEN_3500 : ~_GEN_3575 & _GEN_3500;	// rob.scala:346:{27,69}, :347:31
    _GEN_3630 = _GEN_108 ? ~_GEN_3629 & _GEN_3502 : ~_GEN_3576 & _GEN_3502;	// rob.scala:346:{27,69}, :347:31
    _GEN_3632 = _GEN_108 ? ~_GEN_3631 & _GEN_3504 : ~_GEN_3577 & _GEN_3504;	// rob.scala:346:{27,69}, :347:31
    _GEN_3634 = _GEN_108 ? ~_GEN_3633 & _GEN_3506 : ~_GEN_3578 & _GEN_3506;	// rob.scala:346:{27,69}, :347:31
    _GEN_3636 = _GEN_108 ? ~_GEN_3635 & _GEN_3508 : ~_GEN_3579 & _GEN_3508;	// rob.scala:346:{27,69}, :347:31
    _GEN_3638 = _GEN_108 ? ~_GEN_3637 & _GEN_3510 : ~_GEN_3580 & _GEN_3510;	// rob.scala:346:{27,69}, :347:31
    _GEN_3640 = _GEN_108 ? ~_GEN_3639 & _GEN_3512 : ~_GEN_3581 & _GEN_3512;	// rob.scala:346:{27,69}, :347:31
    _GEN_3642 = _GEN_108 ? ~_GEN_3641 & _GEN_3514 : ~_GEN_3582 & _GEN_3514;	// rob.scala:346:{27,69}, :347:31
    _GEN_3644 = _GEN_108 ? ~_GEN_3643 & _GEN_3516 : ~_GEN_3583 & _GEN_3516;	// rob.scala:346:{27,69}, :347:31
    _GEN_3646 = _GEN_108 ? ~_GEN_3645 & _GEN_3518 : ~_GEN_3584 & _GEN_3518;	// rob.scala:346:{27,69}, :347:31
    _GEN_3648 = _GEN_108 ? ~_GEN_3647 & _GEN_3520 : ~_GEN_3585 & _GEN_3520;	// rob.scala:346:{27,69}, :347:31
    _GEN_3650 = _GEN_108 ? ~_GEN_3649 & _GEN_3522 : ~_GEN_3586 & _GEN_3522;	// rob.scala:346:{27,69}, :347:31
    _GEN_3651 = _GEN_108 ? ~_GEN_3587 & _GEN_3523 : ~_GEN_3555 & _GEN_3523;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3652 = _GEN_108 ? ~_GEN_3589 & _GEN_3524 : ~_GEN_3556 & _GEN_3524;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3653 = _GEN_108 ? ~_GEN_3591 & _GEN_3525 : ~_GEN_3557 & _GEN_3525;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3654 = _GEN_108 ? ~_GEN_3593 & _GEN_3526 : ~_GEN_3558 & _GEN_3526;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3655 = _GEN_108 ? ~_GEN_3595 & _GEN_3527 : ~_GEN_3559 & _GEN_3527;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3656 = _GEN_108 ? ~_GEN_3597 & _GEN_3528 : ~_GEN_3560 & _GEN_3528;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3657 = _GEN_108 ? ~_GEN_3599 & _GEN_3529 : ~_GEN_3561 & _GEN_3529;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3658 = _GEN_108 ? ~_GEN_3601 & _GEN_3530 : ~_GEN_3562 & _GEN_3530;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3659 = _GEN_108 ? ~_GEN_3603 & _GEN_3531 : ~_GEN_3563 & _GEN_3531;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3660 = _GEN_108 ? ~_GEN_3605 & _GEN_3532 : ~_GEN_3564 & _GEN_3532;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3661 = _GEN_108 ? ~_GEN_3607 & _GEN_3533 : ~_GEN_3565 & _GEN_3533;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3662 = _GEN_108 ? ~_GEN_3609 & _GEN_3534 : ~_GEN_3566 & _GEN_3534;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3663 = _GEN_108 ? ~_GEN_3611 & _GEN_3535 : ~_GEN_3567 & _GEN_3535;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3664 = _GEN_108 ? ~_GEN_3613 & _GEN_3536 : ~_GEN_3568 & _GEN_3536;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3665 = _GEN_108 ? ~_GEN_3615 & _GEN_3537 : ~_GEN_3569 & _GEN_3537;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3666 = _GEN_108 ? ~_GEN_3617 & _GEN_3538 : ~_GEN_3570 & _GEN_3538;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3667 = _GEN_108 ? ~_GEN_3619 & _GEN_3539 : ~_GEN_3571 & _GEN_3539;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3668 = _GEN_108 ? ~_GEN_3621 & _GEN_3540 : ~_GEN_3572 & _GEN_3540;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3669 = _GEN_108 ? ~_GEN_3623 & _GEN_3541 : ~_GEN_3573 & _GEN_3541;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3670 = _GEN_108 ? ~_GEN_3625 & _GEN_3542 : ~_GEN_3574 & _GEN_3542;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3671 = _GEN_108 ? ~_GEN_3627 & _GEN_3543 : ~_GEN_3575 & _GEN_3543;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3672 = _GEN_108 ? ~_GEN_3629 & _GEN_3544 : ~_GEN_3576 & _GEN_3544;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3673 = _GEN_108 ? ~_GEN_3631 & _GEN_3545 : ~_GEN_3577 & _GEN_3545;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3674 = _GEN_108 ? ~_GEN_3633 & _GEN_3546 : ~_GEN_3578 & _GEN_3546;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3675 = _GEN_108 ? ~_GEN_3635 & _GEN_3547 : ~_GEN_3579 & _GEN_3547;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3676 = _GEN_108 ? ~_GEN_3637 & _GEN_3548 : ~_GEN_3580 & _GEN_3548;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3677 = _GEN_108 ? ~_GEN_3639 & _GEN_3549 : ~_GEN_3581 & _GEN_3549;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3678 = _GEN_108 ? ~_GEN_3641 & _GEN_3550 : ~_GEN_3582 & _GEN_3550;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3679 = _GEN_108 ? ~_GEN_3643 & _GEN_3551 : ~_GEN_3583 & _GEN_3551;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3680 = _GEN_108 ? ~_GEN_3645 & _GEN_3552 : ~_GEN_3584 & _GEN_3552;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3681 = _GEN_108 ? ~_GEN_3647 & _GEN_3553 : ~_GEN_3585 & _GEN_3553;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3682 = _GEN_108 ? ~_GEN_3649 & _GEN_3554 : ~_GEN_3586 & _GEN_3554;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3716 = _GEN_110 ? ~_GEN_3715 & _GEN_3588 : ~_GEN_3683 & _GEN_3588;	// rob.scala:346:{27,69}, :347:31
    _GEN_3718 = _GEN_110 ? ~_GEN_3717 & _GEN_3590 : ~_GEN_3684 & _GEN_3590;	// rob.scala:346:{27,69}, :347:31
    _GEN_3720 = _GEN_110 ? ~_GEN_3719 & _GEN_3592 : ~_GEN_3685 & _GEN_3592;	// rob.scala:346:{27,69}, :347:31
    _GEN_3722 = _GEN_110 ? ~_GEN_3721 & _GEN_3594 : ~_GEN_3686 & _GEN_3594;	// rob.scala:346:{27,69}, :347:31
    _GEN_3724 = _GEN_110 ? ~_GEN_3723 & _GEN_3596 : ~_GEN_3687 & _GEN_3596;	// rob.scala:346:{27,69}, :347:31
    _GEN_3726 = _GEN_110 ? ~_GEN_3725 & _GEN_3598 : ~_GEN_3688 & _GEN_3598;	// rob.scala:346:{27,69}, :347:31
    _GEN_3728 = _GEN_110 ? ~_GEN_3727 & _GEN_3600 : ~_GEN_3689 & _GEN_3600;	// rob.scala:346:{27,69}, :347:31
    _GEN_3730 = _GEN_110 ? ~_GEN_3729 & _GEN_3602 : ~_GEN_3690 & _GEN_3602;	// rob.scala:346:{27,69}, :347:31
    _GEN_3732 = _GEN_110 ? ~_GEN_3731 & _GEN_3604 : ~_GEN_3691 & _GEN_3604;	// rob.scala:346:{27,69}, :347:31
    _GEN_3734 = _GEN_110 ? ~_GEN_3733 & _GEN_3606 : ~_GEN_3692 & _GEN_3606;	// rob.scala:346:{27,69}, :347:31
    _GEN_3736 = _GEN_110 ? ~_GEN_3735 & _GEN_3608 : ~_GEN_3693 & _GEN_3608;	// rob.scala:346:{27,69}, :347:31
    _GEN_3738 = _GEN_110 ? ~_GEN_3737 & _GEN_3610 : ~_GEN_3694 & _GEN_3610;	// rob.scala:346:{27,69}, :347:31
    _GEN_3740 = _GEN_110 ? ~_GEN_3739 & _GEN_3612 : ~_GEN_3695 & _GEN_3612;	// rob.scala:346:{27,69}, :347:31
    _GEN_3742 = _GEN_110 ? ~_GEN_3741 & _GEN_3614 : ~_GEN_3696 & _GEN_3614;	// rob.scala:346:{27,69}, :347:31
    _GEN_3744 = _GEN_110 ? ~_GEN_3743 & _GEN_3616 : ~_GEN_3697 & _GEN_3616;	// rob.scala:346:{27,69}, :347:31
    _GEN_3746 = _GEN_110 ? ~_GEN_3745 & _GEN_3618 : ~_GEN_3698 & _GEN_3618;	// rob.scala:346:{27,69}, :347:31
    _GEN_3748 = _GEN_110 ? ~_GEN_3747 & _GEN_3620 : ~_GEN_3699 & _GEN_3620;	// rob.scala:346:{27,69}, :347:31
    _GEN_3750 = _GEN_110 ? ~_GEN_3749 & _GEN_3622 : ~_GEN_3700 & _GEN_3622;	// rob.scala:346:{27,69}, :347:31
    _GEN_3752 = _GEN_110 ? ~_GEN_3751 & _GEN_3624 : ~_GEN_3701 & _GEN_3624;	// rob.scala:346:{27,69}, :347:31
    _GEN_3754 = _GEN_110 ? ~_GEN_3753 & _GEN_3626 : ~_GEN_3702 & _GEN_3626;	// rob.scala:346:{27,69}, :347:31
    _GEN_3756 = _GEN_110 ? ~_GEN_3755 & _GEN_3628 : ~_GEN_3703 & _GEN_3628;	// rob.scala:346:{27,69}, :347:31
    _GEN_3758 = _GEN_110 ? ~_GEN_3757 & _GEN_3630 : ~_GEN_3704 & _GEN_3630;	// rob.scala:346:{27,69}, :347:31
    _GEN_3760 = _GEN_110 ? ~_GEN_3759 & _GEN_3632 : ~_GEN_3705 & _GEN_3632;	// rob.scala:346:{27,69}, :347:31
    _GEN_3762 = _GEN_110 ? ~_GEN_3761 & _GEN_3634 : ~_GEN_3706 & _GEN_3634;	// rob.scala:346:{27,69}, :347:31
    _GEN_3764 = _GEN_110 ? ~_GEN_3763 & _GEN_3636 : ~_GEN_3707 & _GEN_3636;	// rob.scala:346:{27,69}, :347:31
    _GEN_3766 = _GEN_110 ? ~_GEN_3765 & _GEN_3638 : ~_GEN_3708 & _GEN_3638;	// rob.scala:346:{27,69}, :347:31
    _GEN_3768 = _GEN_110 ? ~_GEN_3767 & _GEN_3640 : ~_GEN_3709 & _GEN_3640;	// rob.scala:346:{27,69}, :347:31
    _GEN_3770 = _GEN_110 ? ~_GEN_3769 & _GEN_3642 : ~_GEN_3710 & _GEN_3642;	// rob.scala:346:{27,69}, :347:31
    _GEN_3772 = _GEN_110 ? ~_GEN_3771 & _GEN_3644 : ~_GEN_3711 & _GEN_3644;	// rob.scala:346:{27,69}, :347:31
    _GEN_3774 = _GEN_110 ? ~_GEN_3773 & _GEN_3646 : ~_GEN_3712 & _GEN_3646;	// rob.scala:346:{27,69}, :347:31
    _GEN_3776 = _GEN_110 ? ~_GEN_3775 & _GEN_3648 : ~_GEN_3713 & _GEN_3648;	// rob.scala:346:{27,69}, :347:31
    _GEN_3778 = _GEN_110 ? ~_GEN_3777 & _GEN_3650 : ~_GEN_3714 & _GEN_3650;	// rob.scala:346:{27,69}, :347:31
    _GEN_3779 = _GEN_110 ? ~_GEN_3715 & _GEN_3651 : ~_GEN_3683 & _GEN_3651;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3780 = _GEN_110 ? ~_GEN_3717 & _GEN_3652 : ~_GEN_3684 & _GEN_3652;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3781 = _GEN_110 ? ~_GEN_3719 & _GEN_3653 : ~_GEN_3685 & _GEN_3653;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3782 = _GEN_110 ? ~_GEN_3721 & _GEN_3654 : ~_GEN_3686 & _GEN_3654;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3783 = _GEN_110 ? ~_GEN_3723 & _GEN_3655 : ~_GEN_3687 & _GEN_3655;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3784 = _GEN_110 ? ~_GEN_3725 & _GEN_3656 : ~_GEN_3688 & _GEN_3656;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3785 = _GEN_110 ? ~_GEN_3727 & _GEN_3657 : ~_GEN_3689 & _GEN_3657;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3786 = _GEN_110 ? ~_GEN_3729 & _GEN_3658 : ~_GEN_3690 & _GEN_3658;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3787 = _GEN_110 ? ~_GEN_3731 & _GEN_3659 : ~_GEN_3691 & _GEN_3659;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3788 = _GEN_110 ? ~_GEN_3733 & _GEN_3660 : ~_GEN_3692 & _GEN_3660;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3789 = _GEN_110 ? ~_GEN_3735 & _GEN_3661 : ~_GEN_3693 & _GEN_3661;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3790 = _GEN_110 ? ~_GEN_3737 & _GEN_3662 : ~_GEN_3694 & _GEN_3662;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3791 = _GEN_110 ? ~_GEN_3739 & _GEN_3663 : ~_GEN_3695 & _GEN_3663;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3792 = _GEN_110 ? ~_GEN_3741 & _GEN_3664 : ~_GEN_3696 & _GEN_3664;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3793 = _GEN_110 ? ~_GEN_3743 & _GEN_3665 : ~_GEN_3697 & _GEN_3665;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3794 = _GEN_110 ? ~_GEN_3745 & _GEN_3666 : ~_GEN_3698 & _GEN_3666;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3795 = _GEN_110 ? ~_GEN_3747 & _GEN_3667 : ~_GEN_3699 & _GEN_3667;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3796 = _GEN_110 ? ~_GEN_3749 & _GEN_3668 : ~_GEN_3700 & _GEN_3668;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3797 = _GEN_110 ? ~_GEN_3751 & _GEN_3669 : ~_GEN_3701 & _GEN_3669;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3798 = _GEN_110 ? ~_GEN_3753 & _GEN_3670 : ~_GEN_3702 & _GEN_3670;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3799 = _GEN_110 ? ~_GEN_3755 & _GEN_3671 : ~_GEN_3703 & _GEN_3671;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3800 = _GEN_110 ? ~_GEN_3757 & _GEN_3672 : ~_GEN_3704 & _GEN_3672;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3801 = _GEN_110 ? ~_GEN_3759 & _GEN_3673 : ~_GEN_3705 & _GEN_3673;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3802 = _GEN_110 ? ~_GEN_3761 & _GEN_3674 : ~_GEN_3706 & _GEN_3674;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3803 = _GEN_110 ? ~_GEN_3763 & _GEN_3675 : ~_GEN_3707 & _GEN_3675;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3804 = _GEN_110 ? ~_GEN_3765 & _GEN_3676 : ~_GEN_3708 & _GEN_3676;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3805 = _GEN_110 ? ~_GEN_3767 & _GEN_3677 : ~_GEN_3709 & _GEN_3677;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3806 = _GEN_110 ? ~_GEN_3769 & _GEN_3678 : ~_GEN_3710 & _GEN_3678;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3807 = _GEN_110 ? ~_GEN_3771 & _GEN_3679 : ~_GEN_3711 & _GEN_3679;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3808 = _GEN_110 ? ~_GEN_3773 & _GEN_3680 : ~_GEN_3712 & _GEN_3680;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3809 = _GEN_110 ? ~_GEN_3775 & _GEN_3681 : ~_GEN_3713 & _GEN_3681;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3810 = _GEN_110 ? ~_GEN_3777 & _GEN_3682 : ~_GEN_3714 & _GEN_3682;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3844 = _GEN_112 ? ~_GEN_3843 & _GEN_3716 : ~_GEN_3811 & _GEN_3716;	// rob.scala:346:{27,69}, :347:31
    _GEN_3846 = _GEN_112 ? ~_GEN_3845 & _GEN_3718 : ~_GEN_3812 & _GEN_3718;	// rob.scala:346:{27,69}, :347:31
    _GEN_3848 = _GEN_112 ? ~_GEN_3847 & _GEN_3720 : ~_GEN_3813 & _GEN_3720;	// rob.scala:346:{27,69}, :347:31
    _GEN_3850 = _GEN_112 ? ~_GEN_3849 & _GEN_3722 : ~_GEN_3814 & _GEN_3722;	// rob.scala:346:{27,69}, :347:31
    _GEN_3852 = _GEN_112 ? ~_GEN_3851 & _GEN_3724 : ~_GEN_3815 & _GEN_3724;	// rob.scala:346:{27,69}, :347:31
    _GEN_3854 = _GEN_112 ? ~_GEN_3853 & _GEN_3726 : ~_GEN_3816 & _GEN_3726;	// rob.scala:346:{27,69}, :347:31
    _GEN_3856 = _GEN_112 ? ~_GEN_3855 & _GEN_3728 : ~_GEN_3817 & _GEN_3728;	// rob.scala:346:{27,69}, :347:31
    _GEN_3858 = _GEN_112 ? ~_GEN_3857 & _GEN_3730 : ~_GEN_3818 & _GEN_3730;	// rob.scala:346:{27,69}, :347:31
    _GEN_3860 = _GEN_112 ? ~_GEN_3859 & _GEN_3732 : ~_GEN_3819 & _GEN_3732;	// rob.scala:346:{27,69}, :347:31
    _GEN_3862 = _GEN_112 ? ~_GEN_3861 & _GEN_3734 : ~_GEN_3820 & _GEN_3734;	// rob.scala:346:{27,69}, :347:31
    _GEN_3864 = _GEN_112 ? ~_GEN_3863 & _GEN_3736 : ~_GEN_3821 & _GEN_3736;	// rob.scala:346:{27,69}, :347:31
    _GEN_3866 = _GEN_112 ? ~_GEN_3865 & _GEN_3738 : ~_GEN_3822 & _GEN_3738;	// rob.scala:346:{27,69}, :347:31
    _GEN_3868 = _GEN_112 ? ~_GEN_3867 & _GEN_3740 : ~_GEN_3823 & _GEN_3740;	// rob.scala:346:{27,69}, :347:31
    _GEN_3870 = _GEN_112 ? ~_GEN_3869 & _GEN_3742 : ~_GEN_3824 & _GEN_3742;	// rob.scala:346:{27,69}, :347:31
    _GEN_3872 = _GEN_112 ? ~_GEN_3871 & _GEN_3744 : ~_GEN_3825 & _GEN_3744;	// rob.scala:346:{27,69}, :347:31
    _GEN_3874 = _GEN_112 ? ~_GEN_3873 & _GEN_3746 : ~_GEN_3826 & _GEN_3746;	// rob.scala:346:{27,69}, :347:31
    _GEN_3876 = _GEN_112 ? ~_GEN_3875 & _GEN_3748 : ~_GEN_3827 & _GEN_3748;	// rob.scala:346:{27,69}, :347:31
    _GEN_3878 = _GEN_112 ? ~_GEN_3877 & _GEN_3750 : ~_GEN_3828 & _GEN_3750;	// rob.scala:346:{27,69}, :347:31
    _GEN_3880 = _GEN_112 ? ~_GEN_3879 & _GEN_3752 : ~_GEN_3829 & _GEN_3752;	// rob.scala:346:{27,69}, :347:31
    _GEN_3882 = _GEN_112 ? ~_GEN_3881 & _GEN_3754 : ~_GEN_3830 & _GEN_3754;	// rob.scala:346:{27,69}, :347:31
    _GEN_3884 = _GEN_112 ? ~_GEN_3883 & _GEN_3756 : ~_GEN_3831 & _GEN_3756;	// rob.scala:346:{27,69}, :347:31
    _GEN_3886 = _GEN_112 ? ~_GEN_3885 & _GEN_3758 : ~_GEN_3832 & _GEN_3758;	// rob.scala:346:{27,69}, :347:31
    _GEN_3888 = _GEN_112 ? ~_GEN_3887 & _GEN_3760 : ~_GEN_3833 & _GEN_3760;	// rob.scala:346:{27,69}, :347:31
    _GEN_3890 = _GEN_112 ? ~_GEN_3889 & _GEN_3762 : ~_GEN_3834 & _GEN_3762;	// rob.scala:346:{27,69}, :347:31
    _GEN_3892 = _GEN_112 ? ~_GEN_3891 & _GEN_3764 : ~_GEN_3835 & _GEN_3764;	// rob.scala:346:{27,69}, :347:31
    _GEN_3894 = _GEN_112 ? ~_GEN_3893 & _GEN_3766 : ~_GEN_3836 & _GEN_3766;	// rob.scala:346:{27,69}, :347:31
    _GEN_3896 = _GEN_112 ? ~_GEN_3895 & _GEN_3768 : ~_GEN_3837 & _GEN_3768;	// rob.scala:346:{27,69}, :347:31
    _GEN_3898 = _GEN_112 ? ~_GEN_3897 & _GEN_3770 : ~_GEN_3838 & _GEN_3770;	// rob.scala:346:{27,69}, :347:31
    _GEN_3900 = _GEN_112 ? ~_GEN_3899 & _GEN_3772 : ~_GEN_3839 & _GEN_3772;	// rob.scala:346:{27,69}, :347:31
    _GEN_3902 = _GEN_112 ? ~_GEN_3901 & _GEN_3774 : ~_GEN_3840 & _GEN_3774;	// rob.scala:346:{27,69}, :347:31
    _GEN_3904 = _GEN_112 ? ~_GEN_3903 & _GEN_3776 : ~_GEN_3841 & _GEN_3776;	// rob.scala:346:{27,69}, :347:31
    _GEN_3906 = _GEN_112 ? ~_GEN_3905 & _GEN_3778 : ~_GEN_3842 & _GEN_3778;	// rob.scala:346:{27,69}, :347:31
    _GEN_3907 = _GEN_112 ? ~_GEN_3843 & _GEN_3779 : ~_GEN_3811 & _GEN_3779;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3908 = _GEN_112 ? ~_GEN_3845 & _GEN_3780 : ~_GEN_3812 & _GEN_3780;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3909 = _GEN_112 ? ~_GEN_3847 & _GEN_3781 : ~_GEN_3813 & _GEN_3781;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3910 = _GEN_112 ? ~_GEN_3849 & _GEN_3782 : ~_GEN_3814 & _GEN_3782;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3911 = _GEN_112 ? ~_GEN_3851 & _GEN_3783 : ~_GEN_3815 & _GEN_3783;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3912 = _GEN_112 ? ~_GEN_3853 & _GEN_3784 : ~_GEN_3816 & _GEN_3784;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3913 = _GEN_112 ? ~_GEN_3855 & _GEN_3785 : ~_GEN_3817 & _GEN_3785;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3914 = _GEN_112 ? ~_GEN_3857 & _GEN_3786 : ~_GEN_3818 & _GEN_3786;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3915 = _GEN_112 ? ~_GEN_3859 & _GEN_3787 : ~_GEN_3819 & _GEN_3787;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3916 = _GEN_112 ? ~_GEN_3861 & _GEN_3788 : ~_GEN_3820 & _GEN_3788;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3917 = _GEN_112 ? ~_GEN_3863 & _GEN_3789 : ~_GEN_3821 & _GEN_3789;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3918 = _GEN_112 ? ~_GEN_3865 & _GEN_3790 : ~_GEN_3822 & _GEN_3790;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3919 = _GEN_112 ? ~_GEN_3867 & _GEN_3791 : ~_GEN_3823 & _GEN_3791;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3920 = _GEN_112 ? ~_GEN_3869 & _GEN_3792 : ~_GEN_3824 & _GEN_3792;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3921 = _GEN_112 ? ~_GEN_3871 & _GEN_3793 : ~_GEN_3825 & _GEN_3793;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3922 = _GEN_112 ? ~_GEN_3873 & _GEN_3794 : ~_GEN_3826 & _GEN_3794;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3923 = _GEN_112 ? ~_GEN_3875 & _GEN_3795 : ~_GEN_3827 & _GEN_3795;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3924 = _GEN_112 ? ~_GEN_3877 & _GEN_3796 : ~_GEN_3828 & _GEN_3796;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3925 = _GEN_112 ? ~_GEN_3879 & _GEN_3797 : ~_GEN_3829 & _GEN_3797;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3926 = _GEN_112 ? ~_GEN_3881 & _GEN_3798 : ~_GEN_3830 & _GEN_3798;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3927 = _GEN_112 ? ~_GEN_3883 & _GEN_3799 : ~_GEN_3831 & _GEN_3799;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3928 = _GEN_112 ? ~_GEN_3885 & _GEN_3800 : ~_GEN_3832 & _GEN_3800;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3929 = _GEN_112 ? ~_GEN_3887 & _GEN_3801 : ~_GEN_3833 & _GEN_3801;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3930 = _GEN_112 ? ~_GEN_3889 & _GEN_3802 : ~_GEN_3834 & _GEN_3802;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3931 = _GEN_112 ? ~_GEN_3891 & _GEN_3803 : ~_GEN_3835 & _GEN_3803;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3932 = _GEN_112 ? ~_GEN_3893 & _GEN_3804 : ~_GEN_3836 & _GEN_3804;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3933 = _GEN_112 ? ~_GEN_3895 & _GEN_3805 : ~_GEN_3837 & _GEN_3805;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3934 = _GEN_112 ? ~_GEN_3897 & _GEN_3806 : ~_GEN_3838 & _GEN_3806;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3935 = _GEN_112 ? ~_GEN_3899 & _GEN_3807 : ~_GEN_3839 & _GEN_3807;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3936 = _GEN_112 ? ~_GEN_3901 & _GEN_3808 : ~_GEN_3840 & _GEN_3808;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3937 = _GEN_112 ? ~_GEN_3903 & _GEN_3809 : ~_GEN_3841 & _GEN_3809;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3938 = _GEN_112 ? ~_GEN_3905 & _GEN_3810 : ~_GEN_3842 & _GEN_3810;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_3972 = _GEN_114 ? ~_GEN_3971 & _GEN_3844 : ~_GEN_3939 & _GEN_3844;	// rob.scala:346:{27,69}, :347:31
    _GEN_3974 = _GEN_114 ? ~_GEN_3973 & _GEN_3846 : ~_GEN_3940 & _GEN_3846;	// rob.scala:346:{27,69}, :347:31
    _GEN_3976 = _GEN_114 ? ~_GEN_3975 & _GEN_3848 : ~_GEN_3941 & _GEN_3848;	// rob.scala:346:{27,69}, :347:31
    _GEN_3978 = _GEN_114 ? ~_GEN_3977 & _GEN_3850 : ~_GEN_3942 & _GEN_3850;	// rob.scala:346:{27,69}, :347:31
    _GEN_3980 = _GEN_114 ? ~_GEN_3979 & _GEN_3852 : ~_GEN_3943 & _GEN_3852;	// rob.scala:346:{27,69}, :347:31
    _GEN_3982 = _GEN_114 ? ~_GEN_3981 & _GEN_3854 : ~_GEN_3944 & _GEN_3854;	// rob.scala:346:{27,69}, :347:31
    _GEN_3984 = _GEN_114 ? ~_GEN_3983 & _GEN_3856 : ~_GEN_3945 & _GEN_3856;	// rob.scala:346:{27,69}, :347:31
    _GEN_3986 = _GEN_114 ? ~_GEN_3985 & _GEN_3858 : ~_GEN_3946 & _GEN_3858;	// rob.scala:346:{27,69}, :347:31
    _GEN_3988 = _GEN_114 ? ~_GEN_3987 & _GEN_3860 : ~_GEN_3947 & _GEN_3860;	// rob.scala:346:{27,69}, :347:31
    _GEN_3990 = _GEN_114 ? ~_GEN_3989 & _GEN_3862 : ~_GEN_3948 & _GEN_3862;	// rob.scala:346:{27,69}, :347:31
    _GEN_3992 = _GEN_114 ? ~_GEN_3991 & _GEN_3864 : ~_GEN_3949 & _GEN_3864;	// rob.scala:346:{27,69}, :347:31
    _GEN_3994 = _GEN_114 ? ~_GEN_3993 & _GEN_3866 : ~_GEN_3950 & _GEN_3866;	// rob.scala:346:{27,69}, :347:31
    _GEN_3996 = _GEN_114 ? ~_GEN_3995 & _GEN_3868 : ~_GEN_3951 & _GEN_3868;	// rob.scala:346:{27,69}, :347:31
    _GEN_3998 = _GEN_114 ? ~_GEN_3997 & _GEN_3870 : ~_GEN_3952 & _GEN_3870;	// rob.scala:346:{27,69}, :347:31
    _GEN_4000 = _GEN_114 ? ~_GEN_3999 & _GEN_3872 : ~_GEN_3953 & _GEN_3872;	// rob.scala:346:{27,69}, :347:31
    _GEN_4002 = _GEN_114 ? ~_GEN_4001 & _GEN_3874 : ~_GEN_3954 & _GEN_3874;	// rob.scala:346:{27,69}, :347:31
    _GEN_4004 = _GEN_114 ? ~_GEN_4003 & _GEN_3876 : ~_GEN_3955 & _GEN_3876;	// rob.scala:346:{27,69}, :347:31
    _GEN_4006 = _GEN_114 ? ~_GEN_4005 & _GEN_3878 : ~_GEN_3956 & _GEN_3878;	// rob.scala:346:{27,69}, :347:31
    _GEN_4008 = _GEN_114 ? ~_GEN_4007 & _GEN_3880 : ~_GEN_3957 & _GEN_3880;	// rob.scala:346:{27,69}, :347:31
    _GEN_4010 = _GEN_114 ? ~_GEN_4009 & _GEN_3882 : ~_GEN_3958 & _GEN_3882;	// rob.scala:346:{27,69}, :347:31
    _GEN_4012 = _GEN_114 ? ~_GEN_4011 & _GEN_3884 : ~_GEN_3959 & _GEN_3884;	// rob.scala:346:{27,69}, :347:31
    _GEN_4014 = _GEN_114 ? ~_GEN_4013 & _GEN_3886 : ~_GEN_3960 & _GEN_3886;	// rob.scala:346:{27,69}, :347:31
    _GEN_4016 = _GEN_114 ? ~_GEN_4015 & _GEN_3888 : ~_GEN_3961 & _GEN_3888;	// rob.scala:346:{27,69}, :347:31
    _GEN_4018 = _GEN_114 ? ~_GEN_4017 & _GEN_3890 : ~_GEN_3962 & _GEN_3890;	// rob.scala:346:{27,69}, :347:31
    _GEN_4020 = _GEN_114 ? ~_GEN_4019 & _GEN_3892 : ~_GEN_3963 & _GEN_3892;	// rob.scala:346:{27,69}, :347:31
    _GEN_4022 = _GEN_114 ? ~_GEN_4021 & _GEN_3894 : ~_GEN_3964 & _GEN_3894;	// rob.scala:346:{27,69}, :347:31
    _GEN_4024 = _GEN_114 ? ~_GEN_4023 & _GEN_3896 : ~_GEN_3965 & _GEN_3896;	// rob.scala:346:{27,69}, :347:31
    _GEN_4026 = _GEN_114 ? ~_GEN_4025 & _GEN_3898 : ~_GEN_3966 & _GEN_3898;	// rob.scala:346:{27,69}, :347:31
    _GEN_4028 = _GEN_114 ? ~_GEN_4027 & _GEN_3900 : ~_GEN_3967 & _GEN_3900;	// rob.scala:346:{27,69}, :347:31
    _GEN_4030 = _GEN_114 ? ~_GEN_4029 & _GEN_3902 : ~_GEN_3968 & _GEN_3902;	// rob.scala:346:{27,69}, :347:31
    _GEN_4032 = _GEN_114 ? ~_GEN_4031 & _GEN_3904 : ~_GEN_3969 & _GEN_3904;	// rob.scala:346:{27,69}, :347:31
    _GEN_4034 = _GEN_114 ? ~_GEN_4033 & _GEN_3906 : ~_GEN_3970 & _GEN_3906;	// rob.scala:346:{27,69}, :347:31
    _GEN_4035 = _GEN_114 ? ~_GEN_3971 & _GEN_3907 : ~_GEN_3939 & _GEN_3907;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4036 = _GEN_114 ? ~_GEN_3973 & _GEN_3908 : ~_GEN_3940 & _GEN_3908;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4037 = _GEN_114 ? ~_GEN_3975 & _GEN_3909 : ~_GEN_3941 & _GEN_3909;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4038 = _GEN_114 ? ~_GEN_3977 & _GEN_3910 : ~_GEN_3942 & _GEN_3910;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4039 = _GEN_114 ? ~_GEN_3979 & _GEN_3911 : ~_GEN_3943 & _GEN_3911;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4040 = _GEN_114 ? ~_GEN_3981 & _GEN_3912 : ~_GEN_3944 & _GEN_3912;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4041 = _GEN_114 ? ~_GEN_3983 & _GEN_3913 : ~_GEN_3945 & _GEN_3913;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4042 = _GEN_114 ? ~_GEN_3985 & _GEN_3914 : ~_GEN_3946 & _GEN_3914;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4043 = _GEN_114 ? ~_GEN_3987 & _GEN_3915 : ~_GEN_3947 & _GEN_3915;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4044 = _GEN_114 ? ~_GEN_3989 & _GEN_3916 : ~_GEN_3948 & _GEN_3916;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4045 = _GEN_114 ? ~_GEN_3991 & _GEN_3917 : ~_GEN_3949 & _GEN_3917;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4046 = _GEN_114 ? ~_GEN_3993 & _GEN_3918 : ~_GEN_3950 & _GEN_3918;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4047 = _GEN_114 ? ~_GEN_3995 & _GEN_3919 : ~_GEN_3951 & _GEN_3919;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4048 = _GEN_114 ? ~_GEN_3997 & _GEN_3920 : ~_GEN_3952 & _GEN_3920;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4049 = _GEN_114 ? ~_GEN_3999 & _GEN_3921 : ~_GEN_3953 & _GEN_3921;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4050 = _GEN_114 ? ~_GEN_4001 & _GEN_3922 : ~_GEN_3954 & _GEN_3922;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4051 = _GEN_114 ? ~_GEN_4003 & _GEN_3923 : ~_GEN_3955 & _GEN_3923;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4052 = _GEN_114 ? ~_GEN_4005 & _GEN_3924 : ~_GEN_3956 & _GEN_3924;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4053 = _GEN_114 ? ~_GEN_4007 & _GEN_3925 : ~_GEN_3957 & _GEN_3925;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4054 = _GEN_114 ? ~_GEN_4009 & _GEN_3926 : ~_GEN_3958 & _GEN_3926;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4055 = _GEN_114 ? ~_GEN_4011 & _GEN_3927 : ~_GEN_3959 & _GEN_3927;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4056 = _GEN_114 ? ~_GEN_4013 & _GEN_3928 : ~_GEN_3960 & _GEN_3928;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4057 = _GEN_114 ? ~_GEN_4015 & _GEN_3929 : ~_GEN_3961 & _GEN_3929;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4058 = _GEN_114 ? ~_GEN_4017 & _GEN_3930 : ~_GEN_3962 & _GEN_3930;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4059 = _GEN_114 ? ~_GEN_4019 & _GEN_3931 : ~_GEN_3963 & _GEN_3931;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4060 = _GEN_114 ? ~_GEN_4021 & _GEN_3932 : ~_GEN_3964 & _GEN_3932;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4061 = _GEN_114 ? ~_GEN_4023 & _GEN_3933 : ~_GEN_3965 & _GEN_3933;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4062 = _GEN_114 ? ~_GEN_4025 & _GEN_3934 : ~_GEN_3966 & _GEN_3934;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4063 = _GEN_114 ? ~_GEN_4027 & _GEN_3935 : ~_GEN_3967 & _GEN_3935;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4064 = _GEN_114 ? ~_GEN_4029 & _GEN_3936 : ~_GEN_3968 & _GEN_3936;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4065 = _GEN_114 ? ~_GEN_4031 & _GEN_3937 : ~_GEN_3969 & _GEN_3937;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4066 = _GEN_114 ? ~_GEN_4033 & _GEN_3938 : ~_GEN_3970 & _GEN_3938;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_4163 = rbk_row_3 & _GEN_1444;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4164 = rbk_row_3 & _GEN_1446;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4165 = rbk_row_3 & _GEN_1448;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4166 = rbk_row_3 & _GEN_1450;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4167 = rbk_row_3 & _GEN_1452;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4168 = rbk_row_3 & _GEN_1454;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4169 = rbk_row_3 & _GEN_1456;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4170 = rbk_row_3 & _GEN_1458;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4171 = rbk_row_3 & _GEN_1460;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4172 = rbk_row_3 & _GEN_1462;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4173 = rbk_row_3 & _GEN_1464;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4174 = rbk_row_3 & _GEN_1466;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4175 = rbk_row_3 & _GEN_1468;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4176 = rbk_row_3 & _GEN_1470;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4177 = rbk_row_3 & _GEN_1472;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4178 = rbk_row_3 & _GEN_1474;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4179 = rbk_row_3 & _GEN_1476;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4180 = rbk_row_3 & _GEN_1478;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4181 = rbk_row_3 & _GEN_1480;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4182 = rbk_row_3 & _GEN_1482;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4183 = rbk_row_3 & _GEN_1484;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4184 = rbk_row_3 & _GEN_1486;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4185 = rbk_row_3 & _GEN_1488;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4186 = rbk_row_3 & _GEN_1490;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4187 = rbk_row_3 & _GEN_1492;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4188 = rbk_row_3 & _GEN_1494;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4189 = rbk_row_3 & _GEN_1496;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4190 = rbk_row_3 & _GEN_1498;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4191 = rbk_row_3 & _GEN_1500;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4192 = rbk_row_3 & _GEN_1502;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4193 = rbk_row_3 & _GEN_1504;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_4194 = rbk_row_3 & (&com_idx);	// rob.scala:236:20, :323:29, :425:44, :433:20, :434:30
    _GEN_4195 = io_brupdate_b1_mispredict_mask & rob_uop_3_0_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4196 = io_brupdate_b1_mispredict_mask & rob_uop_3_1_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4197 = io_brupdate_b1_mispredict_mask & rob_uop_3_2_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4198 = io_brupdate_b1_mispredict_mask & rob_uop_3_3_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4199 = io_brupdate_b1_mispredict_mask & rob_uop_3_4_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4200 = io_brupdate_b1_mispredict_mask & rob_uop_3_5_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4201 = io_brupdate_b1_mispredict_mask & rob_uop_3_6_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4202 = io_brupdate_b1_mispredict_mask & rob_uop_3_7_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4203 = io_brupdate_b1_mispredict_mask & rob_uop_3_8_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4204 = io_brupdate_b1_mispredict_mask & rob_uop_3_9_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4205 = io_brupdate_b1_mispredict_mask & rob_uop_3_10_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4206 = io_brupdate_b1_mispredict_mask & rob_uop_3_11_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4207 = io_brupdate_b1_mispredict_mask & rob_uop_3_12_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4208 = io_brupdate_b1_mispredict_mask & rob_uop_3_13_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4209 = io_brupdate_b1_mispredict_mask & rob_uop_3_14_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4210 = io_brupdate_b1_mispredict_mask & rob_uop_3_15_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4211 = io_brupdate_b1_mispredict_mask & rob_uop_3_16_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4212 = io_brupdate_b1_mispredict_mask & rob_uop_3_17_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4213 = io_brupdate_b1_mispredict_mask & rob_uop_3_18_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4214 = io_brupdate_b1_mispredict_mask & rob_uop_3_19_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4215 = io_brupdate_b1_mispredict_mask & rob_uop_3_20_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4216 = io_brupdate_b1_mispredict_mask & rob_uop_3_21_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4217 = io_brupdate_b1_mispredict_mask & rob_uop_3_22_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4218 = io_brupdate_b1_mispredict_mask & rob_uop_3_23_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4219 = io_brupdate_b1_mispredict_mask & rob_uop_3_24_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4220 = io_brupdate_b1_mispredict_mask & rob_uop_3_25_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4221 = io_brupdate_b1_mispredict_mask & rob_uop_3_26_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4222 = io_brupdate_b1_mispredict_mask & rob_uop_3_27_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4223 = io_brupdate_b1_mispredict_mask & rob_uop_3_28_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4224 = io_brupdate_b1_mispredict_mask & rob_uop_3_29_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4225 = io_brupdate_b1_mispredict_mask & rob_uop_3_30_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4226 = io_brupdate_b1_mispredict_mask & rob_uop_3_31_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_4227 = ~(_io_flush_valid_output | exception_thrown) & rob_state != 2'h2;	// rob.scala:221:26, :236:31, :545:85, :573:36, :631:{9,26,47,60}
    _GEN_4228 =
      ~r_xcpt_val | io_lxcpt_bits_uop_rob_idx < r_xcpt_uop_rob_idx
      ^ io_lxcpt_bits_uop_rob_idx < rob_head_idx ^ r_xcpt_uop_rob_idx < rob_head_idx;	// Cat.scala:30:58, rob.scala:258:33, :259:29, :635:{13,25}, util.scala:363:{52,64,72,78}
    _GEN_4229 =
      ~r_xcpt_val
      & (enq_xcpts_0 | enq_xcpts_1 | enq_xcpts_2 | io_enq_valids_3
         & io_enq_uops_3_exception);	// rob.scala:258:33, :628:38, :635:13, :641:{30,51}
    idx = enq_xcpts_0 ? 2'h0 : enq_xcpts_1 ? 2'h1 : {1'h1, ~enq_xcpts_2};	// rob.scala:221:26, :540:33, :628:38, :642:37
    next_xcpt_uop_br_mask =
      _GEN_4227
        ? (io_lxcpt_valid
             ? (_GEN_4228 ? io_lxcpt_bits_uop_br_mask : r_xcpt_uop_br_mask)
             : _GEN_4229 ? _GEN_4230[idx] : r_xcpt_uop_br_mask)
        : r_xcpt_uop_br_mask;	// rob.scala:259:29, :625:17, :631:{47,76}, :632:27, :635:{25,93}, :637:33, :641:{30,56}, :642:37, :646:23
    if (reset) begin
      rob_state <= 2'h0;	// rob.scala:221:26
      rob_head <= 5'h0;	// rob.scala:224:29, :236:31, :268:25
      rob_head_lsb <= 2'h0;	// rob.scala:221:26, :225:29
      rob_tail <= 5'h0;	// rob.scala:228:29, :236:31, :268:25
      rob_tail_lsb <= 2'h0;	// rob.scala:221:26, :229:29
      rob_pnr <= 5'h0;	// rob.scala:232:29, :236:31, :268:25
      rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
      maybe_full <= 1'h0;	// rob.scala:239:29, :370:{23,59}, :372:26, :381:32
      r_xcpt_val <= 1'h0;	// rob.scala:258:33, :370:{23,59}, :372:26, :381:32
      rob_val_0 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_4 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_5 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_6 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_7 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_8 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_9 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_10 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_11 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_12 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_13 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_14 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_15 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_16 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_17 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_18 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_19 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_20 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_21 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_22 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_23 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_24 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_25 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_26 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_27 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_28 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_29 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_30 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_31 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_0 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_1 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_2 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_3 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_4 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_5 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_6 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_7 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_8 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_9 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_10 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_11 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_12 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_13 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_14 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_15 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_16 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_17 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_18 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_19 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_20 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_21 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_22 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_23 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_24 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_25 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_26 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_27 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_28 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_29 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_30 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_1_31 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_0 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_1 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_2 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_3 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_4 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_5 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_6 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_7 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_8 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_9 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_10 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_11 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_12 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_13 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_14 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_15 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_16 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_17 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_18 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_19 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_20 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_21 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_22 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_23 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_24 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_25 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_26 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_27 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_28 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_29 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_30 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_2_31 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_0 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_1 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_2 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_3 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_4 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_5 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_6 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_7 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_8 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_9 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_10 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_11 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_12 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_13 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_14 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_15 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_16 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_17 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_18 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_19 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_20 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_21 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_22 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_23 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_24 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_25 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_26 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_27 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_28 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_29 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_30 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      rob_val_3_31 <= 1'h0;	// rob.scala:307:32, :370:{23,59}, :372:26, :381:32
      r_partial_row <= 1'h0;	// rob.scala:370:{23,59}, :372:26, :381:32, :677:30
      pnr_maybe_at_tail <= 1'h0;	// rob.scala:370:{23,59}, :372:26, :381:32, :714:36
    end
    else begin
      automatic logic            _GEN_4232;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4233;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4234;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4235;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4236;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4237;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4238;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4239;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4240;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4241;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4242;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4243;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4244;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4245;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4246;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4247;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4248;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4249;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4250;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4251;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4252;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4253;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4254;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4255;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4256;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4257;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4258;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4259;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4260;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4261;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4262;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4263;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4264;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4265;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4266;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4267;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4268;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4269;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4270;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4271;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4272;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4273;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4274;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4275;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4276;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4277;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4278;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4279;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4280;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4281;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4282;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4283;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4284;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4285;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4286;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4287;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4288;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4289;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4290;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4291;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4292;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4293;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4294;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4295;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4296;	// rob.scala:476:25
      automatic logic            _GEN_4297;	// rob.scala:476:25
      automatic logic            _GEN_4298;	// rob.scala:476:25
      automatic logic            _GEN_4299;	// rob.scala:476:25
      automatic logic            _GEN_4300;	// rob.scala:476:25
      automatic logic            _GEN_4301;	// rob.scala:476:25
      automatic logic            _GEN_4302;	// rob.scala:476:25
      automatic logic            _GEN_4303;	// rob.scala:476:25
      automatic logic            _GEN_4304;	// rob.scala:476:25
      automatic logic            _GEN_4305;	// rob.scala:476:25
      automatic logic            _GEN_4306;	// rob.scala:476:25
      automatic logic            _GEN_4307;	// rob.scala:476:25
      automatic logic            _GEN_4308;	// rob.scala:476:25
      automatic logic            _GEN_4309;	// rob.scala:476:25
      automatic logic            _GEN_4310;	// rob.scala:476:25
      automatic logic            _GEN_4311;	// rob.scala:476:25
      automatic logic            _GEN_4312;	// rob.scala:476:25
      automatic logic            _GEN_4313;	// rob.scala:476:25
      automatic logic            _GEN_4314;	// rob.scala:476:25
      automatic logic            _GEN_4315;	// rob.scala:476:25
      automatic logic            _GEN_4316;	// rob.scala:476:25
      automatic logic            _GEN_4317;	// rob.scala:476:25
      automatic logic            _GEN_4318;	// rob.scala:476:25
      automatic logic            _GEN_4319;	// rob.scala:476:25
      automatic logic            _GEN_4320;	// rob.scala:476:25
      automatic logic            _GEN_4321;	// rob.scala:476:25
      automatic logic            _GEN_4322;	// rob.scala:476:25
      automatic logic            _GEN_4323;	// rob.scala:476:25
      automatic logic            _GEN_4324;	// rob.scala:476:25
      automatic logic            _GEN_4325;	// rob.scala:476:25
      automatic logic            _GEN_4326;	// rob.scala:476:25
      automatic logic            rob_pnr_unsafe_0;	// rob.scala:493:43
      automatic logic            _GEN_4327;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4328;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4329;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4330;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4331;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4332;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4333;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4334;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4335;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4336;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4337;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4338;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4339;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4340;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4341;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4342;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4343;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4344;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4345;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4346;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4347;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4348;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4349;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4350;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4351;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4352;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4353;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4354;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4355;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4356;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4357;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4358;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4359;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4360;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4361;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4362;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4363;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4364;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4365;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4366;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4367;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4368;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4369;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4370;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4371;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4372;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4373;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4374;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4375;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4376;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4377;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4378;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4379;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4380;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4381;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4382;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4383;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4384;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4385;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4386;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4387;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4388;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4389;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4390;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            rob_pnr_unsafe_1;	// rob.scala:493:43
      automatic logic            _GEN_4391;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4392;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4393;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4394;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4395;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4396;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4397;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4398;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4399;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4400;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4401;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4402;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4403;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4404;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4405;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4406;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4407;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4408;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4409;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4410;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4411;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4412;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4413;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4414;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4415;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4416;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4417;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4418;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4419;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4420;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4421;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4422;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4423;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4424;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4425;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4426;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4427;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4428;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4429;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4430;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4431;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4432;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4433;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4434;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4435;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4436;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4437;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4438;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4439;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4440;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4441;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4442;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4443;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4444;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4445;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4446;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4447;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4448;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4449;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4450;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4451;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4452;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4453;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4454;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            rob_pnr_unsafe_2;	// rob.scala:493:43
      automatic logic            _GEN_4455;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4456;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4457;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4458;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4459;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4460;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4461;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4462;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4463;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4464;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4465;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4466;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4467;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4468;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4469;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4470;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4471;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4472;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4473;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4474;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4475;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4476;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4477;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4478;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4479;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4480;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4481;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4482;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4483;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4484;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4485;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4486;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_4487;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4488;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4489;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4490;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4491;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4492;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4493;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4494;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4495;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4496;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4497;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4498;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4499;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4500;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4501;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4502;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4503;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4504;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4505;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4506;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4507;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4508;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4509;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4510;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4511;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4512;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4513;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4514;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4515;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4516;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4517;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_4518;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _do_inc_row_T_4;	// rob.scala:717:64
      automatic logic            do_inc_row;	// rob.scala:717:52
      automatic logic [3:0]      _GEN_4519;	// rob.scala:718:34
      automatic logic            _GEN_4520;	// rob.scala:755:68
      automatic logic            _GEN_4521;	// rob.scala:761:45
      automatic logic [1:0]      _GEN_4522;	// rob.scala:221:26, :819:22, :820:21
      automatic logic [3:0][1:0] _GEN_4523;	// Conditional.scala:37:30, :39:67, :40:58, rob.scala:221:26, :540:61, :804:19, :808:51, :819:22, :824:42
      _GEN_4232 = _GEN_148 | rob_val_0;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4233 = _GEN_150 | rob_val_1;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4234 = _GEN_152 | rob_val_2;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4235 = _GEN_154 | rob_val_3;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4236 = _GEN_156 | rob_val_4;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4237 = _GEN_158 | rob_val_5;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4238 = _GEN_160 | rob_val_6;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4239 = _GEN_162 | rob_val_7;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4240 = _GEN_164 | rob_val_8;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4241 = _GEN_166 | rob_val_9;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4242 = _GEN_168 | rob_val_10;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4243 = _GEN_170 | rob_val_11;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4244 = _GEN_172 | rob_val_12;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4245 = _GEN_174 | rob_val_13;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4246 = _GEN_176 | rob_val_14;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4247 = _GEN_178 | rob_val_15;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4248 = _GEN_180 | rob_val_16;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4249 = _GEN_182 | rob_val_17;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4250 = _GEN_184 | rob_val_18;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4251 = _GEN_186 | rob_val_19;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4252 = _GEN_188 | rob_val_20;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4253 = _GEN_190 | rob_val_21;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4254 = _GEN_192 | rob_val_22;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4255 = _GEN_194 | rob_val_23;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4256 = _GEN_196 | rob_val_24;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4257 = _GEN_198 | rob_val_25;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4258 = _GEN_200 | rob_val_26;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4259 = _GEN_202 | rob_val_27;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4260 = _GEN_204 | rob_val_28;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4261 = _GEN_206 | rob_val_29;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4262 = _GEN_208 | rob_val_30;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4263 = _GEN_209 | rob_val_31;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4264 = (|_GEN_1507) | _GEN_1445;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4265 = (|_GEN_1508) | _GEN_1447;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4266 = (|_GEN_1509) | _GEN_1449;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4267 = (|_GEN_1510) | _GEN_1451;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4268 = (|_GEN_1511) | _GEN_1453;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4269 = (|_GEN_1512) | _GEN_1455;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4270 = (|_GEN_1513) | _GEN_1457;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4271 = (|_GEN_1514) | _GEN_1459;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4272 = (|_GEN_1515) | _GEN_1461;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4273 = (|_GEN_1516) | _GEN_1463;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4274 = (|_GEN_1517) | _GEN_1465;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4275 = (|_GEN_1518) | _GEN_1467;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4276 = (|_GEN_1519) | _GEN_1469;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4277 = (|_GEN_1520) | _GEN_1471;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4278 = (|_GEN_1521) | _GEN_1473;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4279 = (|_GEN_1522) | _GEN_1475;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4280 = (|_GEN_1523) | _GEN_1477;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4281 = (|_GEN_1524) | _GEN_1479;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4282 = (|_GEN_1525) | _GEN_1481;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4283 = (|_GEN_1526) | _GEN_1483;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4284 = (|_GEN_1527) | _GEN_1485;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4285 = (|_GEN_1528) | _GEN_1487;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4286 = (|_GEN_1529) | _GEN_1489;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4287 = (|_GEN_1530) | _GEN_1491;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4288 = (|_GEN_1531) | _GEN_1493;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4289 = (|_GEN_1532) | _GEN_1495;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4290 = (|_GEN_1533) | _GEN_1497;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4291 = (|_GEN_1534) | _GEN_1499;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4292 = (|_GEN_1535) | _GEN_1501;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4293 = (|_GEN_1536) | _GEN_1503;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4294 = (|_GEN_1537) | _GEN_1505;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4295 = (|_GEN_1538) | _GEN_1506;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4296 = rob_head == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :476:25
      _GEN_4297 = rob_head == 5'h1;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4298 = rob_head == 5'h2;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4299 = rob_head == 5'h3;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4300 = rob_head == 5'h4;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4301 = rob_head == 5'h5;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4302 = rob_head == 5'h6;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4303 = rob_head == 5'h7;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4304 = rob_head == 5'h8;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4305 = rob_head == 5'h9;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4306 = rob_head == 5'hA;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4307 = rob_head == 5'hB;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4308 = rob_head == 5'hC;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4309 = rob_head == 5'hD;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4310 = rob_head == 5'hE;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4311 = rob_head == 5'hF;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4312 = rob_head == 5'h10;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4313 = rob_head == 5'h11;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4314 = rob_head == 5'h12;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4315 = rob_head == 5'h13;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4316 = rob_head == 5'h14;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4317 = rob_head == 5'h15;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4318 = rob_head == 5'h16;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4319 = rob_head == 5'h17;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4320 = rob_head == 5'h18;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4321 = rob_head == 5'h19;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4322 = rob_head == 5'h1A;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4323 = rob_head == 5'h1B;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4324 = rob_head == 5'h1C;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4325 = rob_head == 5'h1D;	// rob.scala:224:29, :324:31, :476:25
      _GEN_4326 = rob_head == 5'h1E;	// rob.scala:224:29, :324:31, :476:25
      rob_pnr_unsafe_0 = _GEN[rob_pnr] & (_GEN_15[rob_pnr] | _GEN_16[rob_pnr]);	// rob.scala:232:29, :324:31, :394:15, :398:49, :493:{43,67}
      _GEN_4327 = _GEN_1539 | rob_val_1_0;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4328 = _GEN_1540 | rob_val_1_1;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4329 = _GEN_1541 | rob_val_1_2;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4330 = _GEN_1542 | rob_val_1_3;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4331 = _GEN_1543 | rob_val_1_4;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4332 = _GEN_1544 | rob_val_1_5;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4333 = _GEN_1545 | rob_val_1_6;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4334 = _GEN_1546 | rob_val_1_7;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4335 = _GEN_1547 | rob_val_1_8;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4336 = _GEN_1548 | rob_val_1_9;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4337 = _GEN_1549 | rob_val_1_10;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4338 = _GEN_1550 | rob_val_1_11;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4339 = _GEN_1551 | rob_val_1_12;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4340 = _GEN_1552 | rob_val_1_13;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4341 = _GEN_1553 | rob_val_1_14;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4342 = _GEN_1554 | rob_val_1_15;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4343 = _GEN_1555 | rob_val_1_16;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4344 = _GEN_1556 | rob_val_1_17;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4345 = _GEN_1557 | rob_val_1_18;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4346 = _GEN_1558 | rob_val_1_19;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4347 = _GEN_1559 | rob_val_1_20;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4348 = _GEN_1560 | rob_val_1_21;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4349 = _GEN_1561 | rob_val_1_22;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4350 = _GEN_1562 | rob_val_1_23;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4351 = _GEN_1563 | rob_val_1_24;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4352 = _GEN_1564 | rob_val_1_25;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4353 = _GEN_1565 | rob_val_1_26;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4354 = _GEN_1566 | rob_val_1_27;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4355 = _GEN_1567 | rob_val_1_28;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4356 = _GEN_1568 | rob_val_1_29;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4357 = _GEN_1569 | rob_val_1_30;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4358 = _GEN_1570 | rob_val_1_31;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4359 = (|_GEN_2403) | _GEN_2371;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4360 = (|_GEN_2404) | _GEN_2372;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4361 = (|_GEN_2405) | _GEN_2373;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4362 = (|_GEN_2406) | _GEN_2374;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4363 = (|_GEN_2407) | _GEN_2375;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4364 = (|_GEN_2408) | _GEN_2376;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4365 = (|_GEN_2409) | _GEN_2377;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4366 = (|_GEN_2410) | _GEN_2378;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4367 = (|_GEN_2411) | _GEN_2379;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4368 = (|_GEN_2412) | _GEN_2380;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4369 = (|_GEN_2413) | _GEN_2381;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4370 = (|_GEN_2414) | _GEN_2382;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4371 = (|_GEN_2415) | _GEN_2383;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4372 = (|_GEN_2416) | _GEN_2384;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4373 = (|_GEN_2417) | _GEN_2385;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4374 = (|_GEN_2418) | _GEN_2386;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4375 = (|_GEN_2419) | _GEN_2387;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4376 = (|_GEN_2420) | _GEN_2388;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4377 = (|_GEN_2421) | _GEN_2389;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4378 = (|_GEN_2422) | _GEN_2390;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4379 = (|_GEN_2423) | _GEN_2391;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4380 = (|_GEN_2424) | _GEN_2392;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4381 = (|_GEN_2425) | _GEN_2393;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4382 = (|_GEN_2426) | _GEN_2394;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4383 = (|_GEN_2427) | _GEN_2395;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4384 = (|_GEN_2428) | _GEN_2396;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4385 = (|_GEN_2429) | _GEN_2397;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4386 = (|_GEN_2430) | _GEN_2398;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4387 = (|_GEN_2431) | _GEN_2399;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4388 = (|_GEN_2432) | _GEN_2400;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4389 = (|_GEN_2433) | _GEN_2401;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4390 = (|_GEN_2434) | _GEN_2402;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      rob_pnr_unsafe_1 = _GEN_34[rob_pnr] & (_GEN_50[rob_pnr] | _GEN_51[rob_pnr]);	// rob.scala:232:29, :324:31, :394:15, :398:49, :493:{43,67}
      _GEN_4391 = _GEN_2435 | rob_val_2_0;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4392 = _GEN_2436 | rob_val_2_1;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4393 = _GEN_2437 | rob_val_2_2;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4394 = _GEN_2438 | rob_val_2_3;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4395 = _GEN_2439 | rob_val_2_4;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4396 = _GEN_2440 | rob_val_2_5;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4397 = _GEN_2441 | rob_val_2_6;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4398 = _GEN_2442 | rob_val_2_7;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4399 = _GEN_2443 | rob_val_2_8;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4400 = _GEN_2444 | rob_val_2_9;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4401 = _GEN_2445 | rob_val_2_10;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4402 = _GEN_2446 | rob_val_2_11;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4403 = _GEN_2447 | rob_val_2_12;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4404 = _GEN_2448 | rob_val_2_13;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4405 = _GEN_2449 | rob_val_2_14;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4406 = _GEN_2450 | rob_val_2_15;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4407 = _GEN_2451 | rob_val_2_16;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4408 = _GEN_2452 | rob_val_2_17;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4409 = _GEN_2453 | rob_val_2_18;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4410 = _GEN_2454 | rob_val_2_19;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4411 = _GEN_2455 | rob_val_2_20;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4412 = _GEN_2456 | rob_val_2_21;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4413 = _GEN_2457 | rob_val_2_22;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4414 = _GEN_2458 | rob_val_2_23;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4415 = _GEN_2459 | rob_val_2_24;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4416 = _GEN_2460 | rob_val_2_25;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4417 = _GEN_2461 | rob_val_2_26;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4418 = _GEN_2462 | rob_val_2_27;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4419 = _GEN_2463 | rob_val_2_28;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4420 = _GEN_2464 | rob_val_2_29;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4421 = _GEN_2465 | rob_val_2_30;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4422 = _GEN_2466 | rob_val_2_31;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4423 = (|_GEN_3299) | _GEN_3267;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4424 = (|_GEN_3300) | _GEN_3268;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4425 = (|_GEN_3301) | _GEN_3269;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4426 = (|_GEN_3302) | _GEN_3270;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4427 = (|_GEN_3303) | _GEN_3271;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4428 = (|_GEN_3304) | _GEN_3272;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4429 = (|_GEN_3305) | _GEN_3273;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4430 = (|_GEN_3306) | _GEN_3274;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4431 = (|_GEN_3307) | _GEN_3275;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4432 = (|_GEN_3308) | _GEN_3276;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4433 = (|_GEN_3309) | _GEN_3277;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4434 = (|_GEN_3310) | _GEN_3278;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4435 = (|_GEN_3311) | _GEN_3279;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4436 = (|_GEN_3312) | _GEN_3280;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4437 = (|_GEN_3313) | _GEN_3281;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4438 = (|_GEN_3314) | _GEN_3282;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4439 = (|_GEN_3315) | _GEN_3283;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4440 = (|_GEN_3316) | _GEN_3284;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4441 = (|_GEN_3317) | _GEN_3285;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4442 = (|_GEN_3318) | _GEN_3286;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4443 = (|_GEN_3319) | _GEN_3287;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4444 = (|_GEN_3320) | _GEN_3288;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4445 = (|_GEN_3321) | _GEN_3289;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4446 = (|_GEN_3322) | _GEN_3290;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4447 = (|_GEN_3323) | _GEN_3291;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4448 = (|_GEN_3324) | _GEN_3292;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4449 = (|_GEN_3325) | _GEN_3293;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4450 = (|_GEN_3326) | _GEN_3294;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4451 = (|_GEN_3327) | _GEN_3295;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4452 = (|_GEN_3328) | _GEN_3296;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4453 = (|_GEN_3329) | _GEN_3297;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4454 = (|_GEN_3330) | _GEN_3298;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      rob_pnr_unsafe_2 = _GEN_69[rob_pnr] & (_GEN_85[rob_pnr] | _GEN_86[rob_pnr]);	// rob.scala:232:29, :324:31, :394:15, :398:49, :493:{43,67}
      _GEN_4455 = _GEN_3331 | rob_val_3_0;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4456 = _GEN_3332 | rob_val_3_1;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4457 = _GEN_3333 | rob_val_3_2;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4458 = _GEN_3334 | rob_val_3_3;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4459 = _GEN_3335 | rob_val_3_4;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4460 = _GEN_3336 | rob_val_3_5;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4461 = _GEN_3337 | rob_val_3_6;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4462 = _GEN_3338 | rob_val_3_7;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4463 = _GEN_3339 | rob_val_3_8;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4464 = _GEN_3340 | rob_val_3_9;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4465 = _GEN_3341 | rob_val_3_10;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4466 = _GEN_3342 | rob_val_3_11;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4467 = _GEN_3343 | rob_val_3_12;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4468 = _GEN_3344 | rob_val_3_13;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4469 = _GEN_3345 | rob_val_3_14;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4470 = _GEN_3346 | rob_val_3_15;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4471 = _GEN_3347 | rob_val_3_16;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4472 = _GEN_3348 | rob_val_3_17;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4473 = _GEN_3349 | rob_val_3_18;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4474 = _GEN_3350 | rob_val_3_19;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4475 = _GEN_3351 | rob_val_3_20;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4476 = _GEN_3352 | rob_val_3_21;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4477 = _GEN_3353 | rob_val_3_22;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4478 = _GEN_3354 | rob_val_3_23;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4479 = _GEN_3355 | rob_val_3_24;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4480 = _GEN_3356 | rob_val_3_25;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4481 = _GEN_3357 | rob_val_3_26;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4482 = _GEN_3358 | rob_val_3_27;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4483 = _GEN_3359 | rob_val_3_28;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4484 = _GEN_3360 | rob_val_3_29;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4485 = _GEN_3361 | rob_val_3_30;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4486 = _GEN_3362 | rob_val_3_31;	// rob.scala:307:32, :323:29, :324:31
      _GEN_4487 = (|_GEN_4195) | _GEN_4163;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4488 = (|_GEN_4196) | _GEN_4164;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4489 = (|_GEN_4197) | _GEN_4165;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4490 = (|_GEN_4198) | _GEN_4166;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4491 = (|_GEN_4199) | _GEN_4167;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4492 = (|_GEN_4200) | _GEN_4168;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4493 = (|_GEN_4201) | _GEN_4169;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4494 = (|_GEN_4202) | _GEN_4170;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4495 = (|_GEN_4203) | _GEN_4171;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4496 = (|_GEN_4204) | _GEN_4172;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4497 = (|_GEN_4205) | _GEN_4173;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4498 = (|_GEN_4206) | _GEN_4174;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4499 = (|_GEN_4207) | _GEN_4175;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4500 = (|_GEN_4208) | _GEN_4176;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4501 = (|_GEN_4209) | _GEN_4177;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4502 = (|_GEN_4210) | _GEN_4178;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4503 = (|_GEN_4211) | _GEN_4179;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4504 = (|_GEN_4212) | _GEN_4180;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4505 = (|_GEN_4213) | _GEN_4181;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4506 = (|_GEN_4214) | _GEN_4182;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4507 = (|_GEN_4215) | _GEN_4183;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4508 = (|_GEN_4216) | _GEN_4184;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4509 = (|_GEN_4217) | _GEN_4185;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4510 = (|_GEN_4218) | _GEN_4186;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4511 = (|_GEN_4219) | _GEN_4187;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4512 = (|_GEN_4220) | _GEN_4188;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4513 = (|_GEN_4221) | _GEN_4189;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4514 = (|_GEN_4222) | _GEN_4190;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4515 = (|_GEN_4223) | _GEN_4191;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4516 = (|_GEN_4224) | _GEN_4192;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4517 = (|_GEN_4225) | _GEN_4193;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_4518 = (|_GEN_4226) | _GEN_4194;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _do_inc_row_T_4 = rob_pnr != rob_tail;	// rob.scala:228:29, :232:29, :717:64
      do_inc_row =
        ~(rob_pnr_unsafe_0 | rob_pnr_unsafe_1 | rob_pnr_unsafe_2 | _GEN_104[rob_pnr]
          & (_GEN_120[rob_pnr] | _GEN_121[rob_pnr]))
        & (_do_inc_row_T_4 | full & ~pnr_maybe_at_tail);	// rob.scala:232:29, :324:31, :394:15, :398:49, :493:{43,67}, :714:36, :717:{23,47,52,64,77,86,89}, :787:39
      _GEN_4519 = {io_enq_valids_3, io_enq_valids_2, io_enq_valids_1, io_enq_valids_0};	// rob.scala:718:34
      _GEN_4520 = _io_commit_rollback_T_3 & rob_tail == rob_head & ~maybe_full;	// rob.scala:224:29, :228:29, :236:31, :239:29, :686:49, :755:{54,68}
      _GEN_4521 = (|_GEN_4519) & ~io_enq_partial_stall;	// rob.scala:718:{34,41}, :761:{45,48}
      _GEN_4522 = empty ? 2'h1 : rob_state;	// rob.scala:221:26, :540:33, :788:41, :819:22, :820:21
      _GEN_4523 =
        {{REG_2 ? 2'h2 : _GEN_4522},
         {_GEN_4522},
         {REG_1
            ? 2'h2
            : io_enq_valids_3 & io_enq_uops_3_is_unique | io_enq_valids_2
              & io_enq_uops_2_is_unique | io_enq_valids_1 & io_enq_uops_1_is_unique
              | io_enq_valids_0 & io_enq_uops_0_is_unique
                ? 2'h3
                : rob_state},
         {2'h1}};	// Conditional.scala:37:30, :39:67, :40:58, rob.scala:221:26, :236:31, :419:36, :540:{33,61}, :804:19, :808:{22,51}, :809:21, :812:{36,65}, :813:25, :819:22, :820:21, :824:{22,42}, :825:21, :826:29
      rob_state <= _GEN_4523[rob_state];	// Conditional.scala:37:30, :39:67, :40:58, rob.scala:221:26, :540:61, :804:19, :808:51, :819:22, :824:42
      if (finished_committing_row) begin	// rob.scala:685:59
        rob_head <= rob_head + 5'h1;	// rob.scala:224:29, :324:31, util.scala:203:14
        rob_head_lsb <= 2'h0;	// rob.scala:221:26, :225:29
      end
      else begin	// rob.scala:685:59
        automatic logic [2:0] _lo_T_12 =
          rob_head_vals_0
            ? 3'h0
            : rob_head_vals_1 ? 3'h1 : rob_head_vals_2 ? 3'h2 : {rob_head_vals_3, 2'h0};	// Mux.scala:47:69, rob.scala:174:10, :175:10, :221:26, :398:49
        rob_head_lsb <= {|(_lo_T_12[2:1]), _lo_T_12[2] | _lo_T_12[0]};	// Cat.scala:30:58, Mux.scala:47:69, OneHot.scala:30:18, :31:18, :32:{14,28}, rob.scala:225:29
      end
      if (_GEN_146) begin	// rob.scala:750:34
        rob_tail <= rob_tail - 5'h1;	// rob.scala:228:29, util.scala:220:14
        rob_tail_lsb <= 2'h3;	// rob.scala:229:29, :419:36
      end
      else if (_GEN_4520)	// rob.scala:755:68
        rob_tail_lsb <= rob_head_lsb;	// rob.scala:225:29, :229:29
      else begin	// rob.scala:755:68
        if (io_brupdate_b2_mispredict)
          rob_tail <= io_brupdate_b2_uop_rob_idx[6:2] + 5'h1;	// rob.scala:228:29, :236:31, :268:25, :324:31, util.scala:203:14
        else if (_GEN_4521)	// rob.scala:761:45
          rob_tail <= rob_tail + 5'h1;	// rob.scala:228:29, :324:31, util.scala:203:14
        if (io_brupdate_b2_mispredict | _GEN_4521)	// rob.scala:758:43, :760:18, :761:{45,71}, :763:18, :765:70
          rob_tail_lsb <= 2'h0;	// rob.scala:221:26, :229:29
        else if ((|_GEN_4519) & io_enq_partial_stall) begin	// rob.scala:718:{34,41}, :765:45
          automatic logic [2:0] _GEN_4524 =
            {io_enq_valids_2, io_enq_valids_1, io_enq_valids_0}
            | {io_enq_valids_3, io_enq_valids_2, io_enq_valids_1};	// util.scala:373:{29,45}
          automatic logic [1:0] _GEN_4525 =
            _GEN_4524[1:0] | {io_enq_valids_3, io_enq_valids_2};	// rob.scala:236:31, util.scala:373:{29,45}
          automatic logic [2:0] _lo_T_47;	// rob.scala:766:37
          _lo_T_47 = ~{_GEN_4524[2], _GEN_4525[1], _GEN_4525[0] | io_enq_valids_3};	// rob.scala:236:31, :419:36, :766:37, util.scala:373:{29,45}
          if (_lo_T_47[0])	// OneHot.scala:47:40, rob.scala:766:37
            rob_tail_lsb <= 2'h0;	// rob.scala:221:26, :229:29
          else if (_lo_T_47[1])	// OneHot.scala:47:40, rob.scala:766:37
            rob_tail_lsb <= 2'h1;	// rob.scala:229:29, :540:33
          else	// OneHot.scala:47:40
            rob_tail_lsb <= {1'h1, ~(_lo_T_47[2])};	// Mux.scala:47:69, OneHot.scala:47:40, rob.scala:229:29, :766:37
        end
      end
      if (empty & (|_GEN_4519)) begin	// rob.scala:718:{17,34,41}, :788:41
        rob_pnr <= rob_head;	// rob.scala:224:29, :232:29
        if (io_enq_valids_0)
          rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
        else if (io_enq_valids_1)
          rob_pnr_lsb <= 2'h1;	// rob.scala:233:29, :540:33
        else
          rob_pnr_lsb <= {1'h1, ~io_enq_valids_2};	// Mux.scala:47:69, rob.scala:233:29
      end
      else begin	// rob.scala:718:17
        automatic logic safe_to_inc;	// rob.scala:716:46
        safe_to_inc = _io_ready_T | (&rob_state);	// rob.scala:221:26, :716:{33,46,59}
        if (safe_to_inc & do_inc_row) begin	// rob.scala:716:46, :717:52, :725:30
          rob_pnr <= rob_pnr + 5'h1;	// rob.scala:232:29, :324:31, util.scala:203:14
          rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
        end
        else if (safe_to_inc & (_do_inc_row_T_4 | full & ~pnr_maybe_at_tail)) begin	// rob.scala:714:36, :716:46, :717:{64,89}, :728:{30,55,64}, :787:39
          if (rob_pnr_unsafe_0)	// rob.scala:493:43
            rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
          else if (rob_pnr_unsafe_1)	// rob.scala:493:43
            rob_pnr_lsb <= 2'h1;	// rob.scala:233:29, :540:33
          else	// rob.scala:493:43
            rob_pnr_lsb <= {1'h1, ~rob_pnr_unsafe_2};	// Mux.scala:47:69, rob.scala:233:29, :493:43
        end
        else if (safe_to_inc & ~full & ~empty) begin	// rob.scala:425:47, :716:46, :730:{39,42}, :787:39, :788:41
          automatic logic [2:0] _GEN_4526 =
            {rob_tail_vals_2, rob_tail_vals_1, rob_tail_vals_0}
            | {rob_tail_vals_3, rob_tail_vals_2, rob_tail_vals_1};	// rob.scala:324:31, util.scala:373:{29,45}
          automatic logic [1:0] _GEN_4527 =
            _GEN_4526[1:0] | {rob_tail_vals_3, rob_tail_vals_2};	// rob.scala:236:31, :324:31, util.scala:373:{29,45}
          automatic logic [2:0] _lo_T_31;	// rob.scala:731:60
          _lo_T_31 =
            {rob_pnr_unsafe_2, rob_pnr_unsafe_1, rob_pnr_unsafe_0}
            | ~{_GEN_4526[2], _GEN_4527[1], _GEN_4527[0] | rob_tail_vals_3};	// rob.scala:236:31, :324:31, :419:36, :493:43, :731:{53,60,62}, util.scala:373:{29,45}
          if (_lo_T_31[0])	// OneHot.scala:47:40, rob.scala:731:60
            rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
          else if (_lo_T_31[1])	// OneHot.scala:47:40, rob.scala:731:60
            rob_pnr_lsb <= 2'h1;	// rob.scala:233:29, :540:33
          else	// OneHot.scala:47:40
            rob_pnr_lsb <= {1'h1, ~(_lo_T_31[2])};	// Mux.scala:47:69, OneHot.scala:47:40, rob.scala:233:29, :731:60
        end
        else if (full & pnr_maybe_at_tail)	// rob.scala:714:36, :732:23, :787:39
          rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
      end
      maybe_full <=
        ~rob_deq
        & (~(_GEN_146 | _GEN_4520 | io_brupdate_b2_mispredict) & _GEN_4521 | maybe_full)
        | (|io_brupdate_b1_mispredict_mask);	// rob.scala:239:29, :688:34, :736:26, :750:{34,76}, :754:13, :755:{68,84}, :758:43, :761:{45,71}, :786:{26,38,53,87}
      r_xcpt_val <=
        ~(_io_flush_valid_output
          | (|(io_brupdate_b1_mispredict_mask & next_xcpt_uop_br_mask)))
        & (_GEN_4227
             ? (io_lxcpt_valid ? _GEN_4228 | r_xcpt_val : _GEN_4229 | r_xcpt_val)
             : r_xcpt_val);	// rob.scala:258:33, :573:36, :625:17, :631:{47,76}, :632:27, :635:{25,93}, :636:33, :641:{30,56}, :645:23, :654:{24,73}, :655:16, util.scala:118:{51,59}
      if (will_commit_0) begin	// rob.scala:547:70
        rob_val_0 <= ~(_GEN_4296 | _GEN_4264) & _GEN_4232;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1 <= ~(_GEN_4297 | _GEN_4265) & _GEN_4233;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2 <= ~(_GEN_4298 | _GEN_4266) & _GEN_4234;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3 <= ~(_GEN_4299 | _GEN_4267) & _GEN_4235;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_4 <= ~(_GEN_4300 | _GEN_4268) & _GEN_4236;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_5 <= ~(_GEN_4301 | _GEN_4269) & _GEN_4237;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_6 <= ~(_GEN_4302 | _GEN_4270) & _GEN_4238;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_7 <= ~(_GEN_4303 | _GEN_4271) & _GEN_4239;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_8 <= ~(_GEN_4304 | _GEN_4272) & _GEN_4240;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_9 <= ~(_GEN_4305 | _GEN_4273) & _GEN_4241;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_10 <= ~(_GEN_4306 | _GEN_4274) & _GEN_4242;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_11 <= ~(_GEN_4307 | _GEN_4275) & _GEN_4243;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_12 <= ~(_GEN_4308 | _GEN_4276) & _GEN_4244;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_13 <= ~(_GEN_4309 | _GEN_4277) & _GEN_4245;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_14 <= ~(_GEN_4310 | _GEN_4278) & _GEN_4246;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_15 <= ~(_GEN_4311 | _GEN_4279) & _GEN_4247;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_16 <= ~(_GEN_4312 | _GEN_4280) & _GEN_4248;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_17 <= ~(_GEN_4313 | _GEN_4281) & _GEN_4249;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_18 <= ~(_GEN_4314 | _GEN_4282) & _GEN_4250;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_19 <= ~(_GEN_4315 | _GEN_4283) & _GEN_4251;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_20 <= ~(_GEN_4316 | _GEN_4284) & _GEN_4252;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_21 <= ~(_GEN_4317 | _GEN_4285) & _GEN_4253;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_22 <= ~(_GEN_4318 | _GEN_4286) & _GEN_4254;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_23 <= ~(_GEN_4319 | _GEN_4287) & _GEN_4255;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_24 <= ~(_GEN_4320 | _GEN_4288) & _GEN_4256;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_25 <= ~(_GEN_4321 | _GEN_4289) & _GEN_4257;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_26 <= ~(_GEN_4322 | _GEN_4290) & _GEN_4258;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_27 <= ~(_GEN_4323 | _GEN_4291) & _GEN_4259;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_28 <= ~(_GEN_4324 | _GEN_4292) & _GEN_4260;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_29 <= ~(_GEN_4325 | _GEN_4293) & _GEN_4261;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_30 <= ~(_GEN_4326 | _GEN_4294) & _GEN_4262;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_31 <= ~((&rob_head) | _GEN_4295) & _GEN_4263;	// rob.scala:224:29, :307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
      end
      else begin	// rob.scala:547:70
        rob_val_0 <= ~_GEN_4264 & _GEN_4232;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1 <= ~_GEN_4265 & _GEN_4233;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2 <= ~_GEN_4266 & _GEN_4234;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3 <= ~_GEN_4267 & _GEN_4235;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_4 <= ~_GEN_4268 & _GEN_4236;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_5 <= ~_GEN_4269 & _GEN_4237;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_6 <= ~_GEN_4270 & _GEN_4238;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_7 <= ~_GEN_4271 & _GEN_4239;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_8 <= ~_GEN_4272 & _GEN_4240;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_9 <= ~_GEN_4273 & _GEN_4241;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_10 <= ~_GEN_4274 & _GEN_4242;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_11 <= ~_GEN_4275 & _GEN_4243;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_12 <= ~_GEN_4276 & _GEN_4244;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_13 <= ~_GEN_4277 & _GEN_4245;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_14 <= ~_GEN_4278 & _GEN_4246;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_15 <= ~_GEN_4279 & _GEN_4247;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_16 <= ~_GEN_4280 & _GEN_4248;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_17 <= ~_GEN_4281 & _GEN_4249;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_18 <= ~_GEN_4282 & _GEN_4250;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_19 <= ~_GEN_4283 & _GEN_4251;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_20 <= ~_GEN_4284 & _GEN_4252;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_21 <= ~_GEN_4285 & _GEN_4253;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_22 <= ~_GEN_4286 & _GEN_4254;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_23 <= ~_GEN_4287 & _GEN_4255;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_24 <= ~_GEN_4288 & _GEN_4256;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_25 <= ~_GEN_4289 & _GEN_4257;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_26 <= ~_GEN_4290 & _GEN_4258;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_27 <= ~_GEN_4291 & _GEN_4259;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_28 <= ~_GEN_4292 & _GEN_4260;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_29 <= ~_GEN_4293 & _GEN_4261;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_30 <= ~_GEN_4294 & _GEN_4262;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_31 <= ~_GEN_4295 & _GEN_4263;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
      end
      if (will_commit_1) begin	// rob.scala:547:70
        rob_val_1_0 <= ~(_GEN_4296 | _GEN_4359) & _GEN_4327;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_1 <= ~(_GEN_4297 | _GEN_4360) & _GEN_4328;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_2 <= ~(_GEN_4298 | _GEN_4361) & _GEN_4329;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_3 <= ~(_GEN_4299 | _GEN_4362) & _GEN_4330;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_4 <= ~(_GEN_4300 | _GEN_4363) & _GEN_4331;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_5 <= ~(_GEN_4301 | _GEN_4364) & _GEN_4332;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_6 <= ~(_GEN_4302 | _GEN_4365) & _GEN_4333;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_7 <= ~(_GEN_4303 | _GEN_4366) & _GEN_4334;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_8 <= ~(_GEN_4304 | _GEN_4367) & _GEN_4335;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_9 <= ~(_GEN_4305 | _GEN_4368) & _GEN_4336;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_10 <= ~(_GEN_4306 | _GEN_4369) & _GEN_4337;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_11 <= ~(_GEN_4307 | _GEN_4370) & _GEN_4338;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_12 <= ~(_GEN_4308 | _GEN_4371) & _GEN_4339;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_13 <= ~(_GEN_4309 | _GEN_4372) & _GEN_4340;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_14 <= ~(_GEN_4310 | _GEN_4373) & _GEN_4341;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_15 <= ~(_GEN_4311 | _GEN_4374) & _GEN_4342;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_16 <= ~(_GEN_4312 | _GEN_4375) & _GEN_4343;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_17 <= ~(_GEN_4313 | _GEN_4376) & _GEN_4344;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_18 <= ~(_GEN_4314 | _GEN_4377) & _GEN_4345;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_19 <= ~(_GEN_4315 | _GEN_4378) & _GEN_4346;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_20 <= ~(_GEN_4316 | _GEN_4379) & _GEN_4347;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_21 <= ~(_GEN_4317 | _GEN_4380) & _GEN_4348;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_22 <= ~(_GEN_4318 | _GEN_4381) & _GEN_4349;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_23 <= ~(_GEN_4319 | _GEN_4382) & _GEN_4350;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_24 <= ~(_GEN_4320 | _GEN_4383) & _GEN_4351;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_25 <= ~(_GEN_4321 | _GEN_4384) & _GEN_4352;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_26 <= ~(_GEN_4322 | _GEN_4385) & _GEN_4353;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_27 <= ~(_GEN_4323 | _GEN_4386) & _GEN_4354;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_28 <= ~(_GEN_4324 | _GEN_4387) & _GEN_4355;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_29 <= ~(_GEN_4325 | _GEN_4388) & _GEN_4356;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_30 <= ~(_GEN_4326 | _GEN_4389) & _GEN_4357;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_31 <= ~((&rob_head) | _GEN_4390) & _GEN_4358;	// rob.scala:224:29, :307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
      end
      else begin	// rob.scala:547:70
        rob_val_1_0 <= ~_GEN_4359 & _GEN_4327;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_1 <= ~_GEN_4360 & _GEN_4328;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_2 <= ~_GEN_4361 & _GEN_4329;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_3 <= ~_GEN_4362 & _GEN_4330;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_4 <= ~_GEN_4363 & _GEN_4331;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_5 <= ~_GEN_4364 & _GEN_4332;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_6 <= ~_GEN_4365 & _GEN_4333;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_7 <= ~_GEN_4366 & _GEN_4334;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_8 <= ~_GEN_4367 & _GEN_4335;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_9 <= ~_GEN_4368 & _GEN_4336;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_10 <= ~_GEN_4369 & _GEN_4337;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_11 <= ~_GEN_4370 & _GEN_4338;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_12 <= ~_GEN_4371 & _GEN_4339;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_13 <= ~_GEN_4372 & _GEN_4340;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_14 <= ~_GEN_4373 & _GEN_4341;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_15 <= ~_GEN_4374 & _GEN_4342;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_16 <= ~_GEN_4375 & _GEN_4343;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_17 <= ~_GEN_4376 & _GEN_4344;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_18 <= ~_GEN_4377 & _GEN_4345;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_19 <= ~_GEN_4378 & _GEN_4346;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_20 <= ~_GEN_4379 & _GEN_4347;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_21 <= ~_GEN_4380 & _GEN_4348;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_22 <= ~_GEN_4381 & _GEN_4349;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_23 <= ~_GEN_4382 & _GEN_4350;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_24 <= ~_GEN_4383 & _GEN_4351;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_25 <= ~_GEN_4384 & _GEN_4352;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_26 <= ~_GEN_4385 & _GEN_4353;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_27 <= ~_GEN_4386 & _GEN_4354;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_28 <= ~_GEN_4387 & _GEN_4355;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_29 <= ~_GEN_4388 & _GEN_4356;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_30 <= ~_GEN_4389 & _GEN_4357;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_31 <= ~_GEN_4390 & _GEN_4358;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
      end
      if (will_commit_2) begin	// rob.scala:547:70
        rob_val_2_0 <= ~(_GEN_4296 | _GEN_4423) & _GEN_4391;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_1 <= ~(_GEN_4297 | _GEN_4424) & _GEN_4392;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_2 <= ~(_GEN_4298 | _GEN_4425) & _GEN_4393;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_3 <= ~(_GEN_4299 | _GEN_4426) & _GEN_4394;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_4 <= ~(_GEN_4300 | _GEN_4427) & _GEN_4395;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_5 <= ~(_GEN_4301 | _GEN_4428) & _GEN_4396;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_6 <= ~(_GEN_4302 | _GEN_4429) & _GEN_4397;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_7 <= ~(_GEN_4303 | _GEN_4430) & _GEN_4398;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_8 <= ~(_GEN_4304 | _GEN_4431) & _GEN_4399;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_9 <= ~(_GEN_4305 | _GEN_4432) & _GEN_4400;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_10 <= ~(_GEN_4306 | _GEN_4433) & _GEN_4401;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_11 <= ~(_GEN_4307 | _GEN_4434) & _GEN_4402;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_12 <= ~(_GEN_4308 | _GEN_4435) & _GEN_4403;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_13 <= ~(_GEN_4309 | _GEN_4436) & _GEN_4404;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_14 <= ~(_GEN_4310 | _GEN_4437) & _GEN_4405;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_15 <= ~(_GEN_4311 | _GEN_4438) & _GEN_4406;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_16 <= ~(_GEN_4312 | _GEN_4439) & _GEN_4407;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_17 <= ~(_GEN_4313 | _GEN_4440) & _GEN_4408;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_18 <= ~(_GEN_4314 | _GEN_4441) & _GEN_4409;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_19 <= ~(_GEN_4315 | _GEN_4442) & _GEN_4410;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_20 <= ~(_GEN_4316 | _GEN_4443) & _GEN_4411;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_21 <= ~(_GEN_4317 | _GEN_4444) & _GEN_4412;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_22 <= ~(_GEN_4318 | _GEN_4445) & _GEN_4413;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_23 <= ~(_GEN_4319 | _GEN_4446) & _GEN_4414;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_24 <= ~(_GEN_4320 | _GEN_4447) & _GEN_4415;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_25 <= ~(_GEN_4321 | _GEN_4448) & _GEN_4416;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_26 <= ~(_GEN_4322 | _GEN_4449) & _GEN_4417;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_27 <= ~(_GEN_4323 | _GEN_4450) & _GEN_4418;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_28 <= ~(_GEN_4324 | _GEN_4451) & _GEN_4419;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_29 <= ~(_GEN_4325 | _GEN_4452) & _GEN_4420;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_30 <= ~(_GEN_4326 | _GEN_4453) & _GEN_4421;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_31 <= ~((&rob_head) | _GEN_4454) & _GEN_4422;	// rob.scala:224:29, :307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
      end
      else begin	// rob.scala:547:70
        rob_val_2_0 <= ~_GEN_4423 & _GEN_4391;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_1 <= ~_GEN_4424 & _GEN_4392;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_2 <= ~_GEN_4425 & _GEN_4393;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_3 <= ~_GEN_4426 & _GEN_4394;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_4 <= ~_GEN_4427 & _GEN_4395;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_5 <= ~_GEN_4428 & _GEN_4396;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_6 <= ~_GEN_4429 & _GEN_4397;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_7 <= ~_GEN_4430 & _GEN_4398;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_8 <= ~_GEN_4431 & _GEN_4399;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_9 <= ~_GEN_4432 & _GEN_4400;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_10 <= ~_GEN_4433 & _GEN_4401;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_11 <= ~_GEN_4434 & _GEN_4402;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_12 <= ~_GEN_4435 & _GEN_4403;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_13 <= ~_GEN_4436 & _GEN_4404;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_14 <= ~_GEN_4437 & _GEN_4405;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_15 <= ~_GEN_4438 & _GEN_4406;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_16 <= ~_GEN_4439 & _GEN_4407;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_17 <= ~_GEN_4440 & _GEN_4408;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_18 <= ~_GEN_4441 & _GEN_4409;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_19 <= ~_GEN_4442 & _GEN_4410;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_20 <= ~_GEN_4443 & _GEN_4411;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_21 <= ~_GEN_4444 & _GEN_4412;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_22 <= ~_GEN_4445 & _GEN_4413;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_23 <= ~_GEN_4446 & _GEN_4414;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_24 <= ~_GEN_4447 & _GEN_4415;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_25 <= ~_GEN_4448 & _GEN_4416;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_26 <= ~_GEN_4449 & _GEN_4417;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_27 <= ~_GEN_4450 & _GEN_4418;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_28 <= ~_GEN_4451 & _GEN_4419;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_29 <= ~_GEN_4452 & _GEN_4420;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_30 <= ~_GEN_4453 & _GEN_4421;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_31 <= ~_GEN_4454 & _GEN_4422;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
      end
      if (will_commit_3) begin	// rob.scala:547:70
        rob_val_3_0 <= ~(_GEN_4296 | _GEN_4487) & _GEN_4455;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_1 <= ~(_GEN_4297 | _GEN_4488) & _GEN_4456;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_2 <= ~(_GEN_4298 | _GEN_4489) & _GEN_4457;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_3 <= ~(_GEN_4299 | _GEN_4490) & _GEN_4458;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_4 <= ~(_GEN_4300 | _GEN_4491) & _GEN_4459;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_5 <= ~(_GEN_4301 | _GEN_4492) & _GEN_4460;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_6 <= ~(_GEN_4302 | _GEN_4493) & _GEN_4461;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_7 <= ~(_GEN_4303 | _GEN_4494) & _GEN_4462;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_8 <= ~(_GEN_4304 | _GEN_4495) & _GEN_4463;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_9 <= ~(_GEN_4305 | _GEN_4496) & _GEN_4464;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_10 <= ~(_GEN_4306 | _GEN_4497) & _GEN_4465;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_11 <= ~(_GEN_4307 | _GEN_4498) & _GEN_4466;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_12 <= ~(_GEN_4308 | _GEN_4499) & _GEN_4467;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_13 <= ~(_GEN_4309 | _GEN_4500) & _GEN_4468;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_14 <= ~(_GEN_4310 | _GEN_4501) & _GEN_4469;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_15 <= ~(_GEN_4311 | _GEN_4502) & _GEN_4470;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_16 <= ~(_GEN_4312 | _GEN_4503) & _GEN_4471;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_17 <= ~(_GEN_4313 | _GEN_4504) & _GEN_4472;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_18 <= ~(_GEN_4314 | _GEN_4505) & _GEN_4473;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_19 <= ~(_GEN_4315 | _GEN_4506) & _GEN_4474;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_20 <= ~(_GEN_4316 | _GEN_4507) & _GEN_4475;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_21 <= ~(_GEN_4317 | _GEN_4508) & _GEN_4476;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_22 <= ~(_GEN_4318 | _GEN_4509) & _GEN_4477;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_23 <= ~(_GEN_4319 | _GEN_4510) & _GEN_4478;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_24 <= ~(_GEN_4320 | _GEN_4511) & _GEN_4479;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_25 <= ~(_GEN_4321 | _GEN_4512) & _GEN_4480;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_26 <= ~(_GEN_4322 | _GEN_4513) & _GEN_4481;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_27 <= ~(_GEN_4323 | _GEN_4514) & _GEN_4482;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_28 <= ~(_GEN_4324 | _GEN_4515) & _GEN_4483;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_29 <= ~(_GEN_4325 | _GEN_4516) & _GEN_4484;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_30 <= ~(_GEN_4326 | _GEN_4517) & _GEN_4485;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3_31 <= ~((&rob_head) | _GEN_4518) & _GEN_4486;	// rob.scala:224:29, :307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
      end
      else begin	// rob.scala:547:70
        rob_val_3_0 <= ~_GEN_4487 & _GEN_4455;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_1 <= ~_GEN_4488 & _GEN_4456;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_2 <= ~_GEN_4489 & _GEN_4457;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_3 <= ~_GEN_4490 & _GEN_4458;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_4 <= ~_GEN_4491 & _GEN_4459;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_5 <= ~_GEN_4492 & _GEN_4460;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_6 <= ~_GEN_4493 & _GEN_4461;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_7 <= ~_GEN_4494 & _GEN_4462;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_8 <= ~_GEN_4495 & _GEN_4463;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_9 <= ~_GEN_4496 & _GEN_4464;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_10 <= ~_GEN_4497 & _GEN_4465;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_11 <= ~_GEN_4498 & _GEN_4466;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_12 <= ~_GEN_4499 & _GEN_4467;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_13 <= ~_GEN_4500 & _GEN_4468;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_14 <= ~_GEN_4501 & _GEN_4469;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_15 <= ~_GEN_4502 & _GEN_4470;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_16 <= ~_GEN_4503 & _GEN_4471;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_17 <= ~_GEN_4504 & _GEN_4472;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_18 <= ~_GEN_4505 & _GEN_4473;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_19 <= ~_GEN_4506 & _GEN_4474;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_20 <= ~_GEN_4507 & _GEN_4475;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_21 <= ~_GEN_4508 & _GEN_4476;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_22 <= ~_GEN_4509 & _GEN_4477;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_23 <= ~_GEN_4510 & _GEN_4478;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_24 <= ~_GEN_4511 & _GEN_4479;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_25 <= ~_GEN_4512 & _GEN_4480;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_26 <= ~_GEN_4513 & _GEN_4481;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_27 <= ~_GEN_4514 & _GEN_4482;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_28 <= ~_GEN_4515 & _GEN_4483;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_29 <= ~_GEN_4516 & _GEN_4484;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_30 <= ~_GEN_4517 & _GEN_4485;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3_31 <= ~_GEN_4518 & _GEN_4486;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
      end
      if (io_enq_valids_0 | io_enq_valids_1 | io_enq_valids_2 | io_enq_valids_3)	// rob.scala:679:31
        r_partial_row <= io_enq_partial_stall;	// rob.scala:677:30
      pnr_maybe_at_tail <= ~rob_deq & (do_inc_row | pnr_maybe_at_tail);	// rob.scala:688:34, :714:36, :717:52, :736:{26,35,50}, :750:76, :754:13
    end
    r_xcpt_uop_br_mask <= next_xcpt_uop_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:259:29, :625:17, :631:76, :632:27, util.scala:85:{25,27}
    if (_GEN_4227) begin	// rob.scala:631:47
      if (io_lxcpt_valid) begin
        if (_GEN_4228) begin	// rob.scala:635:25
          r_xcpt_uop_rob_idx <= io_lxcpt_bits_uop_rob_idx;	// rob.scala:259:29
          r_xcpt_uop_exc_cause <= {59'h0, io_lxcpt_bits_cause};	// rob.scala:259:29, :556:50, :638:33
          r_xcpt_badvaddr <= io_lxcpt_bits_badvaddr;	// rob.scala:260:29
        end
      end
      else if (_GEN_4229) begin	// rob.scala:641:30
        automatic logic [3:0][6:0]  _GEN_4528 =
          {{io_enq_uops_3_rob_idx},
           {io_enq_uops_2_rob_idx},
           {io_enq_uops_1_rob_idx},
           {io_enq_uops_0_rob_idx}};	// rob.scala:646:23
        automatic logic [3:0][63:0] _GEN_4529 =
          {{io_enq_uops_3_exc_cause},
           {io_enq_uops_2_exc_cause},
           {io_enq_uops_1_exc_cause},
           {io_enq_uops_0_exc_cause}};	// rob.scala:646:23
        automatic logic [3:0][5:0]  _GEN_4530 =
          {{io_enq_uops_3_pc_lob},
           {io_enq_uops_2_pc_lob},
           {io_enq_uops_1_pc_lob},
           {io_enq_uops_0_pc_lob}};	// rob.scala:646:23
        r_xcpt_uop_rob_idx <= _GEN_4528[idx];	// rob.scala:259:29, :642:37, :646:23
        r_xcpt_uop_exc_cause <= _GEN_4529[idx];	// rob.scala:259:29, :642:37, :646:23
        r_xcpt_badvaddr <= {io_xcpt_fetch_pc[39:6], _GEN_4530[idx]};	// rob.scala:260:29, :642:37, :646:23, :647:76
      end
    end
    rob_bsy_0 <= ~_GEN_1351 & (_GEN_12 ? ~_GEN_1288 & _GEN_1099 : ~_GEN_1225 & _GEN_1099);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1 <= ~_GEN_1353 & (_GEN_12 ? ~_GEN_1290 & _GEN_1102 : ~_GEN_1227 & _GEN_1102);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2 <= ~_GEN_1355 & (_GEN_12 ? ~_GEN_1292 & _GEN_1105 : ~_GEN_1229 & _GEN_1105);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3 <= ~_GEN_1357 & (_GEN_12 ? ~_GEN_1294 & _GEN_1108 : ~_GEN_1231 & _GEN_1108);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_4 <= ~_GEN_1359 & (_GEN_12 ? ~_GEN_1296 & _GEN_1111 : ~_GEN_1233 & _GEN_1111);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_5 <= ~_GEN_1361 & (_GEN_12 ? ~_GEN_1298 & _GEN_1114 : ~_GEN_1235 & _GEN_1114);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_6 <= ~_GEN_1363 & (_GEN_12 ? ~_GEN_1300 & _GEN_1117 : ~_GEN_1237 & _GEN_1117);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_7 <= ~_GEN_1365 & (_GEN_12 ? ~_GEN_1302 & _GEN_1120 : ~_GEN_1239 & _GEN_1120);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_8 <= ~_GEN_1367 & (_GEN_12 ? ~_GEN_1304 & _GEN_1123 : ~_GEN_1241 & _GEN_1123);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_9 <= ~_GEN_1369 & (_GEN_12 ? ~_GEN_1306 & _GEN_1126 : ~_GEN_1243 & _GEN_1126);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_10 <=
      ~_GEN_1371 & (_GEN_12 ? ~_GEN_1308 & _GEN_1129 : ~_GEN_1245 & _GEN_1129);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_11 <=
      ~_GEN_1373 & (_GEN_12 ? ~_GEN_1310 & _GEN_1132 : ~_GEN_1247 & _GEN_1132);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_12 <=
      ~_GEN_1375 & (_GEN_12 ? ~_GEN_1312 & _GEN_1135 : ~_GEN_1249 & _GEN_1135);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_13 <=
      ~_GEN_1377 & (_GEN_12 ? ~_GEN_1314 & _GEN_1138 : ~_GEN_1251 & _GEN_1138);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_14 <=
      ~_GEN_1379 & (_GEN_12 ? ~_GEN_1316 & _GEN_1141 : ~_GEN_1253 & _GEN_1141);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_15 <=
      ~_GEN_1381 & (_GEN_12 ? ~_GEN_1318 & _GEN_1144 : ~_GEN_1255 & _GEN_1144);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_16 <=
      ~_GEN_1383 & (_GEN_12 ? ~_GEN_1320 & _GEN_1147 : ~_GEN_1257 & _GEN_1147);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_17 <=
      ~_GEN_1385 & (_GEN_12 ? ~_GEN_1322 & _GEN_1150 : ~_GEN_1259 & _GEN_1150);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_18 <=
      ~_GEN_1387 & (_GEN_12 ? ~_GEN_1324 & _GEN_1153 : ~_GEN_1261 & _GEN_1153);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_19 <=
      ~_GEN_1389 & (_GEN_12 ? ~_GEN_1326 & _GEN_1156 : ~_GEN_1263 & _GEN_1156);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_20 <=
      ~_GEN_1391 & (_GEN_12 ? ~_GEN_1328 & _GEN_1159 : ~_GEN_1265 & _GEN_1159);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_21 <=
      ~_GEN_1393 & (_GEN_12 ? ~_GEN_1330 & _GEN_1162 : ~_GEN_1267 & _GEN_1162);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_22 <=
      ~_GEN_1395 & (_GEN_12 ? ~_GEN_1332 & _GEN_1165 : ~_GEN_1269 & _GEN_1165);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_23 <=
      ~_GEN_1397 & (_GEN_12 ? ~_GEN_1334 & _GEN_1168 : ~_GEN_1271 & _GEN_1168);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_24 <=
      ~_GEN_1399 & (_GEN_12 ? ~_GEN_1336 & _GEN_1171 : ~_GEN_1273 & _GEN_1171);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_25 <=
      ~_GEN_1401 & (_GEN_12 ? ~_GEN_1338 & _GEN_1174 : ~_GEN_1275 & _GEN_1174);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_26 <=
      ~_GEN_1403 & (_GEN_12 ? ~_GEN_1340 & _GEN_1177 : ~_GEN_1277 & _GEN_1177);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_27 <=
      ~_GEN_1405 & (_GEN_12 ? ~_GEN_1342 & _GEN_1180 : ~_GEN_1279 & _GEN_1180);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_28 <=
      ~_GEN_1407 & (_GEN_12 ? ~_GEN_1344 & _GEN_1183 : ~_GEN_1281 & _GEN_1183);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_29 <=
      ~_GEN_1409 & (_GEN_12 ? ~_GEN_1346 & _GEN_1186 : ~_GEN_1283 & _GEN_1186);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_30 <=
      ~_GEN_1411 & (_GEN_12 ? ~_GEN_1348 & _GEN_1189 : ~_GEN_1285 & _GEN_1189);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_31 <=
      ~_GEN_1412 & (_GEN_12 ? ~_GEN_1349 & _GEN_1191 : ~_GEN_1286 & _GEN_1191);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_unsafe_0 <=
      ~_GEN_1351 & (_GEN_12 ? ~_GEN_1288 & _GEN_1192 : ~_GEN_1225 & _GEN_1192);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1 <=
      ~_GEN_1353 & (_GEN_12 ? ~_GEN_1290 & _GEN_1193 : ~_GEN_1227 & _GEN_1193);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2 <=
      ~_GEN_1355 & (_GEN_12 ? ~_GEN_1292 & _GEN_1194 : ~_GEN_1229 & _GEN_1194);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3 <=
      ~_GEN_1357 & (_GEN_12 ? ~_GEN_1294 & _GEN_1195 : ~_GEN_1231 & _GEN_1195);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_4 <=
      ~_GEN_1359 & (_GEN_12 ? ~_GEN_1296 & _GEN_1196 : ~_GEN_1233 & _GEN_1196);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_5 <=
      ~_GEN_1361 & (_GEN_12 ? ~_GEN_1298 & _GEN_1197 : ~_GEN_1235 & _GEN_1197);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_6 <=
      ~_GEN_1363 & (_GEN_12 ? ~_GEN_1300 & _GEN_1198 : ~_GEN_1237 & _GEN_1198);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_7 <=
      ~_GEN_1365 & (_GEN_12 ? ~_GEN_1302 & _GEN_1199 : ~_GEN_1239 & _GEN_1199);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_8 <=
      ~_GEN_1367 & (_GEN_12 ? ~_GEN_1304 & _GEN_1200 : ~_GEN_1241 & _GEN_1200);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_9 <=
      ~_GEN_1369 & (_GEN_12 ? ~_GEN_1306 & _GEN_1201 : ~_GEN_1243 & _GEN_1201);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_10 <=
      ~_GEN_1371 & (_GEN_12 ? ~_GEN_1308 & _GEN_1202 : ~_GEN_1245 & _GEN_1202);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_11 <=
      ~_GEN_1373 & (_GEN_12 ? ~_GEN_1310 & _GEN_1203 : ~_GEN_1247 & _GEN_1203);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_12 <=
      ~_GEN_1375 & (_GEN_12 ? ~_GEN_1312 & _GEN_1204 : ~_GEN_1249 & _GEN_1204);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_13 <=
      ~_GEN_1377 & (_GEN_12 ? ~_GEN_1314 & _GEN_1205 : ~_GEN_1251 & _GEN_1205);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_14 <=
      ~_GEN_1379 & (_GEN_12 ? ~_GEN_1316 & _GEN_1206 : ~_GEN_1253 & _GEN_1206);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_15 <=
      ~_GEN_1381 & (_GEN_12 ? ~_GEN_1318 & _GEN_1207 : ~_GEN_1255 & _GEN_1207);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_16 <=
      ~_GEN_1383 & (_GEN_12 ? ~_GEN_1320 & _GEN_1208 : ~_GEN_1257 & _GEN_1208);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_17 <=
      ~_GEN_1385 & (_GEN_12 ? ~_GEN_1322 & _GEN_1209 : ~_GEN_1259 & _GEN_1209);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_18 <=
      ~_GEN_1387 & (_GEN_12 ? ~_GEN_1324 & _GEN_1210 : ~_GEN_1261 & _GEN_1210);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_19 <=
      ~_GEN_1389 & (_GEN_12 ? ~_GEN_1326 & _GEN_1211 : ~_GEN_1263 & _GEN_1211);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_20 <=
      ~_GEN_1391 & (_GEN_12 ? ~_GEN_1328 & _GEN_1212 : ~_GEN_1265 & _GEN_1212);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_21 <=
      ~_GEN_1393 & (_GEN_12 ? ~_GEN_1330 & _GEN_1213 : ~_GEN_1267 & _GEN_1213);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_22 <=
      ~_GEN_1395 & (_GEN_12 ? ~_GEN_1332 & _GEN_1214 : ~_GEN_1269 & _GEN_1214);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_23 <=
      ~_GEN_1397 & (_GEN_12 ? ~_GEN_1334 & _GEN_1215 : ~_GEN_1271 & _GEN_1215);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_24 <=
      ~_GEN_1399 & (_GEN_12 ? ~_GEN_1336 & _GEN_1216 : ~_GEN_1273 & _GEN_1216);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_25 <=
      ~_GEN_1401 & (_GEN_12 ? ~_GEN_1338 & _GEN_1217 : ~_GEN_1275 & _GEN_1217);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_26 <=
      ~_GEN_1403 & (_GEN_12 ? ~_GEN_1340 & _GEN_1218 : ~_GEN_1277 & _GEN_1218);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_27 <=
      ~_GEN_1405 & (_GEN_12 ? ~_GEN_1342 & _GEN_1219 : ~_GEN_1279 & _GEN_1219);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_28 <=
      ~_GEN_1407 & (_GEN_12 ? ~_GEN_1344 & _GEN_1220 : ~_GEN_1281 & _GEN_1220);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_29 <=
      ~_GEN_1409 & (_GEN_12 ? ~_GEN_1346 & _GEN_1221 : ~_GEN_1283 & _GEN_1221);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_30 <=
      ~_GEN_1411 & (_GEN_12 ? ~_GEN_1348 & _GEN_1222 : ~_GEN_1285 & _GEN_1222);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_31 <=
      ~_GEN_1412 & (_GEN_12 ? ~_GEN_1349 & _GEN_1223 : ~_GEN_1286 & _GEN_1223);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    if (_GEN_148) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_0_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_0_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_0_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_0_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_0_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_0_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_0_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_0_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_0_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_0_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_0_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_0_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_0_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_0_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_0_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_0_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1507) | ~rob_val_0) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_148)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_0_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_0_br_mask <= rob_uop_0_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_150) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_1_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_1_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_1_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_1_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_1_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_1_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_1_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_1_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_1_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_1_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_1_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_1_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_1_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1508) | ~rob_val_1) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_150)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_br_mask <= rob_uop_1_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_152) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_2_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_2_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_2_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_2_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_2_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_2_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_2_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_2_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_2_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_2_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_2_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_2_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_2_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1509) | ~rob_val_2) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_152)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_br_mask <= rob_uop_2_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_154) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_3_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_3_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_3_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_3_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_3_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_3_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_3_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_3_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_3_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_3_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_3_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_3_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_3_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1510) | ~rob_val_3) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_154)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_br_mask <= rob_uop_3_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_156) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_4_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_4_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_4_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_4_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_4_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_4_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_4_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_4_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_4_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_4_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_4_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_4_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_4_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_4_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_4_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_4_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1511) | ~rob_val_4) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_156)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_4_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_4_br_mask <= rob_uop_4_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_158) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_5_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_5_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_5_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_5_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_5_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_5_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_5_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_5_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_5_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_5_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_5_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_5_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_5_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_5_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_5_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_5_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1512) | ~rob_val_5) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_158)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_5_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_5_br_mask <= rob_uop_5_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_160) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_6_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_6_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_6_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_6_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_6_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_6_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_6_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_6_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_6_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_6_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_6_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_6_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_6_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_6_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_6_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_6_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1513) | ~rob_val_6) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_160)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_6_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_6_br_mask <= rob_uop_6_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_162) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_7_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_7_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_7_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_7_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_7_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_7_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_7_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_7_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_7_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_7_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_7_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_7_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_7_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_7_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_7_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_7_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1514) | ~rob_val_7) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_162)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_7_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_7_br_mask <= rob_uop_7_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_164) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_8_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_8_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_8_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_8_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_8_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_8_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_8_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_8_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_8_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_8_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_8_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_8_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_8_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_8_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_8_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_8_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1515) | ~rob_val_8) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_164)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_8_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_8_br_mask <= rob_uop_8_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_166) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_9_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_9_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_9_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_9_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_9_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_9_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_9_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_9_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_9_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_9_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_9_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_9_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_9_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_9_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_9_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_9_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1516) | ~rob_val_9) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_166)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_9_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_9_br_mask <= rob_uop_9_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_168) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_10_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_10_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_10_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_10_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_10_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_10_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_10_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_10_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_10_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_10_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_10_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_10_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_10_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_10_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_10_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_10_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1517) | ~rob_val_10) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_168)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_10_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_10_br_mask <= rob_uop_10_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_170) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_11_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_11_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_11_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_11_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_11_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_11_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_11_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_11_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_11_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_11_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_11_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_11_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_11_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_11_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_11_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_11_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1518) | ~rob_val_11) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_170)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_11_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_11_br_mask <= rob_uop_11_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_172) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_12_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_12_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_12_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_12_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_12_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_12_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_12_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_12_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_12_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_12_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_12_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_12_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_12_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_12_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_12_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_12_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1519) | ~rob_val_12) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_172)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_12_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_12_br_mask <= rob_uop_12_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_174) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_13_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_13_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_13_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_13_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_13_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_13_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_13_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_13_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_13_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_13_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_13_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_13_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_13_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_13_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_13_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_13_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1520) | ~rob_val_13) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_174)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_13_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_13_br_mask <= rob_uop_13_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_176) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_14_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_14_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_14_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_14_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_14_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_14_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_14_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_14_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_14_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_14_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_14_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_14_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_14_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_14_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_14_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_14_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1521) | ~rob_val_14) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_176)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_14_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_14_br_mask <= rob_uop_14_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_178) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_15_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_15_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_15_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_15_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_15_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_15_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_15_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_15_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_15_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_15_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_15_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_15_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_15_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_15_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_15_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_15_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1522) | ~rob_val_15) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_178)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_15_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_15_br_mask <= rob_uop_15_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_180) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_16_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_16_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_16_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_16_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_16_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_16_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_16_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_16_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_16_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_16_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_16_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_16_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_16_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_16_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_16_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_16_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1523) | ~rob_val_16) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_180)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_16_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_16_br_mask <= rob_uop_16_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_182) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_17_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_17_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_17_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_17_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_17_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_17_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_17_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_17_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_17_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_17_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_17_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_17_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_17_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_17_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_17_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_17_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1524) | ~rob_val_17) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_182)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_17_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_17_br_mask <= rob_uop_17_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_184) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_18_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_18_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_18_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_18_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_18_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_18_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_18_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_18_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_18_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_18_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_18_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_18_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_18_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_18_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_18_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_18_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1525) | ~rob_val_18) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_184)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_18_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_18_br_mask <= rob_uop_18_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_186) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_19_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_19_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_19_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_19_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_19_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_19_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_19_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_19_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_19_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_19_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_19_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_19_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_19_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_19_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_19_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_19_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1526) | ~rob_val_19) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_186)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_19_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_19_br_mask <= rob_uop_19_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_188) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_20_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_20_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_20_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_20_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_20_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_20_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_20_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_20_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_20_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_20_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_20_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_20_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_20_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_20_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_20_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_20_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1527) | ~rob_val_20) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_188)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_20_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_20_br_mask <= rob_uop_20_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_190) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_21_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_21_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_21_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_21_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_21_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_21_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_21_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_21_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_21_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_21_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_21_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_21_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_21_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_21_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_21_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_21_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1528) | ~rob_val_21) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_190)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_21_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_21_br_mask <= rob_uop_21_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_192) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_22_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_22_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_22_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_22_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_22_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_22_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_22_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_22_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_22_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_22_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_22_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_22_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_22_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_22_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_22_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_22_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1529) | ~rob_val_22) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_192)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_22_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_22_br_mask <= rob_uop_22_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_194) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_23_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_23_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_23_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_23_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_23_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_23_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_23_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_23_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_23_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_23_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_23_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_23_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_23_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_23_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_23_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_23_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1530) | ~rob_val_23) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_194)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_23_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_23_br_mask <= rob_uop_23_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_196) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_24_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_24_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_24_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_24_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_24_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_24_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_24_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_24_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_24_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_24_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_24_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_24_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_24_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_24_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_24_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_24_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1531) | ~rob_val_24) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_196)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_24_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_24_br_mask <= rob_uop_24_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_198) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_25_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_25_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_25_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_25_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_25_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_25_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_25_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_25_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_25_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_25_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_25_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_25_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_25_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_25_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_25_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_25_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1532) | ~rob_val_25) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_198)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_25_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_25_br_mask <= rob_uop_25_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_200) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_26_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_26_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_26_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_26_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_26_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_26_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_26_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_26_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_26_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_26_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_26_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_26_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_26_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_26_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_26_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_26_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1533) | ~rob_val_26) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_200)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_26_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_26_br_mask <= rob_uop_26_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_202) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_27_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_27_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_27_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_27_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_27_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_27_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_27_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_27_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_27_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_27_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_27_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_27_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_27_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_27_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_27_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_27_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1534) | ~rob_val_27) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_202)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_27_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_27_br_mask <= rob_uop_27_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_204) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_28_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_28_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_28_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_28_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_28_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_28_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_28_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_28_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_28_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_28_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_28_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_28_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_28_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_28_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_28_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_28_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1535) | ~rob_val_28) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_204)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_28_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_28_br_mask <= rob_uop_28_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_206) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_29_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_29_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_29_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_29_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_29_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_29_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_29_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_29_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_29_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_29_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_29_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_29_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_29_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_29_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_29_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_29_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1536) | ~rob_val_29) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_206)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_29_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_29_br_mask <= rob_uop_29_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_208) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_30_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_30_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_30_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_30_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_30_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_30_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_30_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_30_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_30_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_30_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_30_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_30_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_30_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_30_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_30_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_30_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1537) | ~rob_val_30) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_208)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_30_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_30_br_mask <= rob_uop_30_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_209) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_31_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_31_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_31_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_31_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_31_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_31_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_31_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_31_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_31_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_31_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_31_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_31_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_31_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_31_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_31_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_31_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1538) | ~rob_val_31) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_209)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_31_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_31_br_mask <= rob_uop_31_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    rob_exception_0 <=
      ~_GEN_1445
      & (_GEN_14 & _GEN_1413 | (_GEN_148 ? io_enq_uops_0_exception : rob_exception_0));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1 <=
      ~_GEN_1447
      & (_GEN_14 & _GEN_1414 | (_GEN_150 ? io_enq_uops_0_exception : rob_exception_1));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2 <=
      ~_GEN_1449
      & (_GEN_14 & _GEN_1415 | (_GEN_152 ? io_enq_uops_0_exception : rob_exception_2));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3 <=
      ~_GEN_1451
      & (_GEN_14 & _GEN_1416 | (_GEN_154 ? io_enq_uops_0_exception : rob_exception_3));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_4 <=
      ~_GEN_1453
      & (_GEN_14 & _GEN_1417 | (_GEN_156 ? io_enq_uops_0_exception : rob_exception_4));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_5 <=
      ~_GEN_1455
      & (_GEN_14 & _GEN_1418 | (_GEN_158 ? io_enq_uops_0_exception : rob_exception_5));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_6 <=
      ~_GEN_1457
      & (_GEN_14 & _GEN_1419 | (_GEN_160 ? io_enq_uops_0_exception : rob_exception_6));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_7 <=
      ~_GEN_1459
      & (_GEN_14 & _GEN_1420 | (_GEN_162 ? io_enq_uops_0_exception : rob_exception_7));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_8 <=
      ~_GEN_1461
      & (_GEN_14 & _GEN_1421 | (_GEN_164 ? io_enq_uops_0_exception : rob_exception_8));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_9 <=
      ~_GEN_1463
      & (_GEN_14 & _GEN_1422 | (_GEN_166 ? io_enq_uops_0_exception : rob_exception_9));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_10 <=
      ~_GEN_1465
      & (_GEN_14 & _GEN_1423 | (_GEN_168 ? io_enq_uops_0_exception : rob_exception_10));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_11 <=
      ~_GEN_1467
      & (_GEN_14 & _GEN_1424 | (_GEN_170 ? io_enq_uops_0_exception : rob_exception_11));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_12 <=
      ~_GEN_1469
      & (_GEN_14 & _GEN_1425 | (_GEN_172 ? io_enq_uops_0_exception : rob_exception_12));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_13 <=
      ~_GEN_1471
      & (_GEN_14 & _GEN_1426 | (_GEN_174 ? io_enq_uops_0_exception : rob_exception_13));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_14 <=
      ~_GEN_1473
      & (_GEN_14 & _GEN_1427 | (_GEN_176 ? io_enq_uops_0_exception : rob_exception_14));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_15 <=
      ~_GEN_1475
      & (_GEN_14 & _GEN_1428 | (_GEN_178 ? io_enq_uops_0_exception : rob_exception_15));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_16 <=
      ~_GEN_1477
      & (_GEN_14 & _GEN_1429 | (_GEN_180 ? io_enq_uops_0_exception : rob_exception_16));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_17 <=
      ~_GEN_1479
      & (_GEN_14 & _GEN_1430 | (_GEN_182 ? io_enq_uops_0_exception : rob_exception_17));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_18 <=
      ~_GEN_1481
      & (_GEN_14 & _GEN_1431 | (_GEN_184 ? io_enq_uops_0_exception : rob_exception_18));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_19 <=
      ~_GEN_1483
      & (_GEN_14 & _GEN_1432 | (_GEN_186 ? io_enq_uops_0_exception : rob_exception_19));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_20 <=
      ~_GEN_1485
      & (_GEN_14 & _GEN_1433 | (_GEN_188 ? io_enq_uops_0_exception : rob_exception_20));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_21 <=
      ~_GEN_1487
      & (_GEN_14 & _GEN_1434 | (_GEN_190 ? io_enq_uops_0_exception : rob_exception_21));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_22 <=
      ~_GEN_1489
      & (_GEN_14 & _GEN_1435 | (_GEN_192 ? io_enq_uops_0_exception : rob_exception_22));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_23 <=
      ~_GEN_1491
      & (_GEN_14 & _GEN_1436 | (_GEN_194 ? io_enq_uops_0_exception : rob_exception_23));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_24 <=
      ~_GEN_1493
      & (_GEN_14 & _GEN_1437 | (_GEN_196 ? io_enq_uops_0_exception : rob_exception_24));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_25 <=
      ~_GEN_1495
      & (_GEN_14 & _GEN_1438 | (_GEN_198 ? io_enq_uops_0_exception : rob_exception_25));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_26 <=
      ~_GEN_1497
      & (_GEN_14 & _GEN_1439 | (_GEN_200 ? io_enq_uops_0_exception : rob_exception_26));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_27 <=
      ~_GEN_1499
      & (_GEN_14 & _GEN_1440 | (_GEN_202 ? io_enq_uops_0_exception : rob_exception_27));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_28 <=
      ~_GEN_1501
      & (_GEN_14 & _GEN_1441 | (_GEN_204 ? io_enq_uops_0_exception : rob_exception_28));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_29 <=
      ~_GEN_1503
      & (_GEN_14 & _GEN_1442 | (_GEN_206 ? io_enq_uops_0_exception : rob_exception_29));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_30 <=
      ~_GEN_1505
      & (_GEN_14 & _GEN_1443 | (_GEN_208 ? io_enq_uops_0_exception : rob_exception_30));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_31 <=
      ~_GEN_1506
      & (_GEN_14 & (&(io_lxcpt_bits_uop_rob_idx[6:2]))
         | (_GEN_209 ? io_enq_uops_0_exception : rob_exception_31));	// rob.scala:236:31, :268:25, :307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_predicated_0 <=
      ~(_GEN_9 & _GEN_1097 | _GEN_1035 | _GEN_7 & _GEN_907)
      & (_GEN_845
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_717 | _GEN_655 | _GEN_3 & _GEN_527 | _GEN_465 | _GEN_1
               & _GEN_337)
             & (_GEN_275 ? io_wb_resps_0_bits_predicated : ~_GEN_148 & rob_predicated_0));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1 <=
      ~(_GEN_9 & _GEN_1100 | _GEN_1037 | _GEN_7 & _GEN_910)
      & (_GEN_847
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_720 | _GEN_657 | _GEN_3 & _GEN_530 | _GEN_467 | _GEN_1
               & _GEN_340)
             & (_GEN_277 ? io_wb_resps_0_bits_predicated : ~_GEN_150 & rob_predicated_1));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2 <=
      ~(_GEN_9 & _GEN_1103 | _GEN_1039 | _GEN_7 & _GEN_913)
      & (_GEN_849
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_723 | _GEN_659 | _GEN_3 & _GEN_533 | _GEN_469 | _GEN_1
               & _GEN_343)
             & (_GEN_279 ? io_wb_resps_0_bits_predicated : ~_GEN_152 & rob_predicated_2));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3 <=
      ~(_GEN_9 & _GEN_1106 | _GEN_1041 | _GEN_7 & _GEN_916)
      & (_GEN_851
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_726 | _GEN_661 | _GEN_3 & _GEN_536 | _GEN_471 | _GEN_1
               & _GEN_346)
             & (_GEN_281 ? io_wb_resps_0_bits_predicated : ~_GEN_154 & rob_predicated_3));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_4 <=
      ~(_GEN_9 & _GEN_1109 | _GEN_1043 | _GEN_7 & _GEN_919)
      & (_GEN_853
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_729 | _GEN_663 | _GEN_3 & _GEN_539 | _GEN_473 | _GEN_1
               & _GEN_349)
             & (_GEN_283 ? io_wb_resps_0_bits_predicated : ~_GEN_156 & rob_predicated_4));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_5 <=
      ~(_GEN_9 & _GEN_1112 | _GEN_1045 | _GEN_7 & _GEN_922)
      & (_GEN_855
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_732 | _GEN_665 | _GEN_3 & _GEN_542 | _GEN_475 | _GEN_1
               & _GEN_352)
             & (_GEN_285 ? io_wb_resps_0_bits_predicated : ~_GEN_158 & rob_predicated_5));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_6 <=
      ~(_GEN_9 & _GEN_1115 | _GEN_1047 | _GEN_7 & _GEN_925)
      & (_GEN_857
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_735 | _GEN_667 | _GEN_3 & _GEN_545 | _GEN_477 | _GEN_1
               & _GEN_355)
             & (_GEN_287 ? io_wb_resps_0_bits_predicated : ~_GEN_160 & rob_predicated_6));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_7 <=
      ~(_GEN_9 & _GEN_1118 | _GEN_1049 | _GEN_7 & _GEN_928)
      & (_GEN_859
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_738 | _GEN_669 | _GEN_3 & _GEN_548 | _GEN_479 | _GEN_1
               & _GEN_358)
             & (_GEN_289 ? io_wb_resps_0_bits_predicated : ~_GEN_162 & rob_predicated_7));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_8 <=
      ~(_GEN_9 & _GEN_1121 | _GEN_1051 | _GEN_7 & _GEN_931)
      & (_GEN_861
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_741 | _GEN_671 | _GEN_3 & _GEN_551 | _GEN_481 | _GEN_1
               & _GEN_361)
             & (_GEN_291 ? io_wb_resps_0_bits_predicated : ~_GEN_164 & rob_predicated_8));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_9 <=
      ~(_GEN_9 & _GEN_1124 | _GEN_1053 | _GEN_7 & _GEN_934)
      & (_GEN_863
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_744 | _GEN_673 | _GEN_3 & _GEN_554 | _GEN_483 | _GEN_1
               & _GEN_364)
             & (_GEN_293 ? io_wb_resps_0_bits_predicated : ~_GEN_166 & rob_predicated_9));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_10 <=
      ~(_GEN_9 & _GEN_1127 | _GEN_1055 | _GEN_7 & _GEN_937)
      & (_GEN_865
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_747 | _GEN_675 | _GEN_3 & _GEN_557 | _GEN_485 | _GEN_1
               & _GEN_367)
             & (_GEN_295
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_168 & rob_predicated_10));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_11 <=
      ~(_GEN_9 & _GEN_1130 | _GEN_1057 | _GEN_7 & _GEN_940)
      & (_GEN_867
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_750 | _GEN_677 | _GEN_3 & _GEN_560 | _GEN_487 | _GEN_1
               & _GEN_370)
             & (_GEN_297
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_170 & rob_predicated_11));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_12 <=
      ~(_GEN_9 & _GEN_1133 | _GEN_1059 | _GEN_7 & _GEN_943)
      & (_GEN_869
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_753 | _GEN_679 | _GEN_3 & _GEN_563 | _GEN_489 | _GEN_1
               & _GEN_373)
             & (_GEN_299
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_172 & rob_predicated_12));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_13 <=
      ~(_GEN_9 & _GEN_1136 | _GEN_1061 | _GEN_7 & _GEN_946)
      & (_GEN_871
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_756 | _GEN_681 | _GEN_3 & _GEN_566 | _GEN_491 | _GEN_1
               & _GEN_376)
             & (_GEN_301
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_174 & rob_predicated_13));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_14 <=
      ~(_GEN_9 & _GEN_1139 | _GEN_1063 | _GEN_7 & _GEN_949)
      & (_GEN_873
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_759 | _GEN_683 | _GEN_3 & _GEN_569 | _GEN_493 | _GEN_1
               & _GEN_379)
             & (_GEN_303
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_176 & rob_predicated_14));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_15 <=
      ~(_GEN_9 & _GEN_1142 | _GEN_1065 | _GEN_7 & _GEN_952)
      & (_GEN_875
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_762 | _GEN_685 | _GEN_3 & _GEN_572 | _GEN_495 | _GEN_1
               & _GEN_382)
             & (_GEN_305
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_178 & rob_predicated_15));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_16 <=
      ~(_GEN_9 & _GEN_1145 | _GEN_1067 | _GEN_7 & _GEN_955)
      & (_GEN_877
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_765 | _GEN_687 | _GEN_3 & _GEN_575 | _GEN_497 | _GEN_1
               & _GEN_385)
             & (_GEN_307
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_180 & rob_predicated_16));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_17 <=
      ~(_GEN_9 & _GEN_1148 | _GEN_1069 | _GEN_7 & _GEN_958)
      & (_GEN_879
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_768 | _GEN_689 | _GEN_3 & _GEN_578 | _GEN_499 | _GEN_1
               & _GEN_388)
             & (_GEN_309
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_182 & rob_predicated_17));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_18 <=
      ~(_GEN_9 & _GEN_1151 | _GEN_1071 | _GEN_7 & _GEN_961)
      & (_GEN_881
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_771 | _GEN_691 | _GEN_3 & _GEN_581 | _GEN_501 | _GEN_1
               & _GEN_391)
             & (_GEN_311
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_184 & rob_predicated_18));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_19 <=
      ~(_GEN_9 & _GEN_1154 | _GEN_1073 | _GEN_7 & _GEN_964)
      & (_GEN_883
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_774 | _GEN_693 | _GEN_3 & _GEN_584 | _GEN_503 | _GEN_1
               & _GEN_394)
             & (_GEN_313
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_186 & rob_predicated_19));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_20 <=
      ~(_GEN_9 & _GEN_1157 | _GEN_1075 | _GEN_7 & _GEN_967)
      & (_GEN_885
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_777 | _GEN_695 | _GEN_3 & _GEN_587 | _GEN_505 | _GEN_1
               & _GEN_397)
             & (_GEN_315
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_188 & rob_predicated_20));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_21 <=
      ~(_GEN_9 & _GEN_1160 | _GEN_1077 | _GEN_7 & _GEN_970)
      & (_GEN_887
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_780 | _GEN_697 | _GEN_3 & _GEN_590 | _GEN_507 | _GEN_1
               & _GEN_400)
             & (_GEN_317
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_190 & rob_predicated_21));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_22 <=
      ~(_GEN_9 & _GEN_1163 | _GEN_1079 | _GEN_7 & _GEN_973)
      & (_GEN_889
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_783 | _GEN_699 | _GEN_3 & _GEN_593 | _GEN_509 | _GEN_1
               & _GEN_403)
             & (_GEN_319
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_192 & rob_predicated_22));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_23 <=
      ~(_GEN_9 & _GEN_1166 | _GEN_1081 | _GEN_7 & _GEN_976)
      & (_GEN_891
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_786 | _GEN_701 | _GEN_3 & _GEN_596 | _GEN_511 | _GEN_1
               & _GEN_406)
             & (_GEN_321
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_194 & rob_predicated_23));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_24 <=
      ~(_GEN_9 & _GEN_1169 | _GEN_1083 | _GEN_7 & _GEN_979)
      & (_GEN_893
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_789 | _GEN_703 | _GEN_3 & _GEN_599 | _GEN_513 | _GEN_1
               & _GEN_409)
             & (_GEN_323
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_196 & rob_predicated_24));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_25 <=
      ~(_GEN_9 & _GEN_1172 | _GEN_1085 | _GEN_7 & _GEN_982)
      & (_GEN_895
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_792 | _GEN_705 | _GEN_3 & _GEN_602 | _GEN_515 | _GEN_1
               & _GEN_412)
             & (_GEN_325
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_198 & rob_predicated_25));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_26 <=
      ~(_GEN_9 & _GEN_1175 | _GEN_1087 | _GEN_7 & _GEN_985)
      & (_GEN_897
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_795 | _GEN_707 | _GEN_3 & _GEN_605 | _GEN_517 | _GEN_1
               & _GEN_415)
             & (_GEN_327
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_200 & rob_predicated_26));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_27 <=
      ~(_GEN_9 & _GEN_1178 | _GEN_1089 | _GEN_7 & _GEN_988)
      & (_GEN_899
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_798 | _GEN_709 | _GEN_3 & _GEN_608 | _GEN_519 | _GEN_1
               & _GEN_418)
             & (_GEN_329
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_202 & rob_predicated_27));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_28 <=
      ~(_GEN_9 & _GEN_1181 | _GEN_1091 | _GEN_7 & _GEN_991)
      & (_GEN_901
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_801 | _GEN_711 | _GEN_3 & _GEN_611 | _GEN_521 | _GEN_1
               & _GEN_421)
             & (_GEN_331
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_204 & rob_predicated_28));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_29 <=
      ~(_GEN_9 & _GEN_1184 | _GEN_1093 | _GEN_7 & _GEN_994)
      & (_GEN_903
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_804 | _GEN_713 | _GEN_3 & _GEN_614 | _GEN_523 | _GEN_1
               & _GEN_424)
             & (_GEN_333
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_206 & rob_predicated_29));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_30 <=
      ~(_GEN_9 & _GEN_1187 | _GEN_1095 | _GEN_7 & _GEN_997)
      & (_GEN_905
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & _GEN_807 | _GEN_715 | _GEN_3 & _GEN_617 | _GEN_525 | _GEN_1
               & _GEN_427)
             & (_GEN_335
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_208 & rob_predicated_30));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_31 <=
      ~(_GEN_9 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1096 | _GEN_7
        & (&(io_wb_resps_7_bits_uop_rob_idx[6:2])))
      & (_GEN_906
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_5 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_716 | _GEN_3
               & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_526 | _GEN_1
               & (&(io_wb_resps_1_bits_uop_rob_idx[6:2])))
             & (_GEN_336
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_209 & rob_predicated_31));	// rob.scala:236:31, :268:25, :307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_bsy_1_0 <=
      ~_GEN_2339 & (_GEN_47 ? ~_GEN_2307 & _GEN_2180 : ~_GEN_2275 & _GEN_2180);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_1 <=
      ~_GEN_2340 & (_GEN_47 ? ~_GEN_2308 & _GEN_2182 : ~_GEN_2276 & _GEN_2182);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_2 <=
      ~_GEN_2341 & (_GEN_47 ? ~_GEN_2309 & _GEN_2184 : ~_GEN_2277 & _GEN_2184);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_3 <=
      ~_GEN_2342 & (_GEN_47 ? ~_GEN_2310 & _GEN_2186 : ~_GEN_2278 & _GEN_2186);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_4 <=
      ~_GEN_2343 & (_GEN_47 ? ~_GEN_2311 & _GEN_2188 : ~_GEN_2279 & _GEN_2188);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_5 <=
      ~_GEN_2344 & (_GEN_47 ? ~_GEN_2312 & _GEN_2190 : ~_GEN_2280 & _GEN_2190);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_6 <=
      ~_GEN_2345 & (_GEN_47 ? ~_GEN_2313 & _GEN_2192 : ~_GEN_2281 & _GEN_2192);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_7 <=
      ~_GEN_2346 & (_GEN_47 ? ~_GEN_2314 & _GEN_2194 : ~_GEN_2282 & _GEN_2194);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_8 <=
      ~_GEN_2347 & (_GEN_47 ? ~_GEN_2315 & _GEN_2196 : ~_GEN_2283 & _GEN_2196);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_9 <=
      ~_GEN_2348 & (_GEN_47 ? ~_GEN_2316 & _GEN_2198 : ~_GEN_2284 & _GEN_2198);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_10 <=
      ~_GEN_2349 & (_GEN_47 ? ~_GEN_2317 & _GEN_2200 : ~_GEN_2285 & _GEN_2200);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_11 <=
      ~_GEN_2350 & (_GEN_47 ? ~_GEN_2318 & _GEN_2202 : ~_GEN_2286 & _GEN_2202);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_12 <=
      ~_GEN_2351 & (_GEN_47 ? ~_GEN_2319 & _GEN_2204 : ~_GEN_2287 & _GEN_2204);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_13 <=
      ~_GEN_2352 & (_GEN_47 ? ~_GEN_2320 & _GEN_2206 : ~_GEN_2288 & _GEN_2206);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_14 <=
      ~_GEN_2353 & (_GEN_47 ? ~_GEN_2321 & _GEN_2208 : ~_GEN_2289 & _GEN_2208);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_15 <=
      ~_GEN_2354 & (_GEN_47 ? ~_GEN_2322 & _GEN_2210 : ~_GEN_2290 & _GEN_2210);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_16 <=
      ~_GEN_2355 & (_GEN_47 ? ~_GEN_2323 & _GEN_2212 : ~_GEN_2291 & _GEN_2212);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_17 <=
      ~_GEN_2356 & (_GEN_47 ? ~_GEN_2324 & _GEN_2214 : ~_GEN_2292 & _GEN_2214);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_18 <=
      ~_GEN_2357 & (_GEN_47 ? ~_GEN_2325 & _GEN_2216 : ~_GEN_2293 & _GEN_2216);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_19 <=
      ~_GEN_2358 & (_GEN_47 ? ~_GEN_2326 & _GEN_2218 : ~_GEN_2294 & _GEN_2218);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_20 <=
      ~_GEN_2359 & (_GEN_47 ? ~_GEN_2327 & _GEN_2220 : ~_GEN_2295 & _GEN_2220);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_21 <=
      ~_GEN_2360 & (_GEN_47 ? ~_GEN_2328 & _GEN_2222 : ~_GEN_2296 & _GEN_2222);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_22 <=
      ~_GEN_2361 & (_GEN_47 ? ~_GEN_2329 & _GEN_2224 : ~_GEN_2297 & _GEN_2224);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_23 <=
      ~_GEN_2362 & (_GEN_47 ? ~_GEN_2330 & _GEN_2226 : ~_GEN_2298 & _GEN_2226);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_24 <=
      ~_GEN_2363 & (_GEN_47 ? ~_GEN_2331 & _GEN_2228 : ~_GEN_2299 & _GEN_2228);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_25 <=
      ~_GEN_2364 & (_GEN_47 ? ~_GEN_2332 & _GEN_2230 : ~_GEN_2300 & _GEN_2230);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_26 <=
      ~_GEN_2365 & (_GEN_47 ? ~_GEN_2333 & _GEN_2232 : ~_GEN_2301 & _GEN_2232);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_27 <=
      ~_GEN_2366 & (_GEN_47 ? ~_GEN_2334 & _GEN_2234 : ~_GEN_2302 & _GEN_2234);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_28 <=
      ~_GEN_2367 & (_GEN_47 ? ~_GEN_2335 & _GEN_2236 : ~_GEN_2303 & _GEN_2236);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_29 <=
      ~_GEN_2368 & (_GEN_47 ? ~_GEN_2336 & _GEN_2238 : ~_GEN_2304 & _GEN_2238);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_30 <=
      ~_GEN_2369 & (_GEN_47 ? ~_GEN_2337 & _GEN_2240 : ~_GEN_2305 & _GEN_2240);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_1_31 <=
      ~_GEN_2370 & (_GEN_47 ? ~_GEN_2338 & _GEN_2242 : ~_GEN_2306 & _GEN_2242);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_unsafe_1_0 <=
      ~_GEN_2339 & (_GEN_47 ? ~_GEN_2307 & _GEN_2243 : ~_GEN_2275 & _GEN_2243);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_1 <=
      ~_GEN_2340 & (_GEN_47 ? ~_GEN_2308 & _GEN_2244 : ~_GEN_2276 & _GEN_2244);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_2 <=
      ~_GEN_2341 & (_GEN_47 ? ~_GEN_2309 & _GEN_2245 : ~_GEN_2277 & _GEN_2245);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_3 <=
      ~_GEN_2342 & (_GEN_47 ? ~_GEN_2310 & _GEN_2246 : ~_GEN_2278 & _GEN_2246);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_4 <=
      ~_GEN_2343 & (_GEN_47 ? ~_GEN_2311 & _GEN_2247 : ~_GEN_2279 & _GEN_2247);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_5 <=
      ~_GEN_2344 & (_GEN_47 ? ~_GEN_2312 & _GEN_2248 : ~_GEN_2280 & _GEN_2248);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_6 <=
      ~_GEN_2345 & (_GEN_47 ? ~_GEN_2313 & _GEN_2249 : ~_GEN_2281 & _GEN_2249);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_7 <=
      ~_GEN_2346 & (_GEN_47 ? ~_GEN_2314 & _GEN_2250 : ~_GEN_2282 & _GEN_2250);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_8 <=
      ~_GEN_2347 & (_GEN_47 ? ~_GEN_2315 & _GEN_2251 : ~_GEN_2283 & _GEN_2251);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_9 <=
      ~_GEN_2348 & (_GEN_47 ? ~_GEN_2316 & _GEN_2252 : ~_GEN_2284 & _GEN_2252);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_10 <=
      ~_GEN_2349 & (_GEN_47 ? ~_GEN_2317 & _GEN_2253 : ~_GEN_2285 & _GEN_2253);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_11 <=
      ~_GEN_2350 & (_GEN_47 ? ~_GEN_2318 & _GEN_2254 : ~_GEN_2286 & _GEN_2254);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_12 <=
      ~_GEN_2351 & (_GEN_47 ? ~_GEN_2319 & _GEN_2255 : ~_GEN_2287 & _GEN_2255);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_13 <=
      ~_GEN_2352 & (_GEN_47 ? ~_GEN_2320 & _GEN_2256 : ~_GEN_2288 & _GEN_2256);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_14 <=
      ~_GEN_2353 & (_GEN_47 ? ~_GEN_2321 & _GEN_2257 : ~_GEN_2289 & _GEN_2257);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_15 <=
      ~_GEN_2354 & (_GEN_47 ? ~_GEN_2322 & _GEN_2258 : ~_GEN_2290 & _GEN_2258);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_16 <=
      ~_GEN_2355 & (_GEN_47 ? ~_GEN_2323 & _GEN_2259 : ~_GEN_2291 & _GEN_2259);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_17 <=
      ~_GEN_2356 & (_GEN_47 ? ~_GEN_2324 & _GEN_2260 : ~_GEN_2292 & _GEN_2260);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_18 <=
      ~_GEN_2357 & (_GEN_47 ? ~_GEN_2325 & _GEN_2261 : ~_GEN_2293 & _GEN_2261);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_19 <=
      ~_GEN_2358 & (_GEN_47 ? ~_GEN_2326 & _GEN_2262 : ~_GEN_2294 & _GEN_2262);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_20 <=
      ~_GEN_2359 & (_GEN_47 ? ~_GEN_2327 & _GEN_2263 : ~_GEN_2295 & _GEN_2263);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_21 <=
      ~_GEN_2360 & (_GEN_47 ? ~_GEN_2328 & _GEN_2264 : ~_GEN_2296 & _GEN_2264);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_22 <=
      ~_GEN_2361 & (_GEN_47 ? ~_GEN_2329 & _GEN_2265 : ~_GEN_2297 & _GEN_2265);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_23 <=
      ~_GEN_2362 & (_GEN_47 ? ~_GEN_2330 & _GEN_2266 : ~_GEN_2298 & _GEN_2266);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_24 <=
      ~_GEN_2363 & (_GEN_47 ? ~_GEN_2331 & _GEN_2267 : ~_GEN_2299 & _GEN_2267);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_25 <=
      ~_GEN_2364 & (_GEN_47 ? ~_GEN_2332 & _GEN_2268 : ~_GEN_2300 & _GEN_2268);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_26 <=
      ~_GEN_2365 & (_GEN_47 ? ~_GEN_2333 & _GEN_2269 : ~_GEN_2301 & _GEN_2269);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_27 <=
      ~_GEN_2366 & (_GEN_47 ? ~_GEN_2334 & _GEN_2270 : ~_GEN_2302 & _GEN_2270);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_28 <=
      ~_GEN_2367 & (_GEN_47 ? ~_GEN_2335 & _GEN_2271 : ~_GEN_2303 & _GEN_2271);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_29 <=
      ~_GEN_2368 & (_GEN_47 ? ~_GEN_2336 & _GEN_2272 : ~_GEN_2304 & _GEN_2272);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_30 <=
      ~_GEN_2369 & (_GEN_47 ? ~_GEN_2337 & _GEN_2273 : ~_GEN_2305 & _GEN_2273);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_1_31 <=
      ~_GEN_2370 & (_GEN_47 ? ~_GEN_2338 & _GEN_2274 : ~_GEN_2306 & _GEN_2274);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    if (_GEN_1539) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_0_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_0_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_0_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_0_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_0_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_0_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_0_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_0_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_0_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_0_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_0_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_0_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_0_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_0_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_0_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_0_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2403) | ~rob_val_1_0) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1539)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_0_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_0_br_mask <= rob_uop_1_0_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1540) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_1_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_1_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_1_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_1_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_1_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_1_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_1_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_1_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_1_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_1_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_1_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_1_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_1_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_1_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_1_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_1_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2404) | ~rob_val_1_1) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1540)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_1_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_1_br_mask <= rob_uop_1_1_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1541) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_2_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_2_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_2_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_2_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_2_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_2_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_2_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_2_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_2_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_2_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_2_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_2_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_2_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_2_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_2_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_2_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2405) | ~rob_val_1_2) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1541)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_2_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_2_br_mask <= rob_uop_1_2_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1542) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_3_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_3_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_3_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_3_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_3_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_3_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_3_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_3_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_3_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_3_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_3_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_3_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_3_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_3_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_3_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_3_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2406) | ~rob_val_1_3) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1542)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_3_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_3_br_mask <= rob_uop_1_3_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1543) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_4_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_4_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_4_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_4_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_4_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_4_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_4_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_4_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_4_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_4_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_4_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_4_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_4_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_4_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_4_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_4_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2407) | ~rob_val_1_4) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1543)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_4_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_4_br_mask <= rob_uop_1_4_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1544) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_5_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_5_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_5_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_5_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_5_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_5_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_5_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_5_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_5_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_5_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_5_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_5_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_5_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_5_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_5_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_5_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2408) | ~rob_val_1_5) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1544)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_5_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_5_br_mask <= rob_uop_1_5_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1545) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_6_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_6_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_6_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_6_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_6_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_6_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_6_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_6_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_6_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_6_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_6_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_6_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_6_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_6_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_6_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_6_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2409) | ~rob_val_1_6) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1545)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_6_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_6_br_mask <= rob_uop_1_6_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1546) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_7_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_7_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_7_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_7_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_7_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_7_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_7_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_7_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_7_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_7_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_7_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_7_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_7_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_7_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_7_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_7_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2410) | ~rob_val_1_7) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1546)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_7_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_7_br_mask <= rob_uop_1_7_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1547) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_8_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_8_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_8_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_8_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_8_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_8_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_8_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_8_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_8_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_8_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_8_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_8_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_8_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_8_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_8_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_8_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2411) | ~rob_val_1_8) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1547)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_8_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_8_br_mask <= rob_uop_1_8_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1548) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_9_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_9_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_9_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_9_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_9_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_9_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_9_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_9_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_9_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_9_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_9_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_9_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_9_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_9_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_9_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_9_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2412) | ~rob_val_1_9) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1548)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_9_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_9_br_mask <= rob_uop_1_9_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1549) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_10_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_10_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_10_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_10_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_10_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_10_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_10_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_10_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_10_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_10_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_10_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_10_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_10_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_10_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_10_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_10_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2413) | ~rob_val_1_10) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1549)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_10_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_10_br_mask <= rob_uop_1_10_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1550) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_11_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_11_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_11_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_11_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_11_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_11_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_11_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_11_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_11_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_11_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_11_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_11_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_11_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_11_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_11_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_11_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2414) | ~rob_val_1_11) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1550)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_11_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_11_br_mask <= rob_uop_1_11_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1551) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_12_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_12_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_12_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_12_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_12_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_12_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_12_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_12_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_12_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_12_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_12_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_12_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_12_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_12_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_12_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_12_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2415) | ~rob_val_1_12) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1551)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_12_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_12_br_mask <= rob_uop_1_12_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1552) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_13_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_13_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_13_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_13_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_13_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_13_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_13_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_13_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_13_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_13_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_13_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_13_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_13_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_13_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_13_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_13_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2416) | ~rob_val_1_13) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1552)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_13_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_13_br_mask <= rob_uop_1_13_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1553) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_14_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_14_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_14_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_14_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_14_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_14_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_14_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_14_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_14_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_14_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_14_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_14_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_14_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_14_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_14_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_14_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2417) | ~rob_val_1_14) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1553)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_14_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_14_br_mask <= rob_uop_1_14_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1554) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_15_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_15_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_15_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_15_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_15_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_15_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_15_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_15_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_15_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_15_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_15_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_15_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_15_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_15_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_15_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_15_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2418) | ~rob_val_1_15) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1554)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_15_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_15_br_mask <= rob_uop_1_15_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1555) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_16_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_16_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_16_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_16_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_16_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_16_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_16_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_16_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_16_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_16_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_16_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_16_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_16_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_16_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_16_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_16_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2419) | ~rob_val_1_16) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1555)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_16_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_16_br_mask <= rob_uop_1_16_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1556) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_17_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_17_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_17_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_17_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_17_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_17_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_17_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_17_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_17_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_17_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_17_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_17_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_17_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_17_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_17_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_17_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2420) | ~rob_val_1_17) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1556)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_17_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_17_br_mask <= rob_uop_1_17_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1557) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_18_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_18_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_18_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_18_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_18_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_18_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_18_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_18_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_18_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_18_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_18_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_18_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_18_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_18_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_18_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_18_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2421) | ~rob_val_1_18) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1557)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_18_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_18_br_mask <= rob_uop_1_18_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1558) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_19_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_19_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_19_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_19_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_19_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_19_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_19_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_19_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_19_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_19_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_19_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_19_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_19_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_19_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_19_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_19_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2422) | ~rob_val_1_19) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1558)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_19_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_19_br_mask <= rob_uop_1_19_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1559) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_20_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_20_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_20_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_20_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_20_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_20_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_20_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_20_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_20_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_20_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_20_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_20_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_20_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_20_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_20_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_20_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2423) | ~rob_val_1_20) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1559)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_20_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_20_br_mask <= rob_uop_1_20_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1560) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_21_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_21_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_21_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_21_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_21_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_21_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_21_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_21_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_21_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_21_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_21_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_21_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_21_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_21_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_21_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_21_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2424) | ~rob_val_1_21) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1560)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_21_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_21_br_mask <= rob_uop_1_21_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1561) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_22_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_22_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_22_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_22_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_22_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_22_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_22_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_22_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_22_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_22_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_22_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_22_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_22_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_22_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_22_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_22_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2425) | ~rob_val_1_22) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1561)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_22_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_22_br_mask <= rob_uop_1_22_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1562) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_23_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_23_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_23_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_23_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_23_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_23_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_23_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_23_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_23_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_23_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_23_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_23_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_23_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_23_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_23_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_23_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2426) | ~rob_val_1_23) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1562)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_23_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_23_br_mask <= rob_uop_1_23_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1563) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_24_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_24_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_24_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_24_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_24_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_24_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_24_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_24_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_24_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_24_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_24_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_24_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_24_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_24_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_24_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_24_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2427) | ~rob_val_1_24) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1563)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_24_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_24_br_mask <= rob_uop_1_24_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1564) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_25_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_25_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_25_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_25_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_25_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_25_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_25_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_25_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_25_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_25_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_25_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_25_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_25_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_25_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_25_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_25_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2428) | ~rob_val_1_25) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1564)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_25_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_25_br_mask <= rob_uop_1_25_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1565) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_26_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_26_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_26_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_26_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_26_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_26_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_26_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_26_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_26_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_26_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_26_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_26_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_26_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_26_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_26_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_26_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2429) | ~rob_val_1_26) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1565)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_26_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_26_br_mask <= rob_uop_1_26_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1566) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_27_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_27_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_27_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_27_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_27_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_27_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_27_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_27_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_27_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_27_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_27_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_27_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_27_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_27_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_27_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_27_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2430) | ~rob_val_1_27) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1566)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_27_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_27_br_mask <= rob_uop_1_27_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1567) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_28_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_28_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_28_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_28_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_28_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_28_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_28_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_28_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_28_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_28_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_28_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_28_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_28_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_28_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_28_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_28_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2431) | ~rob_val_1_28) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1567)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_28_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_28_br_mask <= rob_uop_1_28_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1568) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_29_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_29_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_29_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_29_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_29_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_29_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_29_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_29_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_29_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_29_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_29_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_29_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_29_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_29_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_29_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_29_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2432) | ~rob_val_1_29) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1568)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_29_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_29_br_mask <= rob_uop_1_29_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1569) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_30_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_30_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_30_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_30_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_30_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_30_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_30_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_30_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_30_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_30_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_30_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_30_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_30_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_30_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_30_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_30_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2433) | ~rob_val_1_30) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1569)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_30_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_30_br_mask <= rob_uop_1_30_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1570) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_31_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_31_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_31_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_31_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_31_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_31_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_31_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_31_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_31_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_31_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_31_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_31_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_31_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_31_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_31_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_31_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2434) | ~rob_val_1_31) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1570)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_31_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_31_br_mask <= rob_uop_1_31_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    rob_exception_1_0 <=
      ~_GEN_2371
      & (_GEN_49 & _GEN_1413 | (_GEN_1539 ? io_enq_uops_1_exception : rob_exception_1_0));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_1 <=
      ~_GEN_2372
      & (_GEN_49 & _GEN_1414 | (_GEN_1540 ? io_enq_uops_1_exception : rob_exception_1_1));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_2 <=
      ~_GEN_2373
      & (_GEN_49 & _GEN_1415 | (_GEN_1541 ? io_enq_uops_1_exception : rob_exception_1_2));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_3 <=
      ~_GEN_2374
      & (_GEN_49 & _GEN_1416 | (_GEN_1542 ? io_enq_uops_1_exception : rob_exception_1_3));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_4 <=
      ~_GEN_2375
      & (_GEN_49 & _GEN_1417 | (_GEN_1543 ? io_enq_uops_1_exception : rob_exception_1_4));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_5 <=
      ~_GEN_2376
      & (_GEN_49 & _GEN_1418 | (_GEN_1544 ? io_enq_uops_1_exception : rob_exception_1_5));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_6 <=
      ~_GEN_2377
      & (_GEN_49 & _GEN_1419 | (_GEN_1545 ? io_enq_uops_1_exception : rob_exception_1_6));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_7 <=
      ~_GEN_2378
      & (_GEN_49 & _GEN_1420 | (_GEN_1546 ? io_enq_uops_1_exception : rob_exception_1_7));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_8 <=
      ~_GEN_2379
      & (_GEN_49 & _GEN_1421 | (_GEN_1547 ? io_enq_uops_1_exception : rob_exception_1_8));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_9 <=
      ~_GEN_2380
      & (_GEN_49 & _GEN_1422 | (_GEN_1548 ? io_enq_uops_1_exception : rob_exception_1_9));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_10 <=
      ~_GEN_2381
      & (_GEN_49 & _GEN_1423
         | (_GEN_1549 ? io_enq_uops_1_exception : rob_exception_1_10));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_11 <=
      ~_GEN_2382
      & (_GEN_49 & _GEN_1424
         | (_GEN_1550 ? io_enq_uops_1_exception : rob_exception_1_11));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_12 <=
      ~_GEN_2383
      & (_GEN_49 & _GEN_1425
         | (_GEN_1551 ? io_enq_uops_1_exception : rob_exception_1_12));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_13 <=
      ~_GEN_2384
      & (_GEN_49 & _GEN_1426
         | (_GEN_1552 ? io_enq_uops_1_exception : rob_exception_1_13));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_14 <=
      ~_GEN_2385
      & (_GEN_49 & _GEN_1427
         | (_GEN_1553 ? io_enq_uops_1_exception : rob_exception_1_14));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_15 <=
      ~_GEN_2386
      & (_GEN_49 & _GEN_1428
         | (_GEN_1554 ? io_enq_uops_1_exception : rob_exception_1_15));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_16 <=
      ~_GEN_2387
      & (_GEN_49 & _GEN_1429
         | (_GEN_1555 ? io_enq_uops_1_exception : rob_exception_1_16));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_17 <=
      ~_GEN_2388
      & (_GEN_49 & _GEN_1430
         | (_GEN_1556 ? io_enq_uops_1_exception : rob_exception_1_17));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_18 <=
      ~_GEN_2389
      & (_GEN_49 & _GEN_1431
         | (_GEN_1557 ? io_enq_uops_1_exception : rob_exception_1_18));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_19 <=
      ~_GEN_2390
      & (_GEN_49 & _GEN_1432
         | (_GEN_1558 ? io_enq_uops_1_exception : rob_exception_1_19));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_20 <=
      ~_GEN_2391
      & (_GEN_49 & _GEN_1433
         | (_GEN_1559 ? io_enq_uops_1_exception : rob_exception_1_20));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_21 <=
      ~_GEN_2392
      & (_GEN_49 & _GEN_1434
         | (_GEN_1560 ? io_enq_uops_1_exception : rob_exception_1_21));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_22 <=
      ~_GEN_2393
      & (_GEN_49 & _GEN_1435
         | (_GEN_1561 ? io_enq_uops_1_exception : rob_exception_1_22));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_23 <=
      ~_GEN_2394
      & (_GEN_49 & _GEN_1436
         | (_GEN_1562 ? io_enq_uops_1_exception : rob_exception_1_23));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_24 <=
      ~_GEN_2395
      & (_GEN_49 & _GEN_1437
         | (_GEN_1563 ? io_enq_uops_1_exception : rob_exception_1_24));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_25 <=
      ~_GEN_2396
      & (_GEN_49 & _GEN_1438
         | (_GEN_1564 ? io_enq_uops_1_exception : rob_exception_1_25));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_26 <=
      ~_GEN_2397
      & (_GEN_49 & _GEN_1439
         | (_GEN_1565 ? io_enq_uops_1_exception : rob_exception_1_26));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_27 <=
      ~_GEN_2398
      & (_GEN_49 & _GEN_1440
         | (_GEN_1566 ? io_enq_uops_1_exception : rob_exception_1_27));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_28 <=
      ~_GEN_2399
      & (_GEN_49 & _GEN_1441
         | (_GEN_1567 ? io_enq_uops_1_exception : rob_exception_1_28));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_29 <=
      ~_GEN_2400
      & (_GEN_49 & _GEN_1442
         | (_GEN_1568 ? io_enq_uops_1_exception : rob_exception_1_29));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_30 <=
      ~_GEN_2401
      & (_GEN_49 & _GEN_1443
         | (_GEN_1569 ? io_enq_uops_1_exception : rob_exception_1_30));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_31 <=
      ~_GEN_2402
      & (_GEN_49 & (&(io_lxcpt_bits_uop_rob_idx[6:2]))
         | (_GEN_1570 ? io_enq_uops_1_exception : rob_exception_1_31));	// rob.scala:236:31, :268:25, :307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_predicated_1_0 <=
      ~(_GEN_44 & _GEN_1097 | _GEN_2147 | _GEN_42 & _GEN_907)
      & (_GEN_2019
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_717 | _GEN_1891 | _GEN_38 & _GEN_527 | _GEN_1763 | _GEN_36
               & _GEN_337)
             & (_GEN_1635
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1539 & rob_predicated_1_0));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_1 <=
      ~(_GEN_44 & _GEN_1100 | _GEN_2148 | _GEN_42 & _GEN_910)
      & (_GEN_2020
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_720 | _GEN_1892 | _GEN_38 & _GEN_530 | _GEN_1764 | _GEN_36
               & _GEN_340)
             & (_GEN_1636
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1540 & rob_predicated_1_1));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_2 <=
      ~(_GEN_44 & _GEN_1103 | _GEN_2149 | _GEN_42 & _GEN_913)
      & (_GEN_2021
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_723 | _GEN_1893 | _GEN_38 & _GEN_533 | _GEN_1765 | _GEN_36
               & _GEN_343)
             & (_GEN_1637
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1541 & rob_predicated_1_2));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_3 <=
      ~(_GEN_44 & _GEN_1106 | _GEN_2150 | _GEN_42 & _GEN_916)
      & (_GEN_2022
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_726 | _GEN_1894 | _GEN_38 & _GEN_536 | _GEN_1766 | _GEN_36
               & _GEN_346)
             & (_GEN_1638
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1542 & rob_predicated_1_3));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_4 <=
      ~(_GEN_44 & _GEN_1109 | _GEN_2151 | _GEN_42 & _GEN_919)
      & (_GEN_2023
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_729 | _GEN_1895 | _GEN_38 & _GEN_539 | _GEN_1767 | _GEN_36
               & _GEN_349)
             & (_GEN_1639
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1543 & rob_predicated_1_4));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_5 <=
      ~(_GEN_44 & _GEN_1112 | _GEN_2152 | _GEN_42 & _GEN_922)
      & (_GEN_2024
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_732 | _GEN_1896 | _GEN_38 & _GEN_542 | _GEN_1768 | _GEN_36
               & _GEN_352)
             & (_GEN_1640
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1544 & rob_predicated_1_5));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_6 <=
      ~(_GEN_44 & _GEN_1115 | _GEN_2153 | _GEN_42 & _GEN_925)
      & (_GEN_2025
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_735 | _GEN_1897 | _GEN_38 & _GEN_545 | _GEN_1769 | _GEN_36
               & _GEN_355)
             & (_GEN_1641
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1545 & rob_predicated_1_6));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_7 <=
      ~(_GEN_44 & _GEN_1118 | _GEN_2154 | _GEN_42 & _GEN_928)
      & (_GEN_2026
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_738 | _GEN_1898 | _GEN_38 & _GEN_548 | _GEN_1770 | _GEN_36
               & _GEN_358)
             & (_GEN_1642
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1546 & rob_predicated_1_7));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_8 <=
      ~(_GEN_44 & _GEN_1121 | _GEN_2155 | _GEN_42 & _GEN_931)
      & (_GEN_2027
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_741 | _GEN_1899 | _GEN_38 & _GEN_551 | _GEN_1771 | _GEN_36
               & _GEN_361)
             & (_GEN_1643
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1547 & rob_predicated_1_8));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_9 <=
      ~(_GEN_44 & _GEN_1124 | _GEN_2156 | _GEN_42 & _GEN_934)
      & (_GEN_2028
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_744 | _GEN_1900 | _GEN_38 & _GEN_554 | _GEN_1772 | _GEN_36
               & _GEN_364)
             & (_GEN_1644
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1548 & rob_predicated_1_9));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_10 <=
      ~(_GEN_44 & _GEN_1127 | _GEN_2157 | _GEN_42 & _GEN_937)
      & (_GEN_2029
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_747 | _GEN_1901 | _GEN_38 & _GEN_557 | _GEN_1773 | _GEN_36
               & _GEN_367)
             & (_GEN_1645
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1549 & rob_predicated_1_10));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_11 <=
      ~(_GEN_44 & _GEN_1130 | _GEN_2158 | _GEN_42 & _GEN_940)
      & (_GEN_2030
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_750 | _GEN_1902 | _GEN_38 & _GEN_560 | _GEN_1774 | _GEN_36
               & _GEN_370)
             & (_GEN_1646
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1550 & rob_predicated_1_11));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_12 <=
      ~(_GEN_44 & _GEN_1133 | _GEN_2159 | _GEN_42 & _GEN_943)
      & (_GEN_2031
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_753 | _GEN_1903 | _GEN_38 & _GEN_563 | _GEN_1775 | _GEN_36
               & _GEN_373)
             & (_GEN_1647
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1551 & rob_predicated_1_12));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_13 <=
      ~(_GEN_44 & _GEN_1136 | _GEN_2160 | _GEN_42 & _GEN_946)
      & (_GEN_2032
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_756 | _GEN_1904 | _GEN_38 & _GEN_566 | _GEN_1776 | _GEN_36
               & _GEN_376)
             & (_GEN_1648
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1552 & rob_predicated_1_13));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_14 <=
      ~(_GEN_44 & _GEN_1139 | _GEN_2161 | _GEN_42 & _GEN_949)
      & (_GEN_2033
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_759 | _GEN_1905 | _GEN_38 & _GEN_569 | _GEN_1777 | _GEN_36
               & _GEN_379)
             & (_GEN_1649
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1553 & rob_predicated_1_14));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_15 <=
      ~(_GEN_44 & _GEN_1142 | _GEN_2162 | _GEN_42 & _GEN_952)
      & (_GEN_2034
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_762 | _GEN_1906 | _GEN_38 & _GEN_572 | _GEN_1778 | _GEN_36
               & _GEN_382)
             & (_GEN_1650
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1554 & rob_predicated_1_15));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_16 <=
      ~(_GEN_44 & _GEN_1145 | _GEN_2163 | _GEN_42 & _GEN_955)
      & (_GEN_2035
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_765 | _GEN_1907 | _GEN_38 & _GEN_575 | _GEN_1779 | _GEN_36
               & _GEN_385)
             & (_GEN_1651
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1555 & rob_predicated_1_16));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_17 <=
      ~(_GEN_44 & _GEN_1148 | _GEN_2164 | _GEN_42 & _GEN_958)
      & (_GEN_2036
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_768 | _GEN_1908 | _GEN_38 & _GEN_578 | _GEN_1780 | _GEN_36
               & _GEN_388)
             & (_GEN_1652
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1556 & rob_predicated_1_17));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_18 <=
      ~(_GEN_44 & _GEN_1151 | _GEN_2165 | _GEN_42 & _GEN_961)
      & (_GEN_2037
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_771 | _GEN_1909 | _GEN_38 & _GEN_581 | _GEN_1781 | _GEN_36
               & _GEN_391)
             & (_GEN_1653
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1557 & rob_predicated_1_18));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_19 <=
      ~(_GEN_44 & _GEN_1154 | _GEN_2166 | _GEN_42 & _GEN_964)
      & (_GEN_2038
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_774 | _GEN_1910 | _GEN_38 & _GEN_584 | _GEN_1782 | _GEN_36
               & _GEN_394)
             & (_GEN_1654
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1558 & rob_predicated_1_19));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_20 <=
      ~(_GEN_44 & _GEN_1157 | _GEN_2167 | _GEN_42 & _GEN_967)
      & (_GEN_2039
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_777 | _GEN_1911 | _GEN_38 & _GEN_587 | _GEN_1783 | _GEN_36
               & _GEN_397)
             & (_GEN_1655
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1559 & rob_predicated_1_20));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_21 <=
      ~(_GEN_44 & _GEN_1160 | _GEN_2168 | _GEN_42 & _GEN_970)
      & (_GEN_2040
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_780 | _GEN_1912 | _GEN_38 & _GEN_590 | _GEN_1784 | _GEN_36
               & _GEN_400)
             & (_GEN_1656
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1560 & rob_predicated_1_21));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_22 <=
      ~(_GEN_44 & _GEN_1163 | _GEN_2169 | _GEN_42 & _GEN_973)
      & (_GEN_2041
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_783 | _GEN_1913 | _GEN_38 & _GEN_593 | _GEN_1785 | _GEN_36
               & _GEN_403)
             & (_GEN_1657
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1561 & rob_predicated_1_22));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_23 <=
      ~(_GEN_44 & _GEN_1166 | _GEN_2170 | _GEN_42 & _GEN_976)
      & (_GEN_2042
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_786 | _GEN_1914 | _GEN_38 & _GEN_596 | _GEN_1786 | _GEN_36
               & _GEN_406)
             & (_GEN_1658
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1562 & rob_predicated_1_23));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_24 <=
      ~(_GEN_44 & _GEN_1169 | _GEN_2171 | _GEN_42 & _GEN_979)
      & (_GEN_2043
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_789 | _GEN_1915 | _GEN_38 & _GEN_599 | _GEN_1787 | _GEN_36
               & _GEN_409)
             & (_GEN_1659
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1563 & rob_predicated_1_24));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_25 <=
      ~(_GEN_44 & _GEN_1172 | _GEN_2172 | _GEN_42 & _GEN_982)
      & (_GEN_2044
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_792 | _GEN_1916 | _GEN_38 & _GEN_602 | _GEN_1788 | _GEN_36
               & _GEN_412)
             & (_GEN_1660
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1564 & rob_predicated_1_25));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_26 <=
      ~(_GEN_44 & _GEN_1175 | _GEN_2173 | _GEN_42 & _GEN_985)
      & (_GEN_2045
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_795 | _GEN_1917 | _GEN_38 & _GEN_605 | _GEN_1789 | _GEN_36
               & _GEN_415)
             & (_GEN_1661
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1565 & rob_predicated_1_26));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_27 <=
      ~(_GEN_44 & _GEN_1178 | _GEN_2174 | _GEN_42 & _GEN_988)
      & (_GEN_2046
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_798 | _GEN_1918 | _GEN_38 & _GEN_608 | _GEN_1790 | _GEN_36
               & _GEN_418)
             & (_GEN_1662
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1566 & rob_predicated_1_27));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_28 <=
      ~(_GEN_44 & _GEN_1181 | _GEN_2175 | _GEN_42 & _GEN_991)
      & (_GEN_2047
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_801 | _GEN_1919 | _GEN_38 & _GEN_611 | _GEN_1791 | _GEN_36
               & _GEN_421)
             & (_GEN_1663
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1567 & rob_predicated_1_28));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_29 <=
      ~(_GEN_44 & _GEN_1184 | _GEN_2176 | _GEN_42 & _GEN_994)
      & (_GEN_2048
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_804 | _GEN_1920 | _GEN_38 & _GEN_614 | _GEN_1792 | _GEN_36
               & _GEN_424)
             & (_GEN_1664
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1568 & rob_predicated_1_29));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_30 <=
      ~(_GEN_44 & _GEN_1187 | _GEN_2177 | _GEN_42 & _GEN_997)
      & (_GEN_2049
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & _GEN_807 | _GEN_1921 | _GEN_38 & _GEN_617 | _GEN_1793 | _GEN_36
               & _GEN_427)
             & (_GEN_1665
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1569 & rob_predicated_1_30));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_31 <=
      ~(_GEN_44 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_2178 | _GEN_42
        & (&(io_wb_resps_7_bits_uop_rob_idx[6:2])))
      & (_GEN_2050
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_40 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1922 | _GEN_38
               & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1794 | _GEN_36
               & (&(io_wb_resps_1_bits_uop_rob_idx[6:2])))
             & (_GEN_1666
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1570 & rob_predicated_1_31));	// rob.scala:236:31, :268:25, :307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_bsy_2_0 <=
      ~_GEN_3235 & (_GEN_82 ? ~_GEN_3203 & _GEN_3076 : ~_GEN_3171 & _GEN_3076);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_1 <=
      ~_GEN_3236 & (_GEN_82 ? ~_GEN_3204 & _GEN_3078 : ~_GEN_3172 & _GEN_3078);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_2 <=
      ~_GEN_3237 & (_GEN_82 ? ~_GEN_3205 & _GEN_3080 : ~_GEN_3173 & _GEN_3080);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_3 <=
      ~_GEN_3238 & (_GEN_82 ? ~_GEN_3206 & _GEN_3082 : ~_GEN_3174 & _GEN_3082);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_4 <=
      ~_GEN_3239 & (_GEN_82 ? ~_GEN_3207 & _GEN_3084 : ~_GEN_3175 & _GEN_3084);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_5 <=
      ~_GEN_3240 & (_GEN_82 ? ~_GEN_3208 & _GEN_3086 : ~_GEN_3176 & _GEN_3086);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_6 <=
      ~_GEN_3241 & (_GEN_82 ? ~_GEN_3209 & _GEN_3088 : ~_GEN_3177 & _GEN_3088);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_7 <=
      ~_GEN_3242 & (_GEN_82 ? ~_GEN_3210 & _GEN_3090 : ~_GEN_3178 & _GEN_3090);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_8 <=
      ~_GEN_3243 & (_GEN_82 ? ~_GEN_3211 & _GEN_3092 : ~_GEN_3179 & _GEN_3092);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_9 <=
      ~_GEN_3244 & (_GEN_82 ? ~_GEN_3212 & _GEN_3094 : ~_GEN_3180 & _GEN_3094);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_10 <=
      ~_GEN_3245 & (_GEN_82 ? ~_GEN_3213 & _GEN_3096 : ~_GEN_3181 & _GEN_3096);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_11 <=
      ~_GEN_3246 & (_GEN_82 ? ~_GEN_3214 & _GEN_3098 : ~_GEN_3182 & _GEN_3098);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_12 <=
      ~_GEN_3247 & (_GEN_82 ? ~_GEN_3215 & _GEN_3100 : ~_GEN_3183 & _GEN_3100);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_13 <=
      ~_GEN_3248 & (_GEN_82 ? ~_GEN_3216 & _GEN_3102 : ~_GEN_3184 & _GEN_3102);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_14 <=
      ~_GEN_3249 & (_GEN_82 ? ~_GEN_3217 & _GEN_3104 : ~_GEN_3185 & _GEN_3104);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_15 <=
      ~_GEN_3250 & (_GEN_82 ? ~_GEN_3218 & _GEN_3106 : ~_GEN_3186 & _GEN_3106);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_16 <=
      ~_GEN_3251 & (_GEN_82 ? ~_GEN_3219 & _GEN_3108 : ~_GEN_3187 & _GEN_3108);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_17 <=
      ~_GEN_3252 & (_GEN_82 ? ~_GEN_3220 & _GEN_3110 : ~_GEN_3188 & _GEN_3110);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_18 <=
      ~_GEN_3253 & (_GEN_82 ? ~_GEN_3221 & _GEN_3112 : ~_GEN_3189 & _GEN_3112);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_19 <=
      ~_GEN_3254 & (_GEN_82 ? ~_GEN_3222 & _GEN_3114 : ~_GEN_3190 & _GEN_3114);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_20 <=
      ~_GEN_3255 & (_GEN_82 ? ~_GEN_3223 & _GEN_3116 : ~_GEN_3191 & _GEN_3116);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_21 <=
      ~_GEN_3256 & (_GEN_82 ? ~_GEN_3224 & _GEN_3118 : ~_GEN_3192 & _GEN_3118);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_22 <=
      ~_GEN_3257 & (_GEN_82 ? ~_GEN_3225 & _GEN_3120 : ~_GEN_3193 & _GEN_3120);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_23 <=
      ~_GEN_3258 & (_GEN_82 ? ~_GEN_3226 & _GEN_3122 : ~_GEN_3194 & _GEN_3122);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_24 <=
      ~_GEN_3259 & (_GEN_82 ? ~_GEN_3227 & _GEN_3124 : ~_GEN_3195 & _GEN_3124);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_25 <=
      ~_GEN_3260 & (_GEN_82 ? ~_GEN_3228 & _GEN_3126 : ~_GEN_3196 & _GEN_3126);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_26 <=
      ~_GEN_3261 & (_GEN_82 ? ~_GEN_3229 & _GEN_3128 : ~_GEN_3197 & _GEN_3128);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_27 <=
      ~_GEN_3262 & (_GEN_82 ? ~_GEN_3230 & _GEN_3130 : ~_GEN_3198 & _GEN_3130);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_28 <=
      ~_GEN_3263 & (_GEN_82 ? ~_GEN_3231 & _GEN_3132 : ~_GEN_3199 & _GEN_3132);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_29 <=
      ~_GEN_3264 & (_GEN_82 ? ~_GEN_3232 & _GEN_3134 : ~_GEN_3200 & _GEN_3134);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_30 <=
      ~_GEN_3265 & (_GEN_82 ? ~_GEN_3233 & _GEN_3136 : ~_GEN_3201 & _GEN_3136);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_2_31 <=
      ~_GEN_3266 & (_GEN_82 ? ~_GEN_3234 & _GEN_3138 : ~_GEN_3202 & _GEN_3138);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_unsafe_2_0 <=
      ~_GEN_3235 & (_GEN_82 ? ~_GEN_3203 & _GEN_3139 : ~_GEN_3171 & _GEN_3139);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_1 <=
      ~_GEN_3236 & (_GEN_82 ? ~_GEN_3204 & _GEN_3140 : ~_GEN_3172 & _GEN_3140);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_2 <=
      ~_GEN_3237 & (_GEN_82 ? ~_GEN_3205 & _GEN_3141 : ~_GEN_3173 & _GEN_3141);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_3 <=
      ~_GEN_3238 & (_GEN_82 ? ~_GEN_3206 & _GEN_3142 : ~_GEN_3174 & _GEN_3142);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_4 <=
      ~_GEN_3239 & (_GEN_82 ? ~_GEN_3207 & _GEN_3143 : ~_GEN_3175 & _GEN_3143);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_5 <=
      ~_GEN_3240 & (_GEN_82 ? ~_GEN_3208 & _GEN_3144 : ~_GEN_3176 & _GEN_3144);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_6 <=
      ~_GEN_3241 & (_GEN_82 ? ~_GEN_3209 & _GEN_3145 : ~_GEN_3177 & _GEN_3145);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_7 <=
      ~_GEN_3242 & (_GEN_82 ? ~_GEN_3210 & _GEN_3146 : ~_GEN_3178 & _GEN_3146);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_8 <=
      ~_GEN_3243 & (_GEN_82 ? ~_GEN_3211 & _GEN_3147 : ~_GEN_3179 & _GEN_3147);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_9 <=
      ~_GEN_3244 & (_GEN_82 ? ~_GEN_3212 & _GEN_3148 : ~_GEN_3180 & _GEN_3148);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_10 <=
      ~_GEN_3245 & (_GEN_82 ? ~_GEN_3213 & _GEN_3149 : ~_GEN_3181 & _GEN_3149);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_11 <=
      ~_GEN_3246 & (_GEN_82 ? ~_GEN_3214 & _GEN_3150 : ~_GEN_3182 & _GEN_3150);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_12 <=
      ~_GEN_3247 & (_GEN_82 ? ~_GEN_3215 & _GEN_3151 : ~_GEN_3183 & _GEN_3151);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_13 <=
      ~_GEN_3248 & (_GEN_82 ? ~_GEN_3216 & _GEN_3152 : ~_GEN_3184 & _GEN_3152);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_14 <=
      ~_GEN_3249 & (_GEN_82 ? ~_GEN_3217 & _GEN_3153 : ~_GEN_3185 & _GEN_3153);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_15 <=
      ~_GEN_3250 & (_GEN_82 ? ~_GEN_3218 & _GEN_3154 : ~_GEN_3186 & _GEN_3154);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_16 <=
      ~_GEN_3251 & (_GEN_82 ? ~_GEN_3219 & _GEN_3155 : ~_GEN_3187 & _GEN_3155);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_17 <=
      ~_GEN_3252 & (_GEN_82 ? ~_GEN_3220 & _GEN_3156 : ~_GEN_3188 & _GEN_3156);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_18 <=
      ~_GEN_3253 & (_GEN_82 ? ~_GEN_3221 & _GEN_3157 : ~_GEN_3189 & _GEN_3157);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_19 <=
      ~_GEN_3254 & (_GEN_82 ? ~_GEN_3222 & _GEN_3158 : ~_GEN_3190 & _GEN_3158);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_20 <=
      ~_GEN_3255 & (_GEN_82 ? ~_GEN_3223 & _GEN_3159 : ~_GEN_3191 & _GEN_3159);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_21 <=
      ~_GEN_3256 & (_GEN_82 ? ~_GEN_3224 & _GEN_3160 : ~_GEN_3192 & _GEN_3160);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_22 <=
      ~_GEN_3257 & (_GEN_82 ? ~_GEN_3225 & _GEN_3161 : ~_GEN_3193 & _GEN_3161);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_23 <=
      ~_GEN_3258 & (_GEN_82 ? ~_GEN_3226 & _GEN_3162 : ~_GEN_3194 & _GEN_3162);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_24 <=
      ~_GEN_3259 & (_GEN_82 ? ~_GEN_3227 & _GEN_3163 : ~_GEN_3195 & _GEN_3163);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_25 <=
      ~_GEN_3260 & (_GEN_82 ? ~_GEN_3228 & _GEN_3164 : ~_GEN_3196 & _GEN_3164);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_26 <=
      ~_GEN_3261 & (_GEN_82 ? ~_GEN_3229 & _GEN_3165 : ~_GEN_3197 & _GEN_3165);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_27 <=
      ~_GEN_3262 & (_GEN_82 ? ~_GEN_3230 & _GEN_3166 : ~_GEN_3198 & _GEN_3166);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_28 <=
      ~_GEN_3263 & (_GEN_82 ? ~_GEN_3231 & _GEN_3167 : ~_GEN_3199 & _GEN_3167);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_29 <=
      ~_GEN_3264 & (_GEN_82 ? ~_GEN_3232 & _GEN_3168 : ~_GEN_3200 & _GEN_3168);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_30 <=
      ~_GEN_3265 & (_GEN_82 ? ~_GEN_3233 & _GEN_3169 : ~_GEN_3201 & _GEN_3169);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_2_31 <=
      ~_GEN_3266 & (_GEN_82 ? ~_GEN_3234 & _GEN_3170 : ~_GEN_3202 & _GEN_3170);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    if (_GEN_2435) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_0_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_0_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_0_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_0_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_0_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_0_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_0_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_0_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_0_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_0_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_0_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_0_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_0_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_0_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_0_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_0_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3299) | ~rob_val_2_0) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2435)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_0_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_0_br_mask <= rob_uop_2_0_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2436) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_1_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_1_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_1_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_1_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_1_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_1_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_1_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_1_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_1_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_1_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_1_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_1_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_1_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_1_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_1_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_1_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3300) | ~rob_val_2_1) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2436)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_1_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_1_br_mask <= rob_uop_2_1_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2437) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_2_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_2_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_2_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_2_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_2_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_2_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_2_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_2_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_2_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_2_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_2_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_2_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_2_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_2_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_2_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_2_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3301) | ~rob_val_2_2) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2437)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_2_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_2_br_mask <= rob_uop_2_2_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2438) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_3_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_3_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_3_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_3_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_3_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_3_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_3_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_3_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_3_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_3_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_3_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_3_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_3_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_3_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_3_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_3_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3302) | ~rob_val_2_3) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2438)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_3_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_3_br_mask <= rob_uop_2_3_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2439) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_4_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_4_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_4_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_4_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_4_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_4_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_4_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_4_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_4_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_4_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_4_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_4_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_4_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_4_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_4_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_4_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3303) | ~rob_val_2_4) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2439)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_4_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_4_br_mask <= rob_uop_2_4_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2440) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_5_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_5_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_5_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_5_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_5_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_5_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_5_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_5_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_5_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_5_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_5_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_5_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_5_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_5_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_5_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_5_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3304) | ~rob_val_2_5) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2440)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_5_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_5_br_mask <= rob_uop_2_5_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2441) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_6_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_6_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_6_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_6_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_6_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_6_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_6_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_6_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_6_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_6_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_6_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_6_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_6_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_6_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_6_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_6_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3305) | ~rob_val_2_6) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2441)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_6_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_6_br_mask <= rob_uop_2_6_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2442) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_7_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_7_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_7_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_7_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_7_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_7_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_7_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_7_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_7_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_7_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_7_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_7_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_7_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_7_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_7_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_7_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3306) | ~rob_val_2_7) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2442)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_7_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_7_br_mask <= rob_uop_2_7_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2443) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_8_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_8_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_8_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_8_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_8_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_8_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_8_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_8_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_8_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_8_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_8_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_8_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_8_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_8_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_8_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_8_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3307) | ~rob_val_2_8) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2443)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_8_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_8_br_mask <= rob_uop_2_8_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2444) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_9_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_9_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_9_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_9_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_9_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_9_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_9_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_9_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_9_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_9_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_9_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_9_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_9_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_9_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_9_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_9_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3308) | ~rob_val_2_9) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2444)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_9_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_9_br_mask <= rob_uop_2_9_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2445) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_10_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_10_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_10_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_10_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_10_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_10_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_10_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_10_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_10_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_10_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_10_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_10_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_10_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_10_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_10_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_10_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3309) | ~rob_val_2_10) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2445)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_10_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_10_br_mask <= rob_uop_2_10_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2446) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_11_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_11_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_11_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_11_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_11_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_11_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_11_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_11_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_11_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_11_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_11_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_11_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_11_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_11_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_11_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_11_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3310) | ~rob_val_2_11) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2446)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_11_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_11_br_mask <= rob_uop_2_11_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2447) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_12_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_12_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_12_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_12_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_12_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_12_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_12_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_12_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_12_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_12_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_12_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_12_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_12_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_12_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_12_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_12_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3311) | ~rob_val_2_12) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2447)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_12_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_12_br_mask <= rob_uop_2_12_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2448) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_13_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_13_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_13_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_13_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_13_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_13_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_13_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_13_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_13_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_13_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_13_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_13_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_13_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_13_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_13_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_13_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3312) | ~rob_val_2_13) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2448)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_13_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_13_br_mask <= rob_uop_2_13_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2449) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_14_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_14_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_14_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_14_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_14_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_14_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_14_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_14_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_14_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_14_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_14_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_14_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_14_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_14_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_14_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_14_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3313) | ~rob_val_2_14) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2449)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_14_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_14_br_mask <= rob_uop_2_14_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2450) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_15_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_15_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_15_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_15_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_15_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_15_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_15_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_15_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_15_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_15_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_15_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_15_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_15_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_15_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_15_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_15_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3314) | ~rob_val_2_15) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2450)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_15_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_15_br_mask <= rob_uop_2_15_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2451) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_16_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_16_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_16_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_16_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_16_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_16_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_16_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_16_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_16_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_16_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_16_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_16_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_16_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_16_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_16_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_16_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3315) | ~rob_val_2_16) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2451)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_16_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_16_br_mask <= rob_uop_2_16_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2452) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_17_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_17_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_17_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_17_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_17_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_17_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_17_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_17_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_17_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_17_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_17_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_17_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_17_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_17_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_17_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_17_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3316) | ~rob_val_2_17) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2452)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_17_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_17_br_mask <= rob_uop_2_17_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2453) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_18_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_18_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_18_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_18_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_18_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_18_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_18_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_18_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_18_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_18_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_18_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_18_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_18_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_18_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_18_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_18_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3317) | ~rob_val_2_18) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2453)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_18_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_18_br_mask <= rob_uop_2_18_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2454) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_19_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_19_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_19_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_19_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_19_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_19_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_19_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_19_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_19_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_19_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_19_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_19_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_19_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_19_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_19_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_19_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3318) | ~rob_val_2_19) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2454)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_19_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_19_br_mask <= rob_uop_2_19_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2455) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_20_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_20_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_20_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_20_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_20_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_20_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_20_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_20_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_20_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_20_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_20_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_20_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_20_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_20_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_20_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_20_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3319) | ~rob_val_2_20) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2455)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_20_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_20_br_mask <= rob_uop_2_20_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2456) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_21_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_21_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_21_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_21_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_21_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_21_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_21_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_21_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_21_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_21_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_21_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_21_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_21_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_21_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_21_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_21_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3320) | ~rob_val_2_21) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2456)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_21_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_21_br_mask <= rob_uop_2_21_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2457) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_22_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_22_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_22_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_22_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_22_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_22_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_22_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_22_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_22_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_22_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_22_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_22_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_22_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_22_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_22_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_22_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3321) | ~rob_val_2_22) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2457)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_22_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_22_br_mask <= rob_uop_2_22_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2458) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_23_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_23_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_23_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_23_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_23_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_23_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_23_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_23_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_23_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_23_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_23_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_23_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_23_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_23_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_23_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_23_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3322) | ~rob_val_2_23) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2458)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_23_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_23_br_mask <= rob_uop_2_23_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2459) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_24_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_24_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_24_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_24_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_24_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_24_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_24_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_24_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_24_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_24_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_24_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_24_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_24_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_24_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_24_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_24_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3323) | ~rob_val_2_24) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2459)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_24_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_24_br_mask <= rob_uop_2_24_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2460) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_25_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_25_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_25_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_25_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_25_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_25_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_25_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_25_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_25_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_25_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_25_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_25_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_25_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_25_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_25_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_25_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3324) | ~rob_val_2_25) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2460)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_25_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_25_br_mask <= rob_uop_2_25_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2461) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_26_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_26_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_26_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_26_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_26_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_26_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_26_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_26_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_26_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_26_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_26_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_26_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_26_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_26_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_26_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_26_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3325) | ~rob_val_2_26) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2461)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_26_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_26_br_mask <= rob_uop_2_26_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2462) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_27_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_27_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_27_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_27_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_27_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_27_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_27_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_27_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_27_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_27_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_27_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_27_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_27_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_27_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_27_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_27_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3326) | ~rob_val_2_27) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2462)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_27_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_27_br_mask <= rob_uop_2_27_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2463) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_28_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_28_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_28_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_28_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_28_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_28_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_28_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_28_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_28_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_28_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_28_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_28_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_28_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_28_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_28_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_28_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3327) | ~rob_val_2_28) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2463)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_28_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_28_br_mask <= rob_uop_2_28_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2464) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_29_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_29_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_29_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_29_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_29_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_29_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_29_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_29_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_29_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_29_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_29_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_29_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_29_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_29_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_29_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_29_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3328) | ~rob_val_2_29) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2464)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_29_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_29_br_mask <= rob_uop_2_29_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2465) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_30_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_30_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_30_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_30_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_30_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_30_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_30_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_30_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_30_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_30_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_30_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_30_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_30_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_30_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_30_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_30_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3329) | ~rob_val_2_30) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2465)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_30_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_30_br_mask <= rob_uop_2_30_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_2466) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_31_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_31_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_31_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_31_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_31_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_31_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_31_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_31_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_31_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_31_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_31_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_31_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_31_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_31_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_31_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_31_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_3330) | ~rob_val_2_31) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_2466)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_31_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_31_br_mask <= rob_uop_2_31_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    rob_exception_2_0 <=
      ~_GEN_3267
      & (_GEN_84 & _GEN_1413 | (_GEN_2435 ? io_enq_uops_2_exception : rob_exception_2_0));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_1 <=
      ~_GEN_3268
      & (_GEN_84 & _GEN_1414 | (_GEN_2436 ? io_enq_uops_2_exception : rob_exception_2_1));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_2 <=
      ~_GEN_3269
      & (_GEN_84 & _GEN_1415 | (_GEN_2437 ? io_enq_uops_2_exception : rob_exception_2_2));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_3 <=
      ~_GEN_3270
      & (_GEN_84 & _GEN_1416 | (_GEN_2438 ? io_enq_uops_2_exception : rob_exception_2_3));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_4 <=
      ~_GEN_3271
      & (_GEN_84 & _GEN_1417 | (_GEN_2439 ? io_enq_uops_2_exception : rob_exception_2_4));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_5 <=
      ~_GEN_3272
      & (_GEN_84 & _GEN_1418 | (_GEN_2440 ? io_enq_uops_2_exception : rob_exception_2_5));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_6 <=
      ~_GEN_3273
      & (_GEN_84 & _GEN_1419 | (_GEN_2441 ? io_enq_uops_2_exception : rob_exception_2_6));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_7 <=
      ~_GEN_3274
      & (_GEN_84 & _GEN_1420 | (_GEN_2442 ? io_enq_uops_2_exception : rob_exception_2_7));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_8 <=
      ~_GEN_3275
      & (_GEN_84 & _GEN_1421 | (_GEN_2443 ? io_enq_uops_2_exception : rob_exception_2_8));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_9 <=
      ~_GEN_3276
      & (_GEN_84 & _GEN_1422 | (_GEN_2444 ? io_enq_uops_2_exception : rob_exception_2_9));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_10 <=
      ~_GEN_3277
      & (_GEN_84 & _GEN_1423
         | (_GEN_2445 ? io_enq_uops_2_exception : rob_exception_2_10));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_11 <=
      ~_GEN_3278
      & (_GEN_84 & _GEN_1424
         | (_GEN_2446 ? io_enq_uops_2_exception : rob_exception_2_11));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_12 <=
      ~_GEN_3279
      & (_GEN_84 & _GEN_1425
         | (_GEN_2447 ? io_enq_uops_2_exception : rob_exception_2_12));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_13 <=
      ~_GEN_3280
      & (_GEN_84 & _GEN_1426
         | (_GEN_2448 ? io_enq_uops_2_exception : rob_exception_2_13));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_14 <=
      ~_GEN_3281
      & (_GEN_84 & _GEN_1427
         | (_GEN_2449 ? io_enq_uops_2_exception : rob_exception_2_14));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_15 <=
      ~_GEN_3282
      & (_GEN_84 & _GEN_1428
         | (_GEN_2450 ? io_enq_uops_2_exception : rob_exception_2_15));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_16 <=
      ~_GEN_3283
      & (_GEN_84 & _GEN_1429
         | (_GEN_2451 ? io_enq_uops_2_exception : rob_exception_2_16));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_17 <=
      ~_GEN_3284
      & (_GEN_84 & _GEN_1430
         | (_GEN_2452 ? io_enq_uops_2_exception : rob_exception_2_17));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_18 <=
      ~_GEN_3285
      & (_GEN_84 & _GEN_1431
         | (_GEN_2453 ? io_enq_uops_2_exception : rob_exception_2_18));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_19 <=
      ~_GEN_3286
      & (_GEN_84 & _GEN_1432
         | (_GEN_2454 ? io_enq_uops_2_exception : rob_exception_2_19));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_20 <=
      ~_GEN_3287
      & (_GEN_84 & _GEN_1433
         | (_GEN_2455 ? io_enq_uops_2_exception : rob_exception_2_20));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_21 <=
      ~_GEN_3288
      & (_GEN_84 & _GEN_1434
         | (_GEN_2456 ? io_enq_uops_2_exception : rob_exception_2_21));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_22 <=
      ~_GEN_3289
      & (_GEN_84 & _GEN_1435
         | (_GEN_2457 ? io_enq_uops_2_exception : rob_exception_2_22));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_23 <=
      ~_GEN_3290
      & (_GEN_84 & _GEN_1436
         | (_GEN_2458 ? io_enq_uops_2_exception : rob_exception_2_23));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_24 <=
      ~_GEN_3291
      & (_GEN_84 & _GEN_1437
         | (_GEN_2459 ? io_enq_uops_2_exception : rob_exception_2_24));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_25 <=
      ~_GEN_3292
      & (_GEN_84 & _GEN_1438
         | (_GEN_2460 ? io_enq_uops_2_exception : rob_exception_2_25));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_26 <=
      ~_GEN_3293
      & (_GEN_84 & _GEN_1439
         | (_GEN_2461 ? io_enq_uops_2_exception : rob_exception_2_26));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_27 <=
      ~_GEN_3294
      & (_GEN_84 & _GEN_1440
         | (_GEN_2462 ? io_enq_uops_2_exception : rob_exception_2_27));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_28 <=
      ~_GEN_3295
      & (_GEN_84 & _GEN_1441
         | (_GEN_2463 ? io_enq_uops_2_exception : rob_exception_2_28));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_29 <=
      ~_GEN_3296
      & (_GEN_84 & _GEN_1442
         | (_GEN_2464 ? io_enq_uops_2_exception : rob_exception_2_29));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_30 <=
      ~_GEN_3297
      & (_GEN_84 & _GEN_1443
         | (_GEN_2465 ? io_enq_uops_2_exception : rob_exception_2_30));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_31 <=
      ~_GEN_3298
      & (_GEN_84 & (&(io_lxcpt_bits_uop_rob_idx[6:2]))
         | (_GEN_2466 ? io_enq_uops_2_exception : rob_exception_2_31));	// rob.scala:236:31, :268:25, :307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_predicated_2_0 <=
      ~(_GEN_79 & _GEN_1097 | _GEN_3043 | _GEN_77 & _GEN_907)
      & (_GEN_2915
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_717 | _GEN_2787 | _GEN_73 & _GEN_527 | _GEN_2659 | _GEN_71
               & _GEN_337)
             & (_GEN_2531
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2435 & rob_predicated_2_0));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_1 <=
      ~(_GEN_79 & _GEN_1100 | _GEN_3044 | _GEN_77 & _GEN_910)
      & (_GEN_2916
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_720 | _GEN_2788 | _GEN_73 & _GEN_530 | _GEN_2660 | _GEN_71
               & _GEN_340)
             & (_GEN_2532
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2436 & rob_predicated_2_1));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_2 <=
      ~(_GEN_79 & _GEN_1103 | _GEN_3045 | _GEN_77 & _GEN_913)
      & (_GEN_2917
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_723 | _GEN_2789 | _GEN_73 & _GEN_533 | _GEN_2661 | _GEN_71
               & _GEN_343)
             & (_GEN_2533
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2437 & rob_predicated_2_2));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_3 <=
      ~(_GEN_79 & _GEN_1106 | _GEN_3046 | _GEN_77 & _GEN_916)
      & (_GEN_2918
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_726 | _GEN_2790 | _GEN_73 & _GEN_536 | _GEN_2662 | _GEN_71
               & _GEN_346)
             & (_GEN_2534
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2438 & rob_predicated_2_3));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_4 <=
      ~(_GEN_79 & _GEN_1109 | _GEN_3047 | _GEN_77 & _GEN_919)
      & (_GEN_2919
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_729 | _GEN_2791 | _GEN_73 & _GEN_539 | _GEN_2663 | _GEN_71
               & _GEN_349)
             & (_GEN_2535
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2439 & rob_predicated_2_4));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_5 <=
      ~(_GEN_79 & _GEN_1112 | _GEN_3048 | _GEN_77 & _GEN_922)
      & (_GEN_2920
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_732 | _GEN_2792 | _GEN_73 & _GEN_542 | _GEN_2664 | _GEN_71
               & _GEN_352)
             & (_GEN_2536
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2440 & rob_predicated_2_5));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_6 <=
      ~(_GEN_79 & _GEN_1115 | _GEN_3049 | _GEN_77 & _GEN_925)
      & (_GEN_2921
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_735 | _GEN_2793 | _GEN_73 & _GEN_545 | _GEN_2665 | _GEN_71
               & _GEN_355)
             & (_GEN_2537
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2441 & rob_predicated_2_6));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_7 <=
      ~(_GEN_79 & _GEN_1118 | _GEN_3050 | _GEN_77 & _GEN_928)
      & (_GEN_2922
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_738 | _GEN_2794 | _GEN_73 & _GEN_548 | _GEN_2666 | _GEN_71
               & _GEN_358)
             & (_GEN_2538
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2442 & rob_predicated_2_7));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_8 <=
      ~(_GEN_79 & _GEN_1121 | _GEN_3051 | _GEN_77 & _GEN_931)
      & (_GEN_2923
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_741 | _GEN_2795 | _GEN_73 & _GEN_551 | _GEN_2667 | _GEN_71
               & _GEN_361)
             & (_GEN_2539
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2443 & rob_predicated_2_8));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_9 <=
      ~(_GEN_79 & _GEN_1124 | _GEN_3052 | _GEN_77 & _GEN_934)
      & (_GEN_2924
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_744 | _GEN_2796 | _GEN_73 & _GEN_554 | _GEN_2668 | _GEN_71
               & _GEN_364)
             & (_GEN_2540
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2444 & rob_predicated_2_9));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_10 <=
      ~(_GEN_79 & _GEN_1127 | _GEN_3053 | _GEN_77 & _GEN_937)
      & (_GEN_2925
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_747 | _GEN_2797 | _GEN_73 & _GEN_557 | _GEN_2669 | _GEN_71
               & _GEN_367)
             & (_GEN_2541
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2445 & rob_predicated_2_10));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_11 <=
      ~(_GEN_79 & _GEN_1130 | _GEN_3054 | _GEN_77 & _GEN_940)
      & (_GEN_2926
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_750 | _GEN_2798 | _GEN_73 & _GEN_560 | _GEN_2670 | _GEN_71
               & _GEN_370)
             & (_GEN_2542
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2446 & rob_predicated_2_11));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_12 <=
      ~(_GEN_79 & _GEN_1133 | _GEN_3055 | _GEN_77 & _GEN_943)
      & (_GEN_2927
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_753 | _GEN_2799 | _GEN_73 & _GEN_563 | _GEN_2671 | _GEN_71
               & _GEN_373)
             & (_GEN_2543
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2447 & rob_predicated_2_12));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_13 <=
      ~(_GEN_79 & _GEN_1136 | _GEN_3056 | _GEN_77 & _GEN_946)
      & (_GEN_2928
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_756 | _GEN_2800 | _GEN_73 & _GEN_566 | _GEN_2672 | _GEN_71
               & _GEN_376)
             & (_GEN_2544
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2448 & rob_predicated_2_13));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_14 <=
      ~(_GEN_79 & _GEN_1139 | _GEN_3057 | _GEN_77 & _GEN_949)
      & (_GEN_2929
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_759 | _GEN_2801 | _GEN_73 & _GEN_569 | _GEN_2673 | _GEN_71
               & _GEN_379)
             & (_GEN_2545
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2449 & rob_predicated_2_14));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_15 <=
      ~(_GEN_79 & _GEN_1142 | _GEN_3058 | _GEN_77 & _GEN_952)
      & (_GEN_2930
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_762 | _GEN_2802 | _GEN_73 & _GEN_572 | _GEN_2674 | _GEN_71
               & _GEN_382)
             & (_GEN_2546
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2450 & rob_predicated_2_15));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_16 <=
      ~(_GEN_79 & _GEN_1145 | _GEN_3059 | _GEN_77 & _GEN_955)
      & (_GEN_2931
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_765 | _GEN_2803 | _GEN_73 & _GEN_575 | _GEN_2675 | _GEN_71
               & _GEN_385)
             & (_GEN_2547
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2451 & rob_predicated_2_16));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_17 <=
      ~(_GEN_79 & _GEN_1148 | _GEN_3060 | _GEN_77 & _GEN_958)
      & (_GEN_2932
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_768 | _GEN_2804 | _GEN_73 & _GEN_578 | _GEN_2676 | _GEN_71
               & _GEN_388)
             & (_GEN_2548
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2452 & rob_predicated_2_17));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_18 <=
      ~(_GEN_79 & _GEN_1151 | _GEN_3061 | _GEN_77 & _GEN_961)
      & (_GEN_2933
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_771 | _GEN_2805 | _GEN_73 & _GEN_581 | _GEN_2677 | _GEN_71
               & _GEN_391)
             & (_GEN_2549
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2453 & rob_predicated_2_18));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_19 <=
      ~(_GEN_79 & _GEN_1154 | _GEN_3062 | _GEN_77 & _GEN_964)
      & (_GEN_2934
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_774 | _GEN_2806 | _GEN_73 & _GEN_584 | _GEN_2678 | _GEN_71
               & _GEN_394)
             & (_GEN_2550
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2454 & rob_predicated_2_19));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_20 <=
      ~(_GEN_79 & _GEN_1157 | _GEN_3063 | _GEN_77 & _GEN_967)
      & (_GEN_2935
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_777 | _GEN_2807 | _GEN_73 & _GEN_587 | _GEN_2679 | _GEN_71
               & _GEN_397)
             & (_GEN_2551
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2455 & rob_predicated_2_20));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_21 <=
      ~(_GEN_79 & _GEN_1160 | _GEN_3064 | _GEN_77 & _GEN_970)
      & (_GEN_2936
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_780 | _GEN_2808 | _GEN_73 & _GEN_590 | _GEN_2680 | _GEN_71
               & _GEN_400)
             & (_GEN_2552
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2456 & rob_predicated_2_21));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_22 <=
      ~(_GEN_79 & _GEN_1163 | _GEN_3065 | _GEN_77 & _GEN_973)
      & (_GEN_2937
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_783 | _GEN_2809 | _GEN_73 & _GEN_593 | _GEN_2681 | _GEN_71
               & _GEN_403)
             & (_GEN_2553
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2457 & rob_predicated_2_22));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_23 <=
      ~(_GEN_79 & _GEN_1166 | _GEN_3066 | _GEN_77 & _GEN_976)
      & (_GEN_2938
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_786 | _GEN_2810 | _GEN_73 & _GEN_596 | _GEN_2682 | _GEN_71
               & _GEN_406)
             & (_GEN_2554
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2458 & rob_predicated_2_23));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_24 <=
      ~(_GEN_79 & _GEN_1169 | _GEN_3067 | _GEN_77 & _GEN_979)
      & (_GEN_2939
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_789 | _GEN_2811 | _GEN_73 & _GEN_599 | _GEN_2683 | _GEN_71
               & _GEN_409)
             & (_GEN_2555
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2459 & rob_predicated_2_24));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_25 <=
      ~(_GEN_79 & _GEN_1172 | _GEN_3068 | _GEN_77 & _GEN_982)
      & (_GEN_2940
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_792 | _GEN_2812 | _GEN_73 & _GEN_602 | _GEN_2684 | _GEN_71
               & _GEN_412)
             & (_GEN_2556
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2460 & rob_predicated_2_25));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_26 <=
      ~(_GEN_79 & _GEN_1175 | _GEN_3069 | _GEN_77 & _GEN_985)
      & (_GEN_2941
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_795 | _GEN_2813 | _GEN_73 & _GEN_605 | _GEN_2685 | _GEN_71
               & _GEN_415)
             & (_GEN_2557
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2461 & rob_predicated_2_26));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_27 <=
      ~(_GEN_79 & _GEN_1178 | _GEN_3070 | _GEN_77 & _GEN_988)
      & (_GEN_2942
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_798 | _GEN_2814 | _GEN_73 & _GEN_608 | _GEN_2686 | _GEN_71
               & _GEN_418)
             & (_GEN_2558
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2462 & rob_predicated_2_27));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_28 <=
      ~(_GEN_79 & _GEN_1181 | _GEN_3071 | _GEN_77 & _GEN_991)
      & (_GEN_2943
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_801 | _GEN_2815 | _GEN_73 & _GEN_611 | _GEN_2687 | _GEN_71
               & _GEN_421)
             & (_GEN_2559
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2463 & rob_predicated_2_28));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_29 <=
      ~(_GEN_79 & _GEN_1184 | _GEN_3072 | _GEN_77 & _GEN_994)
      & (_GEN_2944
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_804 | _GEN_2816 | _GEN_73 & _GEN_614 | _GEN_2688 | _GEN_71
               & _GEN_424)
             & (_GEN_2560
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2464 & rob_predicated_2_29));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_30 <=
      ~(_GEN_79 & _GEN_1187 | _GEN_3073 | _GEN_77 & _GEN_997)
      & (_GEN_2945
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & _GEN_807 | _GEN_2817 | _GEN_73 & _GEN_617 | _GEN_2689 | _GEN_71
               & _GEN_427)
             & (_GEN_2561
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2465 & rob_predicated_2_30));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_31 <=
      ~(_GEN_79 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_3074 | _GEN_77
        & (&(io_wb_resps_7_bits_uop_rob_idx[6:2])))
      & (_GEN_2946
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_75 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2818 | _GEN_73
               & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_2690 | _GEN_71
               & (&(io_wb_resps_1_bits_uop_rob_idx[6:2])))
             & (_GEN_2562
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_2466 & rob_predicated_2_31));	// rob.scala:236:31, :268:25, :307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_bsy_3_0 <=
      ~_GEN_4131 & (_GEN_117 ? ~_GEN_4099 & _GEN_3972 : ~_GEN_4067 & _GEN_3972);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_1 <=
      ~_GEN_4132 & (_GEN_117 ? ~_GEN_4100 & _GEN_3974 : ~_GEN_4068 & _GEN_3974);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_2 <=
      ~_GEN_4133 & (_GEN_117 ? ~_GEN_4101 & _GEN_3976 : ~_GEN_4069 & _GEN_3976);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_3 <=
      ~_GEN_4134 & (_GEN_117 ? ~_GEN_4102 & _GEN_3978 : ~_GEN_4070 & _GEN_3978);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_4 <=
      ~_GEN_4135 & (_GEN_117 ? ~_GEN_4103 & _GEN_3980 : ~_GEN_4071 & _GEN_3980);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_5 <=
      ~_GEN_4136 & (_GEN_117 ? ~_GEN_4104 & _GEN_3982 : ~_GEN_4072 & _GEN_3982);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_6 <=
      ~_GEN_4137 & (_GEN_117 ? ~_GEN_4105 & _GEN_3984 : ~_GEN_4073 & _GEN_3984);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_7 <=
      ~_GEN_4138 & (_GEN_117 ? ~_GEN_4106 & _GEN_3986 : ~_GEN_4074 & _GEN_3986);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_8 <=
      ~_GEN_4139 & (_GEN_117 ? ~_GEN_4107 & _GEN_3988 : ~_GEN_4075 & _GEN_3988);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_9 <=
      ~_GEN_4140 & (_GEN_117 ? ~_GEN_4108 & _GEN_3990 : ~_GEN_4076 & _GEN_3990);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_10 <=
      ~_GEN_4141 & (_GEN_117 ? ~_GEN_4109 & _GEN_3992 : ~_GEN_4077 & _GEN_3992);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_11 <=
      ~_GEN_4142 & (_GEN_117 ? ~_GEN_4110 & _GEN_3994 : ~_GEN_4078 & _GEN_3994);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_12 <=
      ~_GEN_4143 & (_GEN_117 ? ~_GEN_4111 & _GEN_3996 : ~_GEN_4079 & _GEN_3996);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_13 <=
      ~_GEN_4144 & (_GEN_117 ? ~_GEN_4112 & _GEN_3998 : ~_GEN_4080 & _GEN_3998);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_14 <=
      ~_GEN_4145 & (_GEN_117 ? ~_GEN_4113 & _GEN_4000 : ~_GEN_4081 & _GEN_4000);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_15 <=
      ~_GEN_4146 & (_GEN_117 ? ~_GEN_4114 & _GEN_4002 : ~_GEN_4082 & _GEN_4002);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_16 <=
      ~_GEN_4147 & (_GEN_117 ? ~_GEN_4115 & _GEN_4004 : ~_GEN_4083 & _GEN_4004);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_17 <=
      ~_GEN_4148 & (_GEN_117 ? ~_GEN_4116 & _GEN_4006 : ~_GEN_4084 & _GEN_4006);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_18 <=
      ~_GEN_4149 & (_GEN_117 ? ~_GEN_4117 & _GEN_4008 : ~_GEN_4085 & _GEN_4008);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_19 <=
      ~_GEN_4150 & (_GEN_117 ? ~_GEN_4118 & _GEN_4010 : ~_GEN_4086 & _GEN_4010);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_20 <=
      ~_GEN_4151 & (_GEN_117 ? ~_GEN_4119 & _GEN_4012 : ~_GEN_4087 & _GEN_4012);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_21 <=
      ~_GEN_4152 & (_GEN_117 ? ~_GEN_4120 & _GEN_4014 : ~_GEN_4088 & _GEN_4014);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_22 <=
      ~_GEN_4153 & (_GEN_117 ? ~_GEN_4121 & _GEN_4016 : ~_GEN_4089 & _GEN_4016);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_23 <=
      ~_GEN_4154 & (_GEN_117 ? ~_GEN_4122 & _GEN_4018 : ~_GEN_4090 & _GEN_4018);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_24 <=
      ~_GEN_4155 & (_GEN_117 ? ~_GEN_4123 & _GEN_4020 : ~_GEN_4091 & _GEN_4020);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_25 <=
      ~_GEN_4156 & (_GEN_117 ? ~_GEN_4124 & _GEN_4022 : ~_GEN_4092 & _GEN_4022);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_26 <=
      ~_GEN_4157 & (_GEN_117 ? ~_GEN_4125 & _GEN_4024 : ~_GEN_4093 & _GEN_4024);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_27 <=
      ~_GEN_4158 & (_GEN_117 ? ~_GEN_4126 & _GEN_4026 : ~_GEN_4094 & _GEN_4026);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_28 <=
      ~_GEN_4159 & (_GEN_117 ? ~_GEN_4127 & _GEN_4028 : ~_GEN_4095 & _GEN_4028);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_29 <=
      ~_GEN_4160 & (_GEN_117 ? ~_GEN_4128 & _GEN_4030 : ~_GEN_4096 & _GEN_4030);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_30 <=
      ~_GEN_4161 & (_GEN_117 ? ~_GEN_4129 & _GEN_4032 : ~_GEN_4097 & _GEN_4032);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_bsy_3_31 <=
      ~_GEN_4162 & (_GEN_117 ? ~_GEN_4130 & _GEN_4034 : ~_GEN_4098 & _GEN_4034);	// rob.scala:308:28, :346:69, :347:31, :361:{31,75}, :363:26
    rob_unsafe_3_0 <=
      ~_GEN_4131 & (_GEN_117 ? ~_GEN_4099 & _GEN_4035 : ~_GEN_4067 & _GEN_4035);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_1 <=
      ~_GEN_4132 & (_GEN_117 ? ~_GEN_4100 & _GEN_4036 : ~_GEN_4068 & _GEN_4036);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_2 <=
      ~_GEN_4133 & (_GEN_117 ? ~_GEN_4101 & _GEN_4037 : ~_GEN_4069 & _GEN_4037);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_3 <=
      ~_GEN_4134 & (_GEN_117 ? ~_GEN_4102 & _GEN_4038 : ~_GEN_4070 & _GEN_4038);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_4 <=
      ~_GEN_4135 & (_GEN_117 ? ~_GEN_4103 & _GEN_4039 : ~_GEN_4071 & _GEN_4039);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_5 <=
      ~_GEN_4136 & (_GEN_117 ? ~_GEN_4104 & _GEN_4040 : ~_GEN_4072 & _GEN_4040);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_6 <=
      ~_GEN_4137 & (_GEN_117 ? ~_GEN_4105 & _GEN_4041 : ~_GEN_4073 & _GEN_4041);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_7 <=
      ~_GEN_4138 & (_GEN_117 ? ~_GEN_4106 & _GEN_4042 : ~_GEN_4074 & _GEN_4042);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_8 <=
      ~_GEN_4139 & (_GEN_117 ? ~_GEN_4107 & _GEN_4043 : ~_GEN_4075 & _GEN_4043);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_9 <=
      ~_GEN_4140 & (_GEN_117 ? ~_GEN_4108 & _GEN_4044 : ~_GEN_4076 & _GEN_4044);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_10 <=
      ~_GEN_4141 & (_GEN_117 ? ~_GEN_4109 & _GEN_4045 : ~_GEN_4077 & _GEN_4045);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_11 <=
      ~_GEN_4142 & (_GEN_117 ? ~_GEN_4110 & _GEN_4046 : ~_GEN_4078 & _GEN_4046);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_12 <=
      ~_GEN_4143 & (_GEN_117 ? ~_GEN_4111 & _GEN_4047 : ~_GEN_4079 & _GEN_4047);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_13 <=
      ~_GEN_4144 & (_GEN_117 ? ~_GEN_4112 & _GEN_4048 : ~_GEN_4080 & _GEN_4048);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_14 <=
      ~_GEN_4145 & (_GEN_117 ? ~_GEN_4113 & _GEN_4049 : ~_GEN_4081 & _GEN_4049);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_15 <=
      ~_GEN_4146 & (_GEN_117 ? ~_GEN_4114 & _GEN_4050 : ~_GEN_4082 & _GEN_4050);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_16 <=
      ~_GEN_4147 & (_GEN_117 ? ~_GEN_4115 & _GEN_4051 : ~_GEN_4083 & _GEN_4051);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_17 <=
      ~_GEN_4148 & (_GEN_117 ? ~_GEN_4116 & _GEN_4052 : ~_GEN_4084 & _GEN_4052);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_18 <=
      ~_GEN_4149 & (_GEN_117 ? ~_GEN_4117 & _GEN_4053 : ~_GEN_4085 & _GEN_4053);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_19 <=
      ~_GEN_4150 & (_GEN_117 ? ~_GEN_4118 & _GEN_4054 : ~_GEN_4086 & _GEN_4054);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_20 <=
      ~_GEN_4151 & (_GEN_117 ? ~_GEN_4119 & _GEN_4055 : ~_GEN_4087 & _GEN_4055);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_21 <=
      ~_GEN_4152 & (_GEN_117 ? ~_GEN_4120 & _GEN_4056 : ~_GEN_4088 & _GEN_4056);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_22 <=
      ~_GEN_4153 & (_GEN_117 ? ~_GEN_4121 & _GEN_4057 : ~_GEN_4089 & _GEN_4057);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_23 <=
      ~_GEN_4154 & (_GEN_117 ? ~_GEN_4122 & _GEN_4058 : ~_GEN_4090 & _GEN_4058);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_24 <=
      ~_GEN_4155 & (_GEN_117 ? ~_GEN_4123 & _GEN_4059 : ~_GEN_4091 & _GEN_4059);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_25 <=
      ~_GEN_4156 & (_GEN_117 ? ~_GEN_4124 & _GEN_4060 : ~_GEN_4092 & _GEN_4060);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_26 <=
      ~_GEN_4157 & (_GEN_117 ? ~_GEN_4125 & _GEN_4061 : ~_GEN_4093 & _GEN_4061);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_27 <=
      ~_GEN_4158 & (_GEN_117 ? ~_GEN_4126 & _GEN_4062 : ~_GEN_4094 & _GEN_4062);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_28 <=
      ~_GEN_4159 & (_GEN_117 ? ~_GEN_4127 & _GEN_4063 : ~_GEN_4095 & _GEN_4063);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_29 <=
      ~_GEN_4160 & (_GEN_117 ? ~_GEN_4128 & _GEN_4064 : ~_GEN_4096 & _GEN_4064);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_30 <=
      ~_GEN_4161 & (_GEN_117 ? ~_GEN_4129 & _GEN_4065 : ~_GEN_4097 & _GEN_4065);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    rob_unsafe_3_31 <=
      ~_GEN_4162 & (_GEN_117 ? ~_GEN_4130 & _GEN_4066 : ~_GEN_4098 & _GEN_4066);	// rob.scala:309:28, :346:69, :348:31, :361:{31,75}, :363:26, :364:26
    if (_GEN_3331) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_0_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_0_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_0_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_0_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_0_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_0_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_0_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_0_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_0_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_0_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_0_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_0_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_0_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_0_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_0_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_0_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4195) | ~rob_val_3_0) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3331)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_0_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_0_br_mask <= rob_uop_3_0_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3332) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_1_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_1_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_1_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_1_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_1_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_1_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_1_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_1_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_1_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_1_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_1_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_1_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_1_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_1_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_1_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_1_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4196) | ~rob_val_3_1) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3332)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_1_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_1_br_mask <= rob_uop_3_1_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3333) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_2_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_2_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_2_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_2_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_2_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_2_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_2_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_2_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_2_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_2_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_2_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_2_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_2_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_2_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_2_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_2_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4197) | ~rob_val_3_2) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3333)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_2_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_2_br_mask <= rob_uop_3_2_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3334) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_3_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_3_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_3_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_3_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_3_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_3_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_3_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_3_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_3_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_3_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_3_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_3_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_3_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_3_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_3_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_3_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4198) | ~rob_val_3_3) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3334)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_3_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_3_br_mask <= rob_uop_3_3_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3335) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_4_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_4_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_4_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_4_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_4_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_4_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_4_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_4_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_4_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_4_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_4_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_4_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_4_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_4_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_4_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_4_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4199) | ~rob_val_3_4) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3335)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_4_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_4_br_mask <= rob_uop_3_4_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3336) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_5_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_5_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_5_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_5_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_5_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_5_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_5_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_5_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_5_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_5_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_5_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_5_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_5_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_5_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_5_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_5_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4200) | ~rob_val_3_5) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3336)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_5_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_5_br_mask <= rob_uop_3_5_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3337) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_6_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_6_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_6_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_6_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_6_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_6_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_6_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_6_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_6_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_6_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_6_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_6_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_6_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_6_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_6_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_6_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4201) | ~rob_val_3_6) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3337)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_6_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_6_br_mask <= rob_uop_3_6_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3338) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_7_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_7_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_7_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_7_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_7_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_7_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_7_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_7_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_7_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_7_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_7_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_7_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_7_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_7_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_7_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_7_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4202) | ~rob_val_3_7) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3338)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_7_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_7_br_mask <= rob_uop_3_7_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3339) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_8_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_8_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_8_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_8_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_8_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_8_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_8_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_8_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_8_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_8_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_8_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_8_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_8_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_8_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_8_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_8_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4203) | ~rob_val_3_8) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3339)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_8_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_8_br_mask <= rob_uop_3_8_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3340) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_9_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_9_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_9_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_9_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_9_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_9_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_9_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_9_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_9_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_9_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_9_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_9_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_9_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_9_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_9_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_9_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4204) | ~rob_val_3_9) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3340)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_9_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_9_br_mask <= rob_uop_3_9_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3341) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_10_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_10_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_10_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_10_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_10_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_10_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_10_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_10_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_10_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_10_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_10_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_10_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_10_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_10_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_10_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_10_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4205) | ~rob_val_3_10) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3341)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_10_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_10_br_mask <= rob_uop_3_10_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3342) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_11_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_11_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_11_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_11_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_11_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_11_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_11_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_11_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_11_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_11_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_11_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_11_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_11_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_11_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_11_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_11_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4206) | ~rob_val_3_11) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3342)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_11_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_11_br_mask <= rob_uop_3_11_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3343) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_12_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_12_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_12_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_12_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_12_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_12_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_12_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_12_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_12_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_12_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_12_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_12_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_12_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_12_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_12_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_12_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4207) | ~rob_val_3_12) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3343)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_12_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_12_br_mask <= rob_uop_3_12_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3344) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_13_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_13_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_13_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_13_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_13_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_13_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_13_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_13_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_13_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_13_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_13_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_13_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_13_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_13_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_13_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_13_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4208) | ~rob_val_3_13) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3344)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_13_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_13_br_mask <= rob_uop_3_13_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3345) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_14_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_14_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_14_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_14_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_14_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_14_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_14_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_14_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_14_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_14_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_14_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_14_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_14_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_14_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_14_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_14_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4209) | ~rob_val_3_14) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3345)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_14_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_14_br_mask <= rob_uop_3_14_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3346) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_15_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_15_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_15_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_15_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_15_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_15_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_15_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_15_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_15_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_15_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_15_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_15_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_15_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_15_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_15_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_15_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4210) | ~rob_val_3_15) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3346)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_15_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_15_br_mask <= rob_uop_3_15_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3347) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_16_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_16_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_16_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_16_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_16_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_16_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_16_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_16_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_16_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_16_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_16_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_16_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_16_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_16_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_16_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_16_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4211) | ~rob_val_3_16) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3347)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_16_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_16_br_mask <= rob_uop_3_16_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3348) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_17_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_17_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_17_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_17_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_17_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_17_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_17_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_17_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_17_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_17_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_17_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_17_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_17_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_17_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_17_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_17_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4212) | ~rob_val_3_17) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3348)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_17_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_17_br_mask <= rob_uop_3_17_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3349) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_18_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_18_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_18_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_18_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_18_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_18_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_18_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_18_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_18_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_18_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_18_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_18_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_18_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_18_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_18_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_18_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4213) | ~rob_val_3_18) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3349)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_18_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_18_br_mask <= rob_uop_3_18_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3350) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_19_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_19_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_19_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_19_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_19_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_19_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_19_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_19_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_19_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_19_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_19_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_19_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_19_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_19_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_19_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_19_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4214) | ~rob_val_3_19) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3350)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_19_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_19_br_mask <= rob_uop_3_19_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3351) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_20_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_20_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_20_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_20_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_20_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_20_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_20_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_20_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_20_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_20_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_20_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_20_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_20_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_20_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_20_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_20_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4215) | ~rob_val_3_20) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3351)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_20_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_20_br_mask <= rob_uop_3_20_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3352) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_21_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_21_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_21_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_21_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_21_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_21_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_21_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_21_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_21_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_21_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_21_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_21_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_21_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_21_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_21_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_21_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4216) | ~rob_val_3_21) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3352)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_21_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_21_br_mask <= rob_uop_3_21_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3353) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_22_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_22_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_22_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_22_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_22_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_22_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_22_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_22_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_22_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_22_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_22_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_22_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_22_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_22_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_22_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_22_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4217) | ~rob_val_3_22) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3353)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_22_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_22_br_mask <= rob_uop_3_22_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3354) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_23_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_23_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_23_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_23_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_23_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_23_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_23_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_23_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_23_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_23_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_23_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_23_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_23_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_23_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_23_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_23_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4218) | ~rob_val_3_23) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3354)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_23_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_23_br_mask <= rob_uop_3_23_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3355) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_24_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_24_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_24_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_24_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_24_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_24_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_24_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_24_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_24_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_24_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_24_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_24_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_24_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_24_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_24_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_24_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4219) | ~rob_val_3_24) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3355)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_24_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_24_br_mask <= rob_uop_3_24_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3356) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_25_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_25_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_25_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_25_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_25_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_25_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_25_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_25_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_25_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_25_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_25_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_25_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_25_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_25_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_25_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_25_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4220) | ~rob_val_3_25) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3356)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_25_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_25_br_mask <= rob_uop_3_25_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3357) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_26_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_26_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_26_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_26_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_26_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_26_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_26_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_26_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_26_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_26_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_26_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_26_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_26_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_26_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_26_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_26_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4221) | ~rob_val_3_26) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3357)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_26_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_26_br_mask <= rob_uop_3_26_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3358) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_27_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_27_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_27_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_27_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_27_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_27_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_27_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_27_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_27_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_27_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_27_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_27_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_27_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_27_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_27_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_27_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4222) | ~rob_val_3_27) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3358)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_27_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_27_br_mask <= rob_uop_3_27_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3359) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_28_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_28_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_28_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_28_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_28_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_28_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_28_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_28_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_28_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_28_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_28_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_28_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_28_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_28_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_28_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_28_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4223) | ~rob_val_3_28) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3359)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_28_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_28_br_mask <= rob_uop_3_28_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3360) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_29_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_29_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_29_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_29_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_29_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_29_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_29_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_29_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_29_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_29_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_29_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_29_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_29_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_29_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_29_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_29_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4224) | ~rob_val_3_29) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3360)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_29_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_29_br_mask <= rob_uop_3_29_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3361) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_30_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_30_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_30_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_30_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_30_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_30_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_30_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_30_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_30_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_30_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_30_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_30_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_30_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_30_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_30_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_30_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4225) | ~rob_val_3_30) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3361)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_30_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_30_br_mask <= rob_uop_3_30_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_3362) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_31_uopc <= io_enq_uops_3_uopc;	// rob.scala:310:28
      rob_uop_3_31_is_rvc <= io_enq_uops_3_is_rvc;	// rob.scala:310:28
      rob_uop_3_31_ftq_idx <= io_enq_uops_3_ftq_idx;	// rob.scala:310:28
      rob_uop_3_31_edge_inst <= io_enq_uops_3_edge_inst;	// rob.scala:310:28
      rob_uop_3_31_pc_lob <= io_enq_uops_3_pc_lob;	// rob.scala:310:28
      rob_uop_3_31_pdst <= io_enq_uops_3_pdst;	// rob.scala:310:28
      rob_uop_3_31_stale_pdst <= io_enq_uops_3_stale_pdst;	// rob.scala:310:28
      rob_uop_3_31_is_fencei <= io_enq_uops_3_is_fencei;	// rob.scala:310:28
      rob_uop_3_31_uses_ldq <= io_enq_uops_3_uses_ldq;	// rob.scala:310:28
      rob_uop_3_31_uses_stq <= io_enq_uops_3_uses_stq;	// rob.scala:310:28
      rob_uop_3_31_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_31_flush_on_commit <= io_enq_uops_3_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_31_ldst <= io_enq_uops_3_ldst;	// rob.scala:310:28
      rob_uop_3_31_ldst_val <= io_enq_uops_3_ldst_val;	// rob.scala:310:28
      rob_uop_3_31_dst_rtype <= io_enq_uops_3_dst_rtype;	// rob.scala:310:28
      rob_uop_3_31_fp_val <= io_enq_uops_3_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_4226) | ~rob_val_3_31) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_3362)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_31_br_mask <= io_enq_uops_3_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_31_br_mask <= rob_uop_3_31_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    rob_exception_3_0 <=
      ~_GEN_4163
      & (_GEN_119 & _GEN_1413
         | (_GEN_3331 ? io_enq_uops_3_exception : rob_exception_3_0));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_1 <=
      ~_GEN_4164
      & (_GEN_119 & _GEN_1414
         | (_GEN_3332 ? io_enq_uops_3_exception : rob_exception_3_1));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_2 <=
      ~_GEN_4165
      & (_GEN_119 & _GEN_1415
         | (_GEN_3333 ? io_enq_uops_3_exception : rob_exception_3_2));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_3 <=
      ~_GEN_4166
      & (_GEN_119 & _GEN_1416
         | (_GEN_3334 ? io_enq_uops_3_exception : rob_exception_3_3));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_4 <=
      ~_GEN_4167
      & (_GEN_119 & _GEN_1417
         | (_GEN_3335 ? io_enq_uops_3_exception : rob_exception_3_4));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_5 <=
      ~_GEN_4168
      & (_GEN_119 & _GEN_1418
         | (_GEN_3336 ? io_enq_uops_3_exception : rob_exception_3_5));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_6 <=
      ~_GEN_4169
      & (_GEN_119 & _GEN_1419
         | (_GEN_3337 ? io_enq_uops_3_exception : rob_exception_3_6));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_7 <=
      ~_GEN_4170
      & (_GEN_119 & _GEN_1420
         | (_GEN_3338 ? io_enq_uops_3_exception : rob_exception_3_7));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_8 <=
      ~_GEN_4171
      & (_GEN_119 & _GEN_1421
         | (_GEN_3339 ? io_enq_uops_3_exception : rob_exception_3_8));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_9 <=
      ~_GEN_4172
      & (_GEN_119 & _GEN_1422
         | (_GEN_3340 ? io_enq_uops_3_exception : rob_exception_3_9));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_10 <=
      ~_GEN_4173
      & (_GEN_119 & _GEN_1423
         | (_GEN_3341 ? io_enq_uops_3_exception : rob_exception_3_10));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_11 <=
      ~_GEN_4174
      & (_GEN_119 & _GEN_1424
         | (_GEN_3342 ? io_enq_uops_3_exception : rob_exception_3_11));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_12 <=
      ~_GEN_4175
      & (_GEN_119 & _GEN_1425
         | (_GEN_3343 ? io_enq_uops_3_exception : rob_exception_3_12));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_13 <=
      ~_GEN_4176
      & (_GEN_119 & _GEN_1426
         | (_GEN_3344 ? io_enq_uops_3_exception : rob_exception_3_13));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_14 <=
      ~_GEN_4177
      & (_GEN_119 & _GEN_1427
         | (_GEN_3345 ? io_enq_uops_3_exception : rob_exception_3_14));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_15 <=
      ~_GEN_4178
      & (_GEN_119 & _GEN_1428
         | (_GEN_3346 ? io_enq_uops_3_exception : rob_exception_3_15));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_16 <=
      ~_GEN_4179
      & (_GEN_119 & _GEN_1429
         | (_GEN_3347 ? io_enq_uops_3_exception : rob_exception_3_16));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_17 <=
      ~_GEN_4180
      & (_GEN_119 & _GEN_1430
         | (_GEN_3348 ? io_enq_uops_3_exception : rob_exception_3_17));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_18 <=
      ~_GEN_4181
      & (_GEN_119 & _GEN_1431
         | (_GEN_3349 ? io_enq_uops_3_exception : rob_exception_3_18));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_19 <=
      ~_GEN_4182
      & (_GEN_119 & _GEN_1432
         | (_GEN_3350 ? io_enq_uops_3_exception : rob_exception_3_19));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_20 <=
      ~_GEN_4183
      & (_GEN_119 & _GEN_1433
         | (_GEN_3351 ? io_enq_uops_3_exception : rob_exception_3_20));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_21 <=
      ~_GEN_4184
      & (_GEN_119 & _GEN_1434
         | (_GEN_3352 ? io_enq_uops_3_exception : rob_exception_3_21));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_22 <=
      ~_GEN_4185
      & (_GEN_119 & _GEN_1435
         | (_GEN_3353 ? io_enq_uops_3_exception : rob_exception_3_22));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_23 <=
      ~_GEN_4186
      & (_GEN_119 & _GEN_1436
         | (_GEN_3354 ? io_enq_uops_3_exception : rob_exception_3_23));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_24 <=
      ~_GEN_4187
      & (_GEN_119 & _GEN_1437
         | (_GEN_3355 ? io_enq_uops_3_exception : rob_exception_3_24));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_25 <=
      ~_GEN_4188
      & (_GEN_119 & _GEN_1438
         | (_GEN_3356 ? io_enq_uops_3_exception : rob_exception_3_25));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_26 <=
      ~_GEN_4189
      & (_GEN_119 & _GEN_1439
         | (_GEN_3357 ? io_enq_uops_3_exception : rob_exception_3_26));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_27 <=
      ~_GEN_4190
      & (_GEN_119 & _GEN_1440
         | (_GEN_3358 ? io_enq_uops_3_exception : rob_exception_3_27));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_28 <=
      ~_GEN_4191
      & (_GEN_119 & _GEN_1441
         | (_GEN_3359 ? io_enq_uops_3_exception : rob_exception_3_28));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_29 <=
      ~_GEN_4192
      & (_GEN_119 & _GEN_1442
         | (_GEN_3360 ? io_enq_uops_3_exception : rob_exception_3_29));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_30 <=
      ~_GEN_4193
      & (_GEN_119 & _GEN_1443
         | (_GEN_3361 ? io_enq_uops_3_exception : rob_exception_3_30));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3_31 <=
      ~_GEN_4194
      & (_GEN_119 & (&(io_lxcpt_bits_uop_rob_idx[6:2]))
         | (_GEN_3362 ? io_enq_uops_3_exception : rob_exception_3_31));	// rob.scala:236:31, :268:25, :307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_predicated_3_0 <=
      ~(_GEN_114 & _GEN_1097 | _GEN_3939 | _GEN_112 & _GEN_907)
      & (_GEN_3811
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_717 | _GEN_3683 | _GEN_108 & _GEN_527 | _GEN_3555
               | _GEN_106 & _GEN_337)
             & (_GEN_3427
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3331 & rob_predicated_3_0));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_1 <=
      ~(_GEN_114 & _GEN_1100 | _GEN_3940 | _GEN_112 & _GEN_910)
      & (_GEN_3812
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_720 | _GEN_3684 | _GEN_108 & _GEN_530 | _GEN_3556
               | _GEN_106 & _GEN_340)
             & (_GEN_3428
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3332 & rob_predicated_3_1));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_2 <=
      ~(_GEN_114 & _GEN_1103 | _GEN_3941 | _GEN_112 & _GEN_913)
      & (_GEN_3813
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_723 | _GEN_3685 | _GEN_108 & _GEN_533 | _GEN_3557
               | _GEN_106 & _GEN_343)
             & (_GEN_3429
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3333 & rob_predicated_3_2));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_3 <=
      ~(_GEN_114 & _GEN_1106 | _GEN_3942 | _GEN_112 & _GEN_916)
      & (_GEN_3814
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_726 | _GEN_3686 | _GEN_108 & _GEN_536 | _GEN_3558
               | _GEN_106 & _GEN_346)
             & (_GEN_3430
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3334 & rob_predicated_3_3));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_4 <=
      ~(_GEN_114 & _GEN_1109 | _GEN_3943 | _GEN_112 & _GEN_919)
      & (_GEN_3815
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_729 | _GEN_3687 | _GEN_108 & _GEN_539 | _GEN_3559
               | _GEN_106 & _GEN_349)
             & (_GEN_3431
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3335 & rob_predicated_3_4));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_5 <=
      ~(_GEN_114 & _GEN_1112 | _GEN_3944 | _GEN_112 & _GEN_922)
      & (_GEN_3816
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_732 | _GEN_3688 | _GEN_108 & _GEN_542 | _GEN_3560
               | _GEN_106 & _GEN_352)
             & (_GEN_3432
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3336 & rob_predicated_3_5));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_6 <=
      ~(_GEN_114 & _GEN_1115 | _GEN_3945 | _GEN_112 & _GEN_925)
      & (_GEN_3817
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_735 | _GEN_3689 | _GEN_108 & _GEN_545 | _GEN_3561
               | _GEN_106 & _GEN_355)
             & (_GEN_3433
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3337 & rob_predicated_3_6));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_7 <=
      ~(_GEN_114 & _GEN_1118 | _GEN_3946 | _GEN_112 & _GEN_928)
      & (_GEN_3818
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_738 | _GEN_3690 | _GEN_108 & _GEN_548 | _GEN_3562
               | _GEN_106 & _GEN_358)
             & (_GEN_3434
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3338 & rob_predicated_3_7));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_8 <=
      ~(_GEN_114 & _GEN_1121 | _GEN_3947 | _GEN_112 & _GEN_931)
      & (_GEN_3819
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_741 | _GEN_3691 | _GEN_108 & _GEN_551 | _GEN_3563
               | _GEN_106 & _GEN_361)
             & (_GEN_3435
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3339 & rob_predicated_3_8));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_9 <=
      ~(_GEN_114 & _GEN_1124 | _GEN_3948 | _GEN_112 & _GEN_934)
      & (_GEN_3820
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_744 | _GEN_3692 | _GEN_108 & _GEN_554 | _GEN_3564
               | _GEN_106 & _GEN_364)
             & (_GEN_3436
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3340 & rob_predicated_3_9));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_10 <=
      ~(_GEN_114 & _GEN_1127 | _GEN_3949 | _GEN_112 & _GEN_937)
      & (_GEN_3821
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_747 | _GEN_3693 | _GEN_108 & _GEN_557 | _GEN_3565
               | _GEN_106 & _GEN_367)
             & (_GEN_3437
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3341 & rob_predicated_3_10));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_11 <=
      ~(_GEN_114 & _GEN_1130 | _GEN_3950 | _GEN_112 & _GEN_940)
      & (_GEN_3822
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_750 | _GEN_3694 | _GEN_108 & _GEN_560 | _GEN_3566
               | _GEN_106 & _GEN_370)
             & (_GEN_3438
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3342 & rob_predicated_3_11));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_12 <=
      ~(_GEN_114 & _GEN_1133 | _GEN_3951 | _GEN_112 & _GEN_943)
      & (_GEN_3823
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_753 | _GEN_3695 | _GEN_108 & _GEN_563 | _GEN_3567
               | _GEN_106 & _GEN_373)
             & (_GEN_3439
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3343 & rob_predicated_3_12));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_13 <=
      ~(_GEN_114 & _GEN_1136 | _GEN_3952 | _GEN_112 & _GEN_946)
      & (_GEN_3824
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_756 | _GEN_3696 | _GEN_108 & _GEN_566 | _GEN_3568
               | _GEN_106 & _GEN_376)
             & (_GEN_3440
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3344 & rob_predicated_3_13));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_14 <=
      ~(_GEN_114 & _GEN_1139 | _GEN_3953 | _GEN_112 & _GEN_949)
      & (_GEN_3825
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_759 | _GEN_3697 | _GEN_108 & _GEN_569 | _GEN_3569
               | _GEN_106 & _GEN_379)
             & (_GEN_3441
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3345 & rob_predicated_3_14));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_15 <=
      ~(_GEN_114 & _GEN_1142 | _GEN_3954 | _GEN_112 & _GEN_952)
      & (_GEN_3826
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_762 | _GEN_3698 | _GEN_108 & _GEN_572 | _GEN_3570
               | _GEN_106 & _GEN_382)
             & (_GEN_3442
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3346 & rob_predicated_3_15));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_16 <=
      ~(_GEN_114 & _GEN_1145 | _GEN_3955 | _GEN_112 & _GEN_955)
      & (_GEN_3827
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_765 | _GEN_3699 | _GEN_108 & _GEN_575 | _GEN_3571
               | _GEN_106 & _GEN_385)
             & (_GEN_3443
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3347 & rob_predicated_3_16));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_17 <=
      ~(_GEN_114 & _GEN_1148 | _GEN_3956 | _GEN_112 & _GEN_958)
      & (_GEN_3828
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_768 | _GEN_3700 | _GEN_108 & _GEN_578 | _GEN_3572
               | _GEN_106 & _GEN_388)
             & (_GEN_3444
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3348 & rob_predicated_3_17));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_18 <=
      ~(_GEN_114 & _GEN_1151 | _GEN_3957 | _GEN_112 & _GEN_961)
      & (_GEN_3829
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_771 | _GEN_3701 | _GEN_108 & _GEN_581 | _GEN_3573
               | _GEN_106 & _GEN_391)
             & (_GEN_3445
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3349 & rob_predicated_3_18));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_19 <=
      ~(_GEN_114 & _GEN_1154 | _GEN_3958 | _GEN_112 & _GEN_964)
      & (_GEN_3830
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_774 | _GEN_3702 | _GEN_108 & _GEN_584 | _GEN_3574
               | _GEN_106 & _GEN_394)
             & (_GEN_3446
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3350 & rob_predicated_3_19));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_20 <=
      ~(_GEN_114 & _GEN_1157 | _GEN_3959 | _GEN_112 & _GEN_967)
      & (_GEN_3831
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_777 | _GEN_3703 | _GEN_108 & _GEN_587 | _GEN_3575
               | _GEN_106 & _GEN_397)
             & (_GEN_3447
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3351 & rob_predicated_3_20));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_21 <=
      ~(_GEN_114 & _GEN_1160 | _GEN_3960 | _GEN_112 & _GEN_970)
      & (_GEN_3832
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_780 | _GEN_3704 | _GEN_108 & _GEN_590 | _GEN_3576
               | _GEN_106 & _GEN_400)
             & (_GEN_3448
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3352 & rob_predicated_3_21));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_22 <=
      ~(_GEN_114 & _GEN_1163 | _GEN_3961 | _GEN_112 & _GEN_973)
      & (_GEN_3833
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_783 | _GEN_3705 | _GEN_108 & _GEN_593 | _GEN_3577
               | _GEN_106 & _GEN_403)
             & (_GEN_3449
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3353 & rob_predicated_3_22));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_23 <=
      ~(_GEN_114 & _GEN_1166 | _GEN_3962 | _GEN_112 & _GEN_976)
      & (_GEN_3834
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_786 | _GEN_3706 | _GEN_108 & _GEN_596 | _GEN_3578
               | _GEN_106 & _GEN_406)
             & (_GEN_3450
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3354 & rob_predicated_3_23));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_24 <=
      ~(_GEN_114 & _GEN_1169 | _GEN_3963 | _GEN_112 & _GEN_979)
      & (_GEN_3835
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_789 | _GEN_3707 | _GEN_108 & _GEN_599 | _GEN_3579
               | _GEN_106 & _GEN_409)
             & (_GEN_3451
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3355 & rob_predicated_3_24));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_25 <=
      ~(_GEN_114 & _GEN_1172 | _GEN_3964 | _GEN_112 & _GEN_982)
      & (_GEN_3836
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_792 | _GEN_3708 | _GEN_108 & _GEN_602 | _GEN_3580
               | _GEN_106 & _GEN_412)
             & (_GEN_3452
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3356 & rob_predicated_3_25));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_26 <=
      ~(_GEN_114 & _GEN_1175 | _GEN_3965 | _GEN_112 & _GEN_985)
      & (_GEN_3837
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_795 | _GEN_3709 | _GEN_108 & _GEN_605 | _GEN_3581
               | _GEN_106 & _GEN_415)
             & (_GEN_3453
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3357 & rob_predicated_3_26));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_27 <=
      ~(_GEN_114 & _GEN_1178 | _GEN_3966 | _GEN_112 & _GEN_988)
      & (_GEN_3838
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_798 | _GEN_3710 | _GEN_108 & _GEN_608 | _GEN_3582
               | _GEN_106 & _GEN_418)
             & (_GEN_3454
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3358 & rob_predicated_3_27));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_28 <=
      ~(_GEN_114 & _GEN_1181 | _GEN_3967 | _GEN_112 & _GEN_991)
      & (_GEN_3839
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_801 | _GEN_3711 | _GEN_108 & _GEN_611 | _GEN_3583
               | _GEN_106 & _GEN_421)
             & (_GEN_3455
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3359 & rob_predicated_3_28));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_29 <=
      ~(_GEN_114 & _GEN_1184 | _GEN_3968 | _GEN_112 & _GEN_994)
      & (_GEN_3840
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_804 | _GEN_3712 | _GEN_108 & _GEN_614 | _GEN_3584
               | _GEN_106 & _GEN_424)
             & (_GEN_3456
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3360 & rob_predicated_3_29));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_30 <=
      ~(_GEN_114 & _GEN_1187 | _GEN_3969 | _GEN_112 & _GEN_997)
      & (_GEN_3841
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & _GEN_807 | _GEN_3713 | _GEN_108 & _GEN_617 | _GEN_3585
               | _GEN_106 & _GEN_427)
             & (_GEN_3457
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3361 & rob_predicated_3_30));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3_31 <=
      ~(_GEN_114 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_3970 | _GEN_112
        & (&(io_wb_resps_7_bits_uop_rob_idx[6:2])))
      & (_GEN_3842
           ? io_wb_resps_6_bits_predicated
           : ~(_GEN_110 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_3714 | _GEN_108
               & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_3586 | _GEN_106
               & (&(io_wb_resps_1_bits_uop_rob_idx[6:2])))
             & (_GEN_3458
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_3362 & rob_predicated_3_31));	// rob.scala:236:31, :268:25, :307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    block_commit_REG <= exception_thrown;	// rob.scala:540:94, :545:85
    block_commit_REG_1 <= exception_thrown;	// rob.scala:540:131, :545:85
    block_commit_REG_2 <= block_commit_REG_1;	// rob.scala:540:{123,131}
    REG <= exception_thrown;	// rob.scala:545:85, :808:30
    REG_1 <= REG;	// rob.scala:808:{22,30}
    REG_2 <= exception_thrown;	// rob.scala:545:85, :824:22
    _GEN_4231 =
      {{_GEN_131[rob_head]},
       {_GEN_96[rob_head]},
       {_GEN_61[rob_head]},
       {_GEN_26[rob_head]}};	// rob.scala:224:29, :411:25, :484:26, :865:98
    io_com_load_is_at_rob_head_REG <=
      _GEN_4231[rob_head_vals_0
                  ? 2'h0
                  : rob_head_vals_1 ? 2'h1 : {1'h1, ~rob_head_vals_2}]
      & ~(will_commit_0 | will_commit_1 | will_commit_2 | will_commit_3);	// Mux.scala:47:69, rob.scala:221:26, :398:49, :540:33, :547:70, :865:{40,98}, :866:{41,62}
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:1703];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [10:0] i = 11'h0; i < 11'h6A8; i += 11'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        rob_state = _RANDOM[11'h0][1:0];	// rob.scala:221:26
        rob_head = _RANDOM[11'h0][6:2];	// rob.scala:221:26, :224:29
        rob_head_lsb = _RANDOM[11'h0][8:7];	// rob.scala:221:26, :225:29
        rob_tail = _RANDOM[11'h0][13:9];	// rob.scala:221:26, :228:29
        rob_tail_lsb = _RANDOM[11'h0][15:14];	// rob.scala:221:26, :229:29
        rob_pnr = _RANDOM[11'h0][20:16];	// rob.scala:221:26, :232:29
        rob_pnr_lsb = _RANDOM[11'h0][22:21];	// rob.scala:221:26, :233:29
        maybe_full = _RANDOM[11'h0][23];	// rob.scala:221:26, :239:29
        r_xcpt_val = _RANDOM[11'h0][24];	// rob.scala:221:26, :258:33
        r_xcpt_uop_br_mask = {_RANDOM[11'h5][31:21], _RANDOM[11'h6][8:0]};	// rob.scala:259:29
        r_xcpt_uop_rob_idx = {_RANDOM[11'h7][31:28], _RANDOM[11'h8][2:0]};	// rob.scala:259:29
        r_xcpt_uop_exc_cause =
          {_RANDOM[11'h9][31:29], _RANDOM[11'hA], _RANDOM[11'hB][28:0]};	// rob.scala:259:29
        r_xcpt_badvaddr = {_RANDOM[11'hD][31:26], _RANDOM[11'hE], _RANDOM[11'hF][1:0]};	// rob.scala:260:29
        rob_val_0 = _RANDOM[11'hF][2];	// rob.scala:260:29, :307:32
        rob_val_1 = _RANDOM[11'hF][3];	// rob.scala:260:29, :307:32
        rob_val_2 = _RANDOM[11'hF][4];	// rob.scala:260:29, :307:32
        rob_val_3 = _RANDOM[11'hF][5];	// rob.scala:260:29, :307:32
        rob_val_4 = _RANDOM[11'hF][6];	// rob.scala:260:29, :307:32
        rob_val_5 = _RANDOM[11'hF][7];	// rob.scala:260:29, :307:32
        rob_val_6 = _RANDOM[11'hF][8];	// rob.scala:260:29, :307:32
        rob_val_7 = _RANDOM[11'hF][9];	// rob.scala:260:29, :307:32
        rob_val_8 = _RANDOM[11'hF][10];	// rob.scala:260:29, :307:32
        rob_val_9 = _RANDOM[11'hF][11];	// rob.scala:260:29, :307:32
        rob_val_10 = _RANDOM[11'hF][12];	// rob.scala:260:29, :307:32
        rob_val_11 = _RANDOM[11'hF][13];	// rob.scala:260:29, :307:32
        rob_val_12 = _RANDOM[11'hF][14];	// rob.scala:260:29, :307:32
        rob_val_13 = _RANDOM[11'hF][15];	// rob.scala:260:29, :307:32
        rob_val_14 = _RANDOM[11'hF][16];	// rob.scala:260:29, :307:32
        rob_val_15 = _RANDOM[11'hF][17];	// rob.scala:260:29, :307:32
        rob_val_16 = _RANDOM[11'hF][18];	// rob.scala:260:29, :307:32
        rob_val_17 = _RANDOM[11'hF][19];	// rob.scala:260:29, :307:32
        rob_val_18 = _RANDOM[11'hF][20];	// rob.scala:260:29, :307:32
        rob_val_19 = _RANDOM[11'hF][21];	// rob.scala:260:29, :307:32
        rob_val_20 = _RANDOM[11'hF][22];	// rob.scala:260:29, :307:32
        rob_val_21 = _RANDOM[11'hF][23];	// rob.scala:260:29, :307:32
        rob_val_22 = _RANDOM[11'hF][24];	// rob.scala:260:29, :307:32
        rob_val_23 = _RANDOM[11'hF][25];	// rob.scala:260:29, :307:32
        rob_val_24 = _RANDOM[11'hF][26];	// rob.scala:260:29, :307:32
        rob_val_25 = _RANDOM[11'hF][27];	// rob.scala:260:29, :307:32
        rob_val_26 = _RANDOM[11'hF][28];	// rob.scala:260:29, :307:32
        rob_val_27 = _RANDOM[11'hF][29];	// rob.scala:260:29, :307:32
        rob_val_28 = _RANDOM[11'hF][30];	// rob.scala:260:29, :307:32
        rob_val_29 = _RANDOM[11'hF][31];	// rob.scala:260:29, :307:32
        rob_val_30 = _RANDOM[11'h10][0];	// rob.scala:307:32
        rob_val_31 = _RANDOM[11'h10][1];	// rob.scala:307:32
        rob_bsy_0 = _RANDOM[11'h10][2];	// rob.scala:307:32, :308:28
        rob_bsy_1 = _RANDOM[11'h10][3];	// rob.scala:307:32, :308:28
        rob_bsy_2 = _RANDOM[11'h10][4];	// rob.scala:307:32, :308:28
        rob_bsy_3 = _RANDOM[11'h10][5];	// rob.scala:307:32, :308:28
        rob_bsy_4 = _RANDOM[11'h10][6];	// rob.scala:307:32, :308:28
        rob_bsy_5 = _RANDOM[11'h10][7];	// rob.scala:307:32, :308:28
        rob_bsy_6 = _RANDOM[11'h10][8];	// rob.scala:307:32, :308:28
        rob_bsy_7 = _RANDOM[11'h10][9];	// rob.scala:307:32, :308:28
        rob_bsy_8 = _RANDOM[11'h10][10];	// rob.scala:307:32, :308:28
        rob_bsy_9 = _RANDOM[11'h10][11];	// rob.scala:307:32, :308:28
        rob_bsy_10 = _RANDOM[11'h10][12];	// rob.scala:307:32, :308:28
        rob_bsy_11 = _RANDOM[11'h10][13];	// rob.scala:307:32, :308:28
        rob_bsy_12 = _RANDOM[11'h10][14];	// rob.scala:307:32, :308:28
        rob_bsy_13 = _RANDOM[11'h10][15];	// rob.scala:307:32, :308:28
        rob_bsy_14 = _RANDOM[11'h10][16];	// rob.scala:307:32, :308:28
        rob_bsy_15 = _RANDOM[11'h10][17];	// rob.scala:307:32, :308:28
        rob_bsy_16 = _RANDOM[11'h10][18];	// rob.scala:307:32, :308:28
        rob_bsy_17 = _RANDOM[11'h10][19];	// rob.scala:307:32, :308:28
        rob_bsy_18 = _RANDOM[11'h10][20];	// rob.scala:307:32, :308:28
        rob_bsy_19 = _RANDOM[11'h10][21];	// rob.scala:307:32, :308:28
        rob_bsy_20 = _RANDOM[11'h10][22];	// rob.scala:307:32, :308:28
        rob_bsy_21 = _RANDOM[11'h10][23];	// rob.scala:307:32, :308:28
        rob_bsy_22 = _RANDOM[11'h10][24];	// rob.scala:307:32, :308:28
        rob_bsy_23 = _RANDOM[11'h10][25];	// rob.scala:307:32, :308:28
        rob_bsy_24 = _RANDOM[11'h10][26];	// rob.scala:307:32, :308:28
        rob_bsy_25 = _RANDOM[11'h10][27];	// rob.scala:307:32, :308:28
        rob_bsy_26 = _RANDOM[11'h10][28];	// rob.scala:307:32, :308:28
        rob_bsy_27 = _RANDOM[11'h10][29];	// rob.scala:307:32, :308:28
        rob_bsy_28 = _RANDOM[11'h10][30];	// rob.scala:307:32, :308:28
        rob_bsy_29 = _RANDOM[11'h10][31];	// rob.scala:307:32, :308:28
        rob_bsy_30 = _RANDOM[11'h11][0];	// rob.scala:308:28
        rob_bsy_31 = _RANDOM[11'h11][1];	// rob.scala:308:28
        rob_unsafe_0 = _RANDOM[11'h11][2];	// rob.scala:308:28, :309:28
        rob_unsafe_1 = _RANDOM[11'h11][3];	// rob.scala:308:28, :309:28
        rob_unsafe_2 = _RANDOM[11'h11][4];	// rob.scala:308:28, :309:28
        rob_unsafe_3 = _RANDOM[11'h11][5];	// rob.scala:308:28, :309:28
        rob_unsafe_4 = _RANDOM[11'h11][6];	// rob.scala:308:28, :309:28
        rob_unsafe_5 = _RANDOM[11'h11][7];	// rob.scala:308:28, :309:28
        rob_unsafe_6 = _RANDOM[11'h11][8];	// rob.scala:308:28, :309:28
        rob_unsafe_7 = _RANDOM[11'h11][9];	// rob.scala:308:28, :309:28
        rob_unsafe_8 = _RANDOM[11'h11][10];	// rob.scala:308:28, :309:28
        rob_unsafe_9 = _RANDOM[11'h11][11];	// rob.scala:308:28, :309:28
        rob_unsafe_10 = _RANDOM[11'h11][12];	// rob.scala:308:28, :309:28
        rob_unsafe_11 = _RANDOM[11'h11][13];	// rob.scala:308:28, :309:28
        rob_unsafe_12 = _RANDOM[11'h11][14];	// rob.scala:308:28, :309:28
        rob_unsafe_13 = _RANDOM[11'h11][15];	// rob.scala:308:28, :309:28
        rob_unsafe_14 = _RANDOM[11'h11][16];	// rob.scala:308:28, :309:28
        rob_unsafe_15 = _RANDOM[11'h11][17];	// rob.scala:308:28, :309:28
        rob_unsafe_16 = _RANDOM[11'h11][18];	// rob.scala:308:28, :309:28
        rob_unsafe_17 = _RANDOM[11'h11][19];	// rob.scala:308:28, :309:28
        rob_unsafe_18 = _RANDOM[11'h11][20];	// rob.scala:308:28, :309:28
        rob_unsafe_19 = _RANDOM[11'h11][21];	// rob.scala:308:28, :309:28
        rob_unsafe_20 = _RANDOM[11'h11][22];	// rob.scala:308:28, :309:28
        rob_unsafe_21 = _RANDOM[11'h11][23];	// rob.scala:308:28, :309:28
        rob_unsafe_22 = _RANDOM[11'h11][24];	// rob.scala:308:28, :309:28
        rob_unsafe_23 = _RANDOM[11'h11][25];	// rob.scala:308:28, :309:28
        rob_unsafe_24 = _RANDOM[11'h11][26];	// rob.scala:308:28, :309:28
        rob_unsafe_25 = _RANDOM[11'h11][27];	// rob.scala:308:28, :309:28
        rob_unsafe_26 = _RANDOM[11'h11][28];	// rob.scala:308:28, :309:28
        rob_unsafe_27 = _RANDOM[11'h11][29];	// rob.scala:308:28, :309:28
        rob_unsafe_28 = _RANDOM[11'h11][30];	// rob.scala:308:28, :309:28
        rob_unsafe_29 = _RANDOM[11'h11][31];	// rob.scala:308:28, :309:28
        rob_unsafe_30 = _RANDOM[11'h12][0];	// rob.scala:309:28
        rob_unsafe_31 = _RANDOM[11'h12][1];	// rob.scala:309:28
        rob_uop_0_uopc = _RANDOM[11'h12][8:2];	// rob.scala:309:28, :310:28
        rob_uop_0_is_rvc = _RANDOM[11'h14][9];	// rob.scala:310:28
        rob_uop_0_br_mask = {_RANDOM[11'h16][31:30], _RANDOM[11'h17][17:0]};	// rob.scala:310:28
        rob_uop_0_ftq_idx = _RANDOM[11'h17][28:23];	// rob.scala:310:28
        rob_uop_0_edge_inst = _RANDOM[11'h17][29];	// rob.scala:310:28
        rob_uop_0_pc_lob = {_RANDOM[11'h17][31:30], _RANDOM[11'h18][3:0]};	// rob.scala:310:28
        rob_uop_0_pdst = _RANDOM[11'h19][30:24];	// rob.scala:310:28
        rob_uop_0_stale_pdst = {_RANDOM[11'h1A][31:30], _RANDOM[11'h1B][4:0]};	// rob.scala:310:28
        rob_uop_0_is_fencei = _RANDOM[11'h1D][16];	// rob.scala:310:28
        rob_uop_0_uses_ldq = _RANDOM[11'h1D][18];	// rob.scala:310:28
        rob_uop_0_uses_stq = _RANDOM[11'h1D][19];	// rob.scala:310:28
        rob_uop_0_is_sys_pc2epc = _RANDOM[11'h1D][20];	// rob.scala:310:28
        rob_uop_0_flush_on_commit = _RANDOM[11'h1D][22];	// rob.scala:310:28
        rob_uop_0_ldst = _RANDOM[11'h1D][29:24];	// rob.scala:310:28
        rob_uop_0_ldst_val = _RANDOM[11'h1E][16];	// rob.scala:310:28
        rob_uop_0_dst_rtype = _RANDOM[11'h1E][18:17];	// rob.scala:310:28
        rob_uop_0_fp_val = _RANDOM[11'h1E][24];	// rob.scala:310:28
        rob_uop_1_uopc = _RANDOM[11'h1F][9:3];	// rob.scala:310:28
        rob_uop_1_is_rvc = _RANDOM[11'h21][10];	// rob.scala:310:28
        rob_uop_1_br_mask = {_RANDOM[11'h23][31], _RANDOM[11'h24][18:0]};	// rob.scala:310:28
        rob_uop_1_ftq_idx = _RANDOM[11'h24][29:24];	// rob.scala:310:28
        rob_uop_1_edge_inst = _RANDOM[11'h24][30];	// rob.scala:310:28
        rob_uop_1_pc_lob = {_RANDOM[11'h24][31], _RANDOM[11'h25][4:0]};	// rob.scala:310:28
        rob_uop_1_pdst = _RANDOM[11'h26][31:25];	// rob.scala:310:28
        rob_uop_1_stale_pdst = {_RANDOM[11'h27][31], _RANDOM[11'h28][5:0]};	// rob.scala:310:28
        rob_uop_1_is_fencei = _RANDOM[11'h2A][17];	// rob.scala:310:28
        rob_uop_1_uses_ldq = _RANDOM[11'h2A][19];	// rob.scala:310:28
        rob_uop_1_uses_stq = _RANDOM[11'h2A][20];	// rob.scala:310:28
        rob_uop_1_is_sys_pc2epc = _RANDOM[11'h2A][21];	// rob.scala:310:28
        rob_uop_1_flush_on_commit = _RANDOM[11'h2A][23];	// rob.scala:310:28
        rob_uop_1_ldst = _RANDOM[11'h2A][30:25];	// rob.scala:310:28
        rob_uop_1_ldst_val = _RANDOM[11'h2B][17];	// rob.scala:310:28
        rob_uop_1_dst_rtype = _RANDOM[11'h2B][19:18];	// rob.scala:310:28
        rob_uop_1_fp_val = _RANDOM[11'h2B][25];	// rob.scala:310:28
        rob_uop_2_uopc = _RANDOM[11'h2C][10:4];	// rob.scala:310:28
        rob_uop_2_is_rvc = _RANDOM[11'h2E][11];	// rob.scala:310:28
        rob_uop_2_br_mask = _RANDOM[11'h31][19:0];	// rob.scala:310:28
        rob_uop_2_ftq_idx = _RANDOM[11'h31][30:25];	// rob.scala:310:28
        rob_uop_2_edge_inst = _RANDOM[11'h31][31];	// rob.scala:310:28
        rob_uop_2_pc_lob = _RANDOM[11'h32][5:0];	// rob.scala:310:28
        rob_uop_2_pdst = {_RANDOM[11'h33][31:26], _RANDOM[11'h34][0]};	// rob.scala:310:28
        rob_uop_2_stale_pdst = _RANDOM[11'h35][6:0];	// rob.scala:310:28
        rob_uop_2_is_fencei = _RANDOM[11'h37][18];	// rob.scala:310:28
        rob_uop_2_uses_ldq = _RANDOM[11'h37][20];	// rob.scala:310:28
        rob_uop_2_uses_stq = _RANDOM[11'h37][21];	// rob.scala:310:28
        rob_uop_2_is_sys_pc2epc = _RANDOM[11'h37][22];	// rob.scala:310:28
        rob_uop_2_flush_on_commit = _RANDOM[11'h37][24];	// rob.scala:310:28
        rob_uop_2_ldst = _RANDOM[11'h37][31:26];	// rob.scala:310:28
        rob_uop_2_ldst_val = _RANDOM[11'h38][18];	// rob.scala:310:28
        rob_uop_2_dst_rtype = _RANDOM[11'h38][20:19];	// rob.scala:310:28
        rob_uop_2_fp_val = _RANDOM[11'h38][26];	// rob.scala:310:28
        rob_uop_3_uopc = _RANDOM[11'h39][11:5];	// rob.scala:310:28
        rob_uop_3_is_rvc = _RANDOM[11'h3B][12];	// rob.scala:310:28
        rob_uop_3_br_mask = _RANDOM[11'h3E][20:1];	// rob.scala:310:28
        rob_uop_3_ftq_idx = _RANDOM[11'h3E][31:26];	// rob.scala:310:28
        rob_uop_3_edge_inst = _RANDOM[11'h3F][0];	// rob.scala:310:28
        rob_uop_3_pc_lob = _RANDOM[11'h3F][6:1];	// rob.scala:310:28
        rob_uop_3_pdst = {_RANDOM[11'h40][31:27], _RANDOM[11'h41][1:0]};	// rob.scala:310:28
        rob_uop_3_stale_pdst = _RANDOM[11'h42][7:1];	// rob.scala:310:28
        rob_uop_3_is_fencei = _RANDOM[11'h44][19];	// rob.scala:310:28
        rob_uop_3_uses_ldq = _RANDOM[11'h44][21];	// rob.scala:310:28
        rob_uop_3_uses_stq = _RANDOM[11'h44][22];	// rob.scala:310:28
        rob_uop_3_is_sys_pc2epc = _RANDOM[11'h44][23];	// rob.scala:310:28
        rob_uop_3_flush_on_commit = _RANDOM[11'h44][25];	// rob.scala:310:28
        rob_uop_3_ldst = {_RANDOM[11'h44][31:27], _RANDOM[11'h45][0]};	// rob.scala:310:28
        rob_uop_3_ldst_val = _RANDOM[11'h45][19];	// rob.scala:310:28
        rob_uop_3_dst_rtype = _RANDOM[11'h45][21:20];	// rob.scala:310:28
        rob_uop_3_fp_val = _RANDOM[11'h45][27];	// rob.scala:310:28
        rob_uop_4_uopc = _RANDOM[11'h46][12:6];	// rob.scala:310:28
        rob_uop_4_is_rvc = _RANDOM[11'h48][13];	// rob.scala:310:28
        rob_uop_4_br_mask = _RANDOM[11'h4B][21:2];	// rob.scala:310:28
        rob_uop_4_ftq_idx = {_RANDOM[11'h4B][31:27], _RANDOM[11'h4C][0]};	// rob.scala:310:28
        rob_uop_4_edge_inst = _RANDOM[11'h4C][1];	// rob.scala:310:28
        rob_uop_4_pc_lob = _RANDOM[11'h4C][7:2];	// rob.scala:310:28
        rob_uop_4_pdst = {_RANDOM[11'h4D][31:28], _RANDOM[11'h4E][2:0]};	// rob.scala:310:28
        rob_uop_4_stale_pdst = _RANDOM[11'h4F][8:2];	// rob.scala:310:28
        rob_uop_4_is_fencei = _RANDOM[11'h51][20];	// rob.scala:310:28
        rob_uop_4_uses_ldq = _RANDOM[11'h51][22];	// rob.scala:310:28
        rob_uop_4_uses_stq = _RANDOM[11'h51][23];	// rob.scala:310:28
        rob_uop_4_is_sys_pc2epc = _RANDOM[11'h51][24];	// rob.scala:310:28
        rob_uop_4_flush_on_commit = _RANDOM[11'h51][26];	// rob.scala:310:28
        rob_uop_4_ldst = {_RANDOM[11'h51][31:28], _RANDOM[11'h52][1:0]};	// rob.scala:310:28
        rob_uop_4_ldst_val = _RANDOM[11'h52][20];	// rob.scala:310:28
        rob_uop_4_dst_rtype = _RANDOM[11'h52][22:21];	// rob.scala:310:28
        rob_uop_4_fp_val = _RANDOM[11'h52][28];	// rob.scala:310:28
        rob_uop_5_uopc = _RANDOM[11'h53][13:7];	// rob.scala:310:28
        rob_uop_5_is_rvc = _RANDOM[11'h55][14];	// rob.scala:310:28
        rob_uop_5_br_mask = _RANDOM[11'h58][22:3];	// rob.scala:310:28
        rob_uop_5_ftq_idx = {_RANDOM[11'h58][31:28], _RANDOM[11'h59][1:0]};	// rob.scala:310:28
        rob_uop_5_edge_inst = _RANDOM[11'h59][2];	// rob.scala:310:28
        rob_uop_5_pc_lob = _RANDOM[11'h59][8:3];	// rob.scala:310:28
        rob_uop_5_pdst = {_RANDOM[11'h5A][31:29], _RANDOM[11'h5B][3:0]};	// rob.scala:310:28
        rob_uop_5_stale_pdst = _RANDOM[11'h5C][9:3];	// rob.scala:310:28
        rob_uop_5_is_fencei = _RANDOM[11'h5E][21];	// rob.scala:310:28
        rob_uop_5_uses_ldq = _RANDOM[11'h5E][23];	// rob.scala:310:28
        rob_uop_5_uses_stq = _RANDOM[11'h5E][24];	// rob.scala:310:28
        rob_uop_5_is_sys_pc2epc = _RANDOM[11'h5E][25];	// rob.scala:310:28
        rob_uop_5_flush_on_commit = _RANDOM[11'h5E][27];	// rob.scala:310:28
        rob_uop_5_ldst = {_RANDOM[11'h5E][31:29], _RANDOM[11'h5F][2:0]};	// rob.scala:310:28
        rob_uop_5_ldst_val = _RANDOM[11'h5F][21];	// rob.scala:310:28
        rob_uop_5_dst_rtype = _RANDOM[11'h5F][23:22];	// rob.scala:310:28
        rob_uop_5_fp_val = _RANDOM[11'h5F][29];	// rob.scala:310:28
        rob_uop_6_uopc = _RANDOM[11'h60][14:8];	// rob.scala:310:28
        rob_uop_6_is_rvc = _RANDOM[11'h62][15];	// rob.scala:310:28
        rob_uop_6_br_mask = _RANDOM[11'h65][23:4];	// rob.scala:310:28
        rob_uop_6_ftq_idx = {_RANDOM[11'h65][31:29], _RANDOM[11'h66][2:0]};	// rob.scala:310:28
        rob_uop_6_edge_inst = _RANDOM[11'h66][3];	// rob.scala:310:28
        rob_uop_6_pc_lob = _RANDOM[11'h66][9:4];	// rob.scala:310:28
        rob_uop_6_pdst = {_RANDOM[11'h67][31:30], _RANDOM[11'h68][4:0]};	// rob.scala:310:28
        rob_uop_6_stale_pdst = _RANDOM[11'h69][10:4];	// rob.scala:310:28
        rob_uop_6_is_fencei = _RANDOM[11'h6B][22];	// rob.scala:310:28
        rob_uop_6_uses_ldq = _RANDOM[11'h6B][24];	// rob.scala:310:28
        rob_uop_6_uses_stq = _RANDOM[11'h6B][25];	// rob.scala:310:28
        rob_uop_6_is_sys_pc2epc = _RANDOM[11'h6B][26];	// rob.scala:310:28
        rob_uop_6_flush_on_commit = _RANDOM[11'h6B][28];	// rob.scala:310:28
        rob_uop_6_ldst = {_RANDOM[11'h6B][31:30], _RANDOM[11'h6C][3:0]};	// rob.scala:310:28
        rob_uop_6_ldst_val = _RANDOM[11'h6C][22];	// rob.scala:310:28
        rob_uop_6_dst_rtype = _RANDOM[11'h6C][24:23];	// rob.scala:310:28
        rob_uop_6_fp_val = _RANDOM[11'h6C][30];	// rob.scala:310:28
        rob_uop_7_uopc = _RANDOM[11'h6D][15:9];	// rob.scala:310:28
        rob_uop_7_is_rvc = _RANDOM[11'h6F][16];	// rob.scala:310:28
        rob_uop_7_br_mask = _RANDOM[11'h72][24:5];	// rob.scala:310:28
        rob_uop_7_ftq_idx = {_RANDOM[11'h72][31:30], _RANDOM[11'h73][3:0]};	// rob.scala:310:28
        rob_uop_7_edge_inst = _RANDOM[11'h73][4];	// rob.scala:310:28
        rob_uop_7_pc_lob = _RANDOM[11'h73][10:5];	// rob.scala:310:28
        rob_uop_7_pdst = {_RANDOM[11'h74][31], _RANDOM[11'h75][5:0]};	// rob.scala:310:28
        rob_uop_7_stale_pdst = _RANDOM[11'h76][11:5];	// rob.scala:310:28
        rob_uop_7_is_fencei = _RANDOM[11'h78][23];	// rob.scala:310:28
        rob_uop_7_uses_ldq = _RANDOM[11'h78][25];	// rob.scala:310:28
        rob_uop_7_uses_stq = _RANDOM[11'h78][26];	// rob.scala:310:28
        rob_uop_7_is_sys_pc2epc = _RANDOM[11'h78][27];	// rob.scala:310:28
        rob_uop_7_flush_on_commit = _RANDOM[11'h78][29];	// rob.scala:310:28
        rob_uop_7_ldst = {_RANDOM[11'h78][31], _RANDOM[11'h79][4:0]};	// rob.scala:310:28
        rob_uop_7_ldst_val = _RANDOM[11'h79][23];	// rob.scala:310:28
        rob_uop_7_dst_rtype = _RANDOM[11'h79][25:24];	// rob.scala:310:28
        rob_uop_7_fp_val = _RANDOM[11'h79][31];	// rob.scala:310:28
        rob_uop_8_uopc = _RANDOM[11'h7A][16:10];	// rob.scala:310:28
        rob_uop_8_is_rvc = _RANDOM[11'h7C][17];	// rob.scala:310:28
        rob_uop_8_br_mask = _RANDOM[11'h7F][25:6];	// rob.scala:310:28
        rob_uop_8_ftq_idx = {_RANDOM[11'h7F][31], _RANDOM[11'h80][4:0]};	// rob.scala:310:28
        rob_uop_8_edge_inst = _RANDOM[11'h80][5];	// rob.scala:310:28
        rob_uop_8_pc_lob = _RANDOM[11'h80][11:6];	// rob.scala:310:28
        rob_uop_8_pdst = _RANDOM[11'h82][6:0];	// rob.scala:310:28
        rob_uop_8_stale_pdst = _RANDOM[11'h83][12:6];	// rob.scala:310:28
        rob_uop_8_is_fencei = _RANDOM[11'h85][24];	// rob.scala:310:28
        rob_uop_8_uses_ldq = _RANDOM[11'h85][26];	// rob.scala:310:28
        rob_uop_8_uses_stq = _RANDOM[11'h85][27];	// rob.scala:310:28
        rob_uop_8_is_sys_pc2epc = _RANDOM[11'h85][28];	// rob.scala:310:28
        rob_uop_8_flush_on_commit = _RANDOM[11'h85][30];	// rob.scala:310:28
        rob_uop_8_ldst = _RANDOM[11'h86][5:0];	// rob.scala:310:28
        rob_uop_8_ldst_val = _RANDOM[11'h86][24];	// rob.scala:310:28
        rob_uop_8_dst_rtype = _RANDOM[11'h86][26:25];	// rob.scala:310:28
        rob_uop_8_fp_val = _RANDOM[11'h87][0];	// rob.scala:310:28
        rob_uop_9_uopc = _RANDOM[11'h87][17:11];	// rob.scala:310:28
        rob_uop_9_is_rvc = _RANDOM[11'h89][18];	// rob.scala:310:28
        rob_uop_9_br_mask = _RANDOM[11'h8C][26:7];	// rob.scala:310:28
        rob_uop_9_ftq_idx = _RANDOM[11'h8D][5:0];	// rob.scala:310:28
        rob_uop_9_edge_inst = _RANDOM[11'h8D][6];	// rob.scala:310:28
        rob_uop_9_pc_lob = _RANDOM[11'h8D][12:7];	// rob.scala:310:28
        rob_uop_9_pdst = _RANDOM[11'h8F][7:1];	// rob.scala:310:28
        rob_uop_9_stale_pdst = _RANDOM[11'h90][13:7];	// rob.scala:310:28
        rob_uop_9_is_fencei = _RANDOM[11'h92][25];	// rob.scala:310:28
        rob_uop_9_uses_ldq = _RANDOM[11'h92][27];	// rob.scala:310:28
        rob_uop_9_uses_stq = _RANDOM[11'h92][28];	// rob.scala:310:28
        rob_uop_9_is_sys_pc2epc = _RANDOM[11'h92][29];	// rob.scala:310:28
        rob_uop_9_flush_on_commit = _RANDOM[11'h92][31];	// rob.scala:310:28
        rob_uop_9_ldst = _RANDOM[11'h93][6:1];	// rob.scala:310:28
        rob_uop_9_ldst_val = _RANDOM[11'h93][25];	// rob.scala:310:28
        rob_uop_9_dst_rtype = _RANDOM[11'h93][27:26];	// rob.scala:310:28
        rob_uop_9_fp_val = _RANDOM[11'h94][1];	// rob.scala:310:28
        rob_uop_10_uopc = _RANDOM[11'h94][18:12];	// rob.scala:310:28
        rob_uop_10_is_rvc = _RANDOM[11'h96][19];	// rob.scala:310:28
        rob_uop_10_br_mask = _RANDOM[11'h99][27:8];	// rob.scala:310:28
        rob_uop_10_ftq_idx = _RANDOM[11'h9A][6:1];	// rob.scala:310:28
        rob_uop_10_edge_inst = _RANDOM[11'h9A][7];	// rob.scala:310:28
        rob_uop_10_pc_lob = _RANDOM[11'h9A][13:8];	// rob.scala:310:28
        rob_uop_10_pdst = _RANDOM[11'h9C][8:2];	// rob.scala:310:28
        rob_uop_10_stale_pdst = _RANDOM[11'h9D][14:8];	// rob.scala:310:28
        rob_uop_10_is_fencei = _RANDOM[11'h9F][26];	// rob.scala:310:28
        rob_uop_10_uses_ldq = _RANDOM[11'h9F][28];	// rob.scala:310:28
        rob_uop_10_uses_stq = _RANDOM[11'h9F][29];	// rob.scala:310:28
        rob_uop_10_is_sys_pc2epc = _RANDOM[11'h9F][30];	// rob.scala:310:28
        rob_uop_10_flush_on_commit = _RANDOM[11'hA0][0];	// rob.scala:310:28
        rob_uop_10_ldst = _RANDOM[11'hA0][7:2];	// rob.scala:310:28
        rob_uop_10_ldst_val = _RANDOM[11'hA0][26];	// rob.scala:310:28
        rob_uop_10_dst_rtype = _RANDOM[11'hA0][28:27];	// rob.scala:310:28
        rob_uop_10_fp_val = _RANDOM[11'hA1][2];	// rob.scala:310:28
        rob_uop_11_uopc = _RANDOM[11'hA1][19:13];	// rob.scala:310:28
        rob_uop_11_is_rvc = _RANDOM[11'hA3][20];	// rob.scala:310:28
        rob_uop_11_br_mask = _RANDOM[11'hA6][28:9];	// rob.scala:310:28
        rob_uop_11_ftq_idx = _RANDOM[11'hA7][7:2];	// rob.scala:310:28
        rob_uop_11_edge_inst = _RANDOM[11'hA7][8];	// rob.scala:310:28
        rob_uop_11_pc_lob = _RANDOM[11'hA7][14:9];	// rob.scala:310:28
        rob_uop_11_pdst = _RANDOM[11'hA9][9:3];	// rob.scala:310:28
        rob_uop_11_stale_pdst = _RANDOM[11'hAA][15:9];	// rob.scala:310:28
        rob_uop_11_is_fencei = _RANDOM[11'hAC][27];	// rob.scala:310:28
        rob_uop_11_uses_ldq = _RANDOM[11'hAC][29];	// rob.scala:310:28
        rob_uop_11_uses_stq = _RANDOM[11'hAC][30];	// rob.scala:310:28
        rob_uop_11_is_sys_pc2epc = _RANDOM[11'hAC][31];	// rob.scala:310:28
        rob_uop_11_flush_on_commit = _RANDOM[11'hAD][1];	// rob.scala:310:28
        rob_uop_11_ldst = _RANDOM[11'hAD][8:3];	// rob.scala:310:28
        rob_uop_11_ldst_val = _RANDOM[11'hAD][27];	// rob.scala:310:28
        rob_uop_11_dst_rtype = _RANDOM[11'hAD][29:28];	// rob.scala:310:28
        rob_uop_11_fp_val = _RANDOM[11'hAE][3];	// rob.scala:310:28
        rob_uop_12_uopc = _RANDOM[11'hAE][20:14];	// rob.scala:310:28
        rob_uop_12_is_rvc = _RANDOM[11'hB0][21];	// rob.scala:310:28
        rob_uop_12_br_mask = _RANDOM[11'hB3][29:10];	// rob.scala:310:28
        rob_uop_12_ftq_idx = _RANDOM[11'hB4][8:3];	// rob.scala:310:28
        rob_uop_12_edge_inst = _RANDOM[11'hB4][9];	// rob.scala:310:28
        rob_uop_12_pc_lob = _RANDOM[11'hB4][15:10];	// rob.scala:310:28
        rob_uop_12_pdst = _RANDOM[11'hB6][10:4];	// rob.scala:310:28
        rob_uop_12_stale_pdst = _RANDOM[11'hB7][16:10];	// rob.scala:310:28
        rob_uop_12_is_fencei = _RANDOM[11'hB9][28];	// rob.scala:310:28
        rob_uop_12_uses_ldq = _RANDOM[11'hB9][30];	// rob.scala:310:28
        rob_uop_12_uses_stq = _RANDOM[11'hB9][31];	// rob.scala:310:28
        rob_uop_12_is_sys_pc2epc = _RANDOM[11'hBA][0];	// rob.scala:310:28
        rob_uop_12_flush_on_commit = _RANDOM[11'hBA][2];	// rob.scala:310:28
        rob_uop_12_ldst = _RANDOM[11'hBA][9:4];	// rob.scala:310:28
        rob_uop_12_ldst_val = _RANDOM[11'hBA][28];	// rob.scala:310:28
        rob_uop_12_dst_rtype = _RANDOM[11'hBA][30:29];	// rob.scala:310:28
        rob_uop_12_fp_val = _RANDOM[11'hBB][4];	// rob.scala:310:28
        rob_uop_13_uopc = _RANDOM[11'hBB][21:15];	// rob.scala:310:28
        rob_uop_13_is_rvc = _RANDOM[11'hBD][22];	// rob.scala:310:28
        rob_uop_13_br_mask = _RANDOM[11'hC0][30:11];	// rob.scala:310:28
        rob_uop_13_ftq_idx = _RANDOM[11'hC1][9:4];	// rob.scala:310:28
        rob_uop_13_edge_inst = _RANDOM[11'hC1][10];	// rob.scala:310:28
        rob_uop_13_pc_lob = _RANDOM[11'hC1][16:11];	// rob.scala:310:28
        rob_uop_13_pdst = _RANDOM[11'hC3][11:5];	// rob.scala:310:28
        rob_uop_13_stale_pdst = _RANDOM[11'hC4][17:11];	// rob.scala:310:28
        rob_uop_13_is_fencei = _RANDOM[11'hC6][29];	// rob.scala:310:28
        rob_uop_13_uses_ldq = _RANDOM[11'hC6][31];	// rob.scala:310:28
        rob_uop_13_uses_stq = _RANDOM[11'hC7][0];	// rob.scala:310:28
        rob_uop_13_is_sys_pc2epc = _RANDOM[11'hC7][1];	// rob.scala:310:28
        rob_uop_13_flush_on_commit = _RANDOM[11'hC7][3];	// rob.scala:310:28
        rob_uop_13_ldst = _RANDOM[11'hC7][10:5];	// rob.scala:310:28
        rob_uop_13_ldst_val = _RANDOM[11'hC7][29];	// rob.scala:310:28
        rob_uop_13_dst_rtype = _RANDOM[11'hC7][31:30];	// rob.scala:310:28
        rob_uop_13_fp_val = _RANDOM[11'hC8][5];	// rob.scala:310:28
        rob_uop_14_uopc = _RANDOM[11'hC8][22:16];	// rob.scala:310:28
        rob_uop_14_is_rvc = _RANDOM[11'hCA][23];	// rob.scala:310:28
        rob_uop_14_br_mask = _RANDOM[11'hCD][31:12];	// rob.scala:310:28
        rob_uop_14_ftq_idx = _RANDOM[11'hCE][10:5];	// rob.scala:310:28
        rob_uop_14_edge_inst = _RANDOM[11'hCE][11];	// rob.scala:310:28
        rob_uop_14_pc_lob = _RANDOM[11'hCE][17:12];	// rob.scala:310:28
        rob_uop_14_pdst = _RANDOM[11'hD0][12:6];	// rob.scala:310:28
        rob_uop_14_stale_pdst = _RANDOM[11'hD1][18:12];	// rob.scala:310:28
        rob_uop_14_is_fencei = _RANDOM[11'hD3][30];	// rob.scala:310:28
        rob_uop_14_uses_ldq = _RANDOM[11'hD4][0];	// rob.scala:310:28
        rob_uop_14_uses_stq = _RANDOM[11'hD4][1];	// rob.scala:310:28
        rob_uop_14_is_sys_pc2epc = _RANDOM[11'hD4][2];	// rob.scala:310:28
        rob_uop_14_flush_on_commit = _RANDOM[11'hD4][4];	// rob.scala:310:28
        rob_uop_14_ldst = _RANDOM[11'hD4][11:6];	// rob.scala:310:28
        rob_uop_14_ldst_val = _RANDOM[11'hD4][30];	// rob.scala:310:28
        rob_uop_14_dst_rtype = {_RANDOM[11'hD4][31], _RANDOM[11'hD5][0]};	// rob.scala:310:28
        rob_uop_14_fp_val = _RANDOM[11'hD5][6];	// rob.scala:310:28
        rob_uop_15_uopc = _RANDOM[11'hD5][23:17];	// rob.scala:310:28
        rob_uop_15_is_rvc = _RANDOM[11'hD7][24];	// rob.scala:310:28
        rob_uop_15_br_mask = {_RANDOM[11'hDA][31:13], _RANDOM[11'hDB][0]};	// rob.scala:310:28
        rob_uop_15_ftq_idx = _RANDOM[11'hDB][11:6];	// rob.scala:310:28
        rob_uop_15_edge_inst = _RANDOM[11'hDB][12];	// rob.scala:310:28
        rob_uop_15_pc_lob = _RANDOM[11'hDB][18:13];	// rob.scala:310:28
        rob_uop_15_pdst = _RANDOM[11'hDD][13:7];	// rob.scala:310:28
        rob_uop_15_stale_pdst = _RANDOM[11'hDE][19:13];	// rob.scala:310:28
        rob_uop_15_is_fencei = _RANDOM[11'hE0][31];	// rob.scala:310:28
        rob_uop_15_uses_ldq = _RANDOM[11'hE1][1];	// rob.scala:310:28
        rob_uop_15_uses_stq = _RANDOM[11'hE1][2];	// rob.scala:310:28
        rob_uop_15_is_sys_pc2epc = _RANDOM[11'hE1][3];	// rob.scala:310:28
        rob_uop_15_flush_on_commit = _RANDOM[11'hE1][5];	// rob.scala:310:28
        rob_uop_15_ldst = _RANDOM[11'hE1][12:7];	// rob.scala:310:28
        rob_uop_15_ldst_val = _RANDOM[11'hE1][31];	// rob.scala:310:28
        rob_uop_15_dst_rtype = _RANDOM[11'hE2][1:0];	// rob.scala:310:28
        rob_uop_15_fp_val = _RANDOM[11'hE2][7];	// rob.scala:310:28
        rob_uop_16_uopc = _RANDOM[11'hE2][24:18];	// rob.scala:310:28
        rob_uop_16_is_rvc = _RANDOM[11'hE4][25];	// rob.scala:310:28
        rob_uop_16_br_mask = {_RANDOM[11'hE7][31:14], _RANDOM[11'hE8][1:0]};	// rob.scala:310:28
        rob_uop_16_ftq_idx = _RANDOM[11'hE8][12:7];	// rob.scala:310:28
        rob_uop_16_edge_inst = _RANDOM[11'hE8][13];	// rob.scala:310:28
        rob_uop_16_pc_lob = _RANDOM[11'hE8][19:14];	// rob.scala:310:28
        rob_uop_16_pdst = _RANDOM[11'hEA][14:8];	// rob.scala:310:28
        rob_uop_16_stale_pdst = _RANDOM[11'hEB][20:14];	// rob.scala:310:28
        rob_uop_16_is_fencei = _RANDOM[11'hEE][0];	// rob.scala:310:28
        rob_uop_16_uses_ldq = _RANDOM[11'hEE][2];	// rob.scala:310:28
        rob_uop_16_uses_stq = _RANDOM[11'hEE][3];	// rob.scala:310:28
        rob_uop_16_is_sys_pc2epc = _RANDOM[11'hEE][4];	// rob.scala:310:28
        rob_uop_16_flush_on_commit = _RANDOM[11'hEE][6];	// rob.scala:310:28
        rob_uop_16_ldst = _RANDOM[11'hEE][13:8];	// rob.scala:310:28
        rob_uop_16_ldst_val = _RANDOM[11'hEF][0];	// rob.scala:310:28
        rob_uop_16_dst_rtype = _RANDOM[11'hEF][2:1];	// rob.scala:310:28
        rob_uop_16_fp_val = _RANDOM[11'hEF][8];	// rob.scala:310:28
        rob_uop_17_uopc = _RANDOM[11'hEF][25:19];	// rob.scala:310:28
        rob_uop_17_is_rvc = _RANDOM[11'hF1][26];	// rob.scala:310:28
        rob_uop_17_br_mask = {_RANDOM[11'hF4][31:15], _RANDOM[11'hF5][2:0]};	// rob.scala:310:28
        rob_uop_17_ftq_idx = _RANDOM[11'hF5][13:8];	// rob.scala:310:28
        rob_uop_17_edge_inst = _RANDOM[11'hF5][14];	// rob.scala:310:28
        rob_uop_17_pc_lob = _RANDOM[11'hF5][20:15];	// rob.scala:310:28
        rob_uop_17_pdst = _RANDOM[11'hF7][15:9];	// rob.scala:310:28
        rob_uop_17_stale_pdst = _RANDOM[11'hF8][21:15];	// rob.scala:310:28
        rob_uop_17_is_fencei = _RANDOM[11'hFB][1];	// rob.scala:310:28
        rob_uop_17_uses_ldq = _RANDOM[11'hFB][3];	// rob.scala:310:28
        rob_uop_17_uses_stq = _RANDOM[11'hFB][4];	// rob.scala:310:28
        rob_uop_17_is_sys_pc2epc = _RANDOM[11'hFB][5];	// rob.scala:310:28
        rob_uop_17_flush_on_commit = _RANDOM[11'hFB][7];	// rob.scala:310:28
        rob_uop_17_ldst = _RANDOM[11'hFB][14:9];	// rob.scala:310:28
        rob_uop_17_ldst_val = _RANDOM[11'hFC][1];	// rob.scala:310:28
        rob_uop_17_dst_rtype = _RANDOM[11'hFC][3:2];	// rob.scala:310:28
        rob_uop_17_fp_val = _RANDOM[11'hFC][9];	// rob.scala:310:28
        rob_uop_18_uopc = _RANDOM[11'hFC][26:20];	// rob.scala:310:28
        rob_uop_18_is_rvc = _RANDOM[11'hFE][27];	// rob.scala:310:28
        rob_uop_18_br_mask = {_RANDOM[11'h101][31:16], _RANDOM[11'h102][3:0]};	// rob.scala:310:28
        rob_uop_18_ftq_idx = _RANDOM[11'h102][14:9];	// rob.scala:310:28
        rob_uop_18_edge_inst = _RANDOM[11'h102][15];	// rob.scala:310:28
        rob_uop_18_pc_lob = _RANDOM[11'h102][21:16];	// rob.scala:310:28
        rob_uop_18_pdst = _RANDOM[11'h104][16:10];	// rob.scala:310:28
        rob_uop_18_stale_pdst = _RANDOM[11'h105][22:16];	// rob.scala:310:28
        rob_uop_18_is_fencei = _RANDOM[11'h108][2];	// rob.scala:310:28
        rob_uop_18_uses_ldq = _RANDOM[11'h108][4];	// rob.scala:310:28
        rob_uop_18_uses_stq = _RANDOM[11'h108][5];	// rob.scala:310:28
        rob_uop_18_is_sys_pc2epc = _RANDOM[11'h108][6];	// rob.scala:310:28
        rob_uop_18_flush_on_commit = _RANDOM[11'h108][8];	// rob.scala:310:28
        rob_uop_18_ldst = _RANDOM[11'h108][15:10];	// rob.scala:310:28
        rob_uop_18_ldst_val = _RANDOM[11'h109][2];	// rob.scala:310:28
        rob_uop_18_dst_rtype = _RANDOM[11'h109][4:3];	// rob.scala:310:28
        rob_uop_18_fp_val = _RANDOM[11'h109][10];	// rob.scala:310:28
        rob_uop_19_uopc = _RANDOM[11'h109][27:21];	// rob.scala:310:28
        rob_uop_19_is_rvc = _RANDOM[11'h10B][28];	// rob.scala:310:28
        rob_uop_19_br_mask = {_RANDOM[11'h10E][31:17], _RANDOM[11'h10F][4:0]};	// rob.scala:310:28
        rob_uop_19_ftq_idx = _RANDOM[11'h10F][15:10];	// rob.scala:310:28
        rob_uop_19_edge_inst = _RANDOM[11'h10F][16];	// rob.scala:310:28
        rob_uop_19_pc_lob = _RANDOM[11'h10F][22:17];	// rob.scala:310:28
        rob_uop_19_pdst = _RANDOM[11'h111][17:11];	// rob.scala:310:28
        rob_uop_19_stale_pdst = _RANDOM[11'h112][23:17];	// rob.scala:310:28
        rob_uop_19_is_fencei = _RANDOM[11'h115][3];	// rob.scala:310:28
        rob_uop_19_uses_ldq = _RANDOM[11'h115][5];	// rob.scala:310:28
        rob_uop_19_uses_stq = _RANDOM[11'h115][6];	// rob.scala:310:28
        rob_uop_19_is_sys_pc2epc = _RANDOM[11'h115][7];	// rob.scala:310:28
        rob_uop_19_flush_on_commit = _RANDOM[11'h115][9];	// rob.scala:310:28
        rob_uop_19_ldst = _RANDOM[11'h115][16:11];	// rob.scala:310:28
        rob_uop_19_ldst_val = _RANDOM[11'h116][3];	// rob.scala:310:28
        rob_uop_19_dst_rtype = _RANDOM[11'h116][5:4];	// rob.scala:310:28
        rob_uop_19_fp_val = _RANDOM[11'h116][11];	// rob.scala:310:28
        rob_uop_20_uopc = _RANDOM[11'h116][28:22];	// rob.scala:310:28
        rob_uop_20_is_rvc = _RANDOM[11'h118][29];	// rob.scala:310:28
        rob_uop_20_br_mask = {_RANDOM[11'h11B][31:18], _RANDOM[11'h11C][5:0]};	// rob.scala:310:28
        rob_uop_20_ftq_idx = _RANDOM[11'h11C][16:11];	// rob.scala:310:28
        rob_uop_20_edge_inst = _RANDOM[11'h11C][17];	// rob.scala:310:28
        rob_uop_20_pc_lob = _RANDOM[11'h11C][23:18];	// rob.scala:310:28
        rob_uop_20_pdst = _RANDOM[11'h11E][18:12];	// rob.scala:310:28
        rob_uop_20_stale_pdst = _RANDOM[11'h11F][24:18];	// rob.scala:310:28
        rob_uop_20_is_fencei = _RANDOM[11'h122][4];	// rob.scala:310:28
        rob_uop_20_uses_ldq = _RANDOM[11'h122][6];	// rob.scala:310:28
        rob_uop_20_uses_stq = _RANDOM[11'h122][7];	// rob.scala:310:28
        rob_uop_20_is_sys_pc2epc = _RANDOM[11'h122][8];	// rob.scala:310:28
        rob_uop_20_flush_on_commit = _RANDOM[11'h122][10];	// rob.scala:310:28
        rob_uop_20_ldst = _RANDOM[11'h122][17:12];	// rob.scala:310:28
        rob_uop_20_ldst_val = _RANDOM[11'h123][4];	// rob.scala:310:28
        rob_uop_20_dst_rtype = _RANDOM[11'h123][6:5];	// rob.scala:310:28
        rob_uop_20_fp_val = _RANDOM[11'h123][12];	// rob.scala:310:28
        rob_uop_21_uopc = _RANDOM[11'h123][29:23];	// rob.scala:310:28
        rob_uop_21_is_rvc = _RANDOM[11'h125][30];	// rob.scala:310:28
        rob_uop_21_br_mask = {_RANDOM[11'h128][31:19], _RANDOM[11'h129][6:0]};	// rob.scala:310:28
        rob_uop_21_ftq_idx = _RANDOM[11'h129][17:12];	// rob.scala:310:28
        rob_uop_21_edge_inst = _RANDOM[11'h129][18];	// rob.scala:310:28
        rob_uop_21_pc_lob = _RANDOM[11'h129][24:19];	// rob.scala:310:28
        rob_uop_21_pdst = _RANDOM[11'h12B][19:13];	// rob.scala:310:28
        rob_uop_21_stale_pdst = _RANDOM[11'h12C][25:19];	// rob.scala:310:28
        rob_uop_21_is_fencei = _RANDOM[11'h12F][5];	// rob.scala:310:28
        rob_uop_21_uses_ldq = _RANDOM[11'h12F][7];	// rob.scala:310:28
        rob_uop_21_uses_stq = _RANDOM[11'h12F][8];	// rob.scala:310:28
        rob_uop_21_is_sys_pc2epc = _RANDOM[11'h12F][9];	// rob.scala:310:28
        rob_uop_21_flush_on_commit = _RANDOM[11'h12F][11];	// rob.scala:310:28
        rob_uop_21_ldst = _RANDOM[11'h12F][18:13];	// rob.scala:310:28
        rob_uop_21_ldst_val = _RANDOM[11'h130][5];	// rob.scala:310:28
        rob_uop_21_dst_rtype = _RANDOM[11'h130][7:6];	// rob.scala:310:28
        rob_uop_21_fp_val = _RANDOM[11'h130][13];	// rob.scala:310:28
        rob_uop_22_uopc = _RANDOM[11'h130][30:24];	// rob.scala:310:28
        rob_uop_22_is_rvc = _RANDOM[11'h132][31];	// rob.scala:310:28
        rob_uop_22_br_mask = {_RANDOM[11'h135][31:20], _RANDOM[11'h136][7:0]};	// rob.scala:310:28
        rob_uop_22_ftq_idx = _RANDOM[11'h136][18:13];	// rob.scala:310:28
        rob_uop_22_edge_inst = _RANDOM[11'h136][19];	// rob.scala:310:28
        rob_uop_22_pc_lob = _RANDOM[11'h136][25:20];	// rob.scala:310:28
        rob_uop_22_pdst = _RANDOM[11'h138][20:14];	// rob.scala:310:28
        rob_uop_22_stale_pdst = _RANDOM[11'h139][26:20];	// rob.scala:310:28
        rob_uop_22_is_fencei = _RANDOM[11'h13C][6];	// rob.scala:310:28
        rob_uop_22_uses_ldq = _RANDOM[11'h13C][8];	// rob.scala:310:28
        rob_uop_22_uses_stq = _RANDOM[11'h13C][9];	// rob.scala:310:28
        rob_uop_22_is_sys_pc2epc = _RANDOM[11'h13C][10];	// rob.scala:310:28
        rob_uop_22_flush_on_commit = _RANDOM[11'h13C][12];	// rob.scala:310:28
        rob_uop_22_ldst = _RANDOM[11'h13C][19:14];	// rob.scala:310:28
        rob_uop_22_ldst_val = _RANDOM[11'h13D][6];	// rob.scala:310:28
        rob_uop_22_dst_rtype = _RANDOM[11'h13D][8:7];	// rob.scala:310:28
        rob_uop_22_fp_val = _RANDOM[11'h13D][14];	// rob.scala:310:28
        rob_uop_23_uopc = _RANDOM[11'h13D][31:25];	// rob.scala:310:28
        rob_uop_23_is_rvc = _RANDOM[11'h140][0];	// rob.scala:310:28
        rob_uop_23_br_mask = {_RANDOM[11'h142][31:21], _RANDOM[11'h143][8:0]};	// rob.scala:310:28
        rob_uop_23_ftq_idx = _RANDOM[11'h143][19:14];	// rob.scala:310:28
        rob_uop_23_edge_inst = _RANDOM[11'h143][20];	// rob.scala:310:28
        rob_uop_23_pc_lob = _RANDOM[11'h143][26:21];	// rob.scala:310:28
        rob_uop_23_pdst = _RANDOM[11'h145][21:15];	// rob.scala:310:28
        rob_uop_23_stale_pdst = _RANDOM[11'h146][27:21];	// rob.scala:310:28
        rob_uop_23_is_fencei = _RANDOM[11'h149][7];	// rob.scala:310:28
        rob_uop_23_uses_ldq = _RANDOM[11'h149][9];	// rob.scala:310:28
        rob_uop_23_uses_stq = _RANDOM[11'h149][10];	// rob.scala:310:28
        rob_uop_23_is_sys_pc2epc = _RANDOM[11'h149][11];	// rob.scala:310:28
        rob_uop_23_flush_on_commit = _RANDOM[11'h149][13];	// rob.scala:310:28
        rob_uop_23_ldst = _RANDOM[11'h149][20:15];	// rob.scala:310:28
        rob_uop_23_ldst_val = _RANDOM[11'h14A][7];	// rob.scala:310:28
        rob_uop_23_dst_rtype = _RANDOM[11'h14A][9:8];	// rob.scala:310:28
        rob_uop_23_fp_val = _RANDOM[11'h14A][15];	// rob.scala:310:28
        rob_uop_24_uopc = {_RANDOM[11'h14A][31:26], _RANDOM[11'h14B][0]};	// rob.scala:310:28
        rob_uop_24_is_rvc = _RANDOM[11'h14D][1];	// rob.scala:310:28
        rob_uop_24_br_mask = {_RANDOM[11'h14F][31:22], _RANDOM[11'h150][9:0]};	// rob.scala:310:28
        rob_uop_24_ftq_idx = _RANDOM[11'h150][20:15];	// rob.scala:310:28
        rob_uop_24_edge_inst = _RANDOM[11'h150][21];	// rob.scala:310:28
        rob_uop_24_pc_lob = _RANDOM[11'h150][27:22];	// rob.scala:310:28
        rob_uop_24_pdst = _RANDOM[11'h152][22:16];	// rob.scala:310:28
        rob_uop_24_stale_pdst = _RANDOM[11'h153][28:22];	// rob.scala:310:28
        rob_uop_24_is_fencei = _RANDOM[11'h156][8];	// rob.scala:310:28
        rob_uop_24_uses_ldq = _RANDOM[11'h156][10];	// rob.scala:310:28
        rob_uop_24_uses_stq = _RANDOM[11'h156][11];	// rob.scala:310:28
        rob_uop_24_is_sys_pc2epc = _RANDOM[11'h156][12];	// rob.scala:310:28
        rob_uop_24_flush_on_commit = _RANDOM[11'h156][14];	// rob.scala:310:28
        rob_uop_24_ldst = _RANDOM[11'h156][21:16];	// rob.scala:310:28
        rob_uop_24_ldst_val = _RANDOM[11'h157][8];	// rob.scala:310:28
        rob_uop_24_dst_rtype = _RANDOM[11'h157][10:9];	// rob.scala:310:28
        rob_uop_24_fp_val = _RANDOM[11'h157][16];	// rob.scala:310:28
        rob_uop_25_uopc = {_RANDOM[11'h157][31:27], _RANDOM[11'h158][1:0]};	// rob.scala:310:28
        rob_uop_25_is_rvc = _RANDOM[11'h15A][2];	// rob.scala:310:28
        rob_uop_25_br_mask = {_RANDOM[11'h15C][31:23], _RANDOM[11'h15D][10:0]};	// rob.scala:310:28
        rob_uop_25_ftq_idx = _RANDOM[11'h15D][21:16];	// rob.scala:310:28
        rob_uop_25_edge_inst = _RANDOM[11'h15D][22];	// rob.scala:310:28
        rob_uop_25_pc_lob = _RANDOM[11'h15D][28:23];	// rob.scala:310:28
        rob_uop_25_pdst = _RANDOM[11'h15F][23:17];	// rob.scala:310:28
        rob_uop_25_stale_pdst = _RANDOM[11'h160][29:23];	// rob.scala:310:28
        rob_uop_25_is_fencei = _RANDOM[11'h163][9];	// rob.scala:310:28
        rob_uop_25_uses_ldq = _RANDOM[11'h163][11];	// rob.scala:310:28
        rob_uop_25_uses_stq = _RANDOM[11'h163][12];	// rob.scala:310:28
        rob_uop_25_is_sys_pc2epc = _RANDOM[11'h163][13];	// rob.scala:310:28
        rob_uop_25_flush_on_commit = _RANDOM[11'h163][15];	// rob.scala:310:28
        rob_uop_25_ldst = _RANDOM[11'h163][22:17];	// rob.scala:310:28
        rob_uop_25_ldst_val = _RANDOM[11'h164][9];	// rob.scala:310:28
        rob_uop_25_dst_rtype = _RANDOM[11'h164][11:10];	// rob.scala:310:28
        rob_uop_25_fp_val = _RANDOM[11'h164][17];	// rob.scala:310:28
        rob_uop_26_uopc = {_RANDOM[11'h164][31:28], _RANDOM[11'h165][2:0]};	// rob.scala:310:28
        rob_uop_26_is_rvc = _RANDOM[11'h167][3];	// rob.scala:310:28
        rob_uop_26_br_mask = {_RANDOM[11'h169][31:24], _RANDOM[11'h16A][11:0]};	// rob.scala:310:28
        rob_uop_26_ftq_idx = _RANDOM[11'h16A][22:17];	// rob.scala:310:28
        rob_uop_26_edge_inst = _RANDOM[11'h16A][23];	// rob.scala:310:28
        rob_uop_26_pc_lob = _RANDOM[11'h16A][29:24];	// rob.scala:310:28
        rob_uop_26_pdst = _RANDOM[11'h16C][24:18];	// rob.scala:310:28
        rob_uop_26_stale_pdst = _RANDOM[11'h16D][30:24];	// rob.scala:310:28
        rob_uop_26_is_fencei = _RANDOM[11'h170][10];	// rob.scala:310:28
        rob_uop_26_uses_ldq = _RANDOM[11'h170][12];	// rob.scala:310:28
        rob_uop_26_uses_stq = _RANDOM[11'h170][13];	// rob.scala:310:28
        rob_uop_26_is_sys_pc2epc = _RANDOM[11'h170][14];	// rob.scala:310:28
        rob_uop_26_flush_on_commit = _RANDOM[11'h170][16];	// rob.scala:310:28
        rob_uop_26_ldst = _RANDOM[11'h170][23:18];	// rob.scala:310:28
        rob_uop_26_ldst_val = _RANDOM[11'h171][10];	// rob.scala:310:28
        rob_uop_26_dst_rtype = _RANDOM[11'h171][12:11];	// rob.scala:310:28
        rob_uop_26_fp_val = _RANDOM[11'h171][18];	// rob.scala:310:28
        rob_uop_27_uopc = {_RANDOM[11'h171][31:29], _RANDOM[11'h172][3:0]};	// rob.scala:310:28
        rob_uop_27_is_rvc = _RANDOM[11'h174][4];	// rob.scala:310:28
        rob_uop_27_br_mask = {_RANDOM[11'h176][31:25], _RANDOM[11'h177][12:0]};	// rob.scala:310:28
        rob_uop_27_ftq_idx = _RANDOM[11'h177][23:18];	// rob.scala:310:28
        rob_uop_27_edge_inst = _RANDOM[11'h177][24];	// rob.scala:310:28
        rob_uop_27_pc_lob = _RANDOM[11'h177][30:25];	// rob.scala:310:28
        rob_uop_27_pdst = _RANDOM[11'h179][25:19];	// rob.scala:310:28
        rob_uop_27_stale_pdst = _RANDOM[11'h17A][31:25];	// rob.scala:310:28
        rob_uop_27_is_fencei = _RANDOM[11'h17D][11];	// rob.scala:310:28
        rob_uop_27_uses_ldq = _RANDOM[11'h17D][13];	// rob.scala:310:28
        rob_uop_27_uses_stq = _RANDOM[11'h17D][14];	// rob.scala:310:28
        rob_uop_27_is_sys_pc2epc = _RANDOM[11'h17D][15];	// rob.scala:310:28
        rob_uop_27_flush_on_commit = _RANDOM[11'h17D][17];	// rob.scala:310:28
        rob_uop_27_ldst = _RANDOM[11'h17D][24:19];	// rob.scala:310:28
        rob_uop_27_ldst_val = _RANDOM[11'h17E][11];	// rob.scala:310:28
        rob_uop_27_dst_rtype = _RANDOM[11'h17E][13:12];	// rob.scala:310:28
        rob_uop_27_fp_val = _RANDOM[11'h17E][19];	// rob.scala:310:28
        rob_uop_28_uopc = {_RANDOM[11'h17E][31:30], _RANDOM[11'h17F][4:0]};	// rob.scala:310:28
        rob_uop_28_is_rvc = _RANDOM[11'h181][5];	// rob.scala:310:28
        rob_uop_28_br_mask = {_RANDOM[11'h183][31:26], _RANDOM[11'h184][13:0]};	// rob.scala:310:28
        rob_uop_28_ftq_idx = _RANDOM[11'h184][24:19];	// rob.scala:310:28
        rob_uop_28_edge_inst = _RANDOM[11'h184][25];	// rob.scala:310:28
        rob_uop_28_pc_lob = _RANDOM[11'h184][31:26];	// rob.scala:310:28
        rob_uop_28_pdst = _RANDOM[11'h186][26:20];	// rob.scala:310:28
        rob_uop_28_stale_pdst = {_RANDOM[11'h187][31:26], _RANDOM[11'h188][0]};	// rob.scala:310:28
        rob_uop_28_is_fencei = _RANDOM[11'h18A][12];	// rob.scala:310:28
        rob_uop_28_uses_ldq = _RANDOM[11'h18A][14];	// rob.scala:310:28
        rob_uop_28_uses_stq = _RANDOM[11'h18A][15];	// rob.scala:310:28
        rob_uop_28_is_sys_pc2epc = _RANDOM[11'h18A][16];	// rob.scala:310:28
        rob_uop_28_flush_on_commit = _RANDOM[11'h18A][18];	// rob.scala:310:28
        rob_uop_28_ldst = _RANDOM[11'h18A][25:20];	// rob.scala:310:28
        rob_uop_28_ldst_val = _RANDOM[11'h18B][12];	// rob.scala:310:28
        rob_uop_28_dst_rtype = _RANDOM[11'h18B][14:13];	// rob.scala:310:28
        rob_uop_28_fp_val = _RANDOM[11'h18B][20];	// rob.scala:310:28
        rob_uop_29_uopc = {_RANDOM[11'h18B][31], _RANDOM[11'h18C][5:0]};	// rob.scala:310:28
        rob_uop_29_is_rvc = _RANDOM[11'h18E][6];	// rob.scala:310:28
        rob_uop_29_br_mask = {_RANDOM[11'h190][31:27], _RANDOM[11'h191][14:0]};	// rob.scala:310:28
        rob_uop_29_ftq_idx = _RANDOM[11'h191][25:20];	// rob.scala:310:28
        rob_uop_29_edge_inst = _RANDOM[11'h191][26];	// rob.scala:310:28
        rob_uop_29_pc_lob = {_RANDOM[11'h191][31:27], _RANDOM[11'h192][0]};	// rob.scala:310:28
        rob_uop_29_pdst = _RANDOM[11'h193][27:21];	// rob.scala:310:28
        rob_uop_29_stale_pdst = {_RANDOM[11'h194][31:27], _RANDOM[11'h195][1:0]};	// rob.scala:310:28
        rob_uop_29_is_fencei = _RANDOM[11'h197][13];	// rob.scala:310:28
        rob_uop_29_uses_ldq = _RANDOM[11'h197][15];	// rob.scala:310:28
        rob_uop_29_uses_stq = _RANDOM[11'h197][16];	// rob.scala:310:28
        rob_uop_29_is_sys_pc2epc = _RANDOM[11'h197][17];	// rob.scala:310:28
        rob_uop_29_flush_on_commit = _RANDOM[11'h197][19];	// rob.scala:310:28
        rob_uop_29_ldst = _RANDOM[11'h197][26:21];	// rob.scala:310:28
        rob_uop_29_ldst_val = _RANDOM[11'h198][13];	// rob.scala:310:28
        rob_uop_29_dst_rtype = _RANDOM[11'h198][15:14];	// rob.scala:310:28
        rob_uop_29_fp_val = _RANDOM[11'h198][21];	// rob.scala:310:28
        rob_uop_30_uopc = _RANDOM[11'h199][6:0];	// rob.scala:310:28
        rob_uop_30_is_rvc = _RANDOM[11'h19B][7];	// rob.scala:310:28
        rob_uop_30_br_mask = {_RANDOM[11'h19D][31:28], _RANDOM[11'h19E][15:0]};	// rob.scala:310:28
        rob_uop_30_ftq_idx = _RANDOM[11'h19E][26:21];	// rob.scala:310:28
        rob_uop_30_edge_inst = _RANDOM[11'h19E][27];	// rob.scala:310:28
        rob_uop_30_pc_lob = {_RANDOM[11'h19E][31:28], _RANDOM[11'h19F][1:0]};	// rob.scala:310:28
        rob_uop_30_pdst = _RANDOM[11'h1A0][28:22];	// rob.scala:310:28
        rob_uop_30_stale_pdst = {_RANDOM[11'h1A1][31:28], _RANDOM[11'h1A2][2:0]};	// rob.scala:310:28
        rob_uop_30_is_fencei = _RANDOM[11'h1A4][14];	// rob.scala:310:28
        rob_uop_30_uses_ldq = _RANDOM[11'h1A4][16];	// rob.scala:310:28
        rob_uop_30_uses_stq = _RANDOM[11'h1A4][17];	// rob.scala:310:28
        rob_uop_30_is_sys_pc2epc = _RANDOM[11'h1A4][18];	// rob.scala:310:28
        rob_uop_30_flush_on_commit = _RANDOM[11'h1A4][20];	// rob.scala:310:28
        rob_uop_30_ldst = _RANDOM[11'h1A4][27:22];	// rob.scala:310:28
        rob_uop_30_ldst_val = _RANDOM[11'h1A5][14];	// rob.scala:310:28
        rob_uop_30_dst_rtype = _RANDOM[11'h1A5][16:15];	// rob.scala:310:28
        rob_uop_30_fp_val = _RANDOM[11'h1A5][22];	// rob.scala:310:28
        rob_uop_31_uopc = _RANDOM[11'h1A6][7:1];	// rob.scala:310:28
        rob_uop_31_is_rvc = _RANDOM[11'h1A8][8];	// rob.scala:310:28
        rob_uop_31_br_mask = {_RANDOM[11'h1AA][31:29], _RANDOM[11'h1AB][16:0]};	// rob.scala:310:28
        rob_uop_31_ftq_idx = _RANDOM[11'h1AB][27:22];	// rob.scala:310:28
        rob_uop_31_edge_inst = _RANDOM[11'h1AB][28];	// rob.scala:310:28
        rob_uop_31_pc_lob = {_RANDOM[11'h1AB][31:29], _RANDOM[11'h1AC][2:0]};	// rob.scala:310:28
        rob_uop_31_pdst = _RANDOM[11'h1AD][29:23];	// rob.scala:310:28
        rob_uop_31_stale_pdst = {_RANDOM[11'h1AE][31:29], _RANDOM[11'h1AF][3:0]};	// rob.scala:310:28
        rob_uop_31_is_fencei = _RANDOM[11'h1B1][15];	// rob.scala:310:28
        rob_uop_31_uses_ldq = _RANDOM[11'h1B1][17];	// rob.scala:310:28
        rob_uop_31_uses_stq = _RANDOM[11'h1B1][18];	// rob.scala:310:28
        rob_uop_31_is_sys_pc2epc = _RANDOM[11'h1B1][19];	// rob.scala:310:28
        rob_uop_31_flush_on_commit = _RANDOM[11'h1B1][21];	// rob.scala:310:28
        rob_uop_31_ldst = _RANDOM[11'h1B1][28:23];	// rob.scala:310:28
        rob_uop_31_ldst_val = _RANDOM[11'h1B2][15];	// rob.scala:310:28
        rob_uop_31_dst_rtype = _RANDOM[11'h1B2][17:16];	// rob.scala:310:28
        rob_uop_31_fp_val = _RANDOM[11'h1B2][23];	// rob.scala:310:28
        rob_exception_0 = _RANDOM[11'h1B3][2];	// rob.scala:311:28
        rob_exception_1 = _RANDOM[11'h1B3][3];	// rob.scala:311:28
        rob_exception_2 = _RANDOM[11'h1B3][4];	// rob.scala:311:28
        rob_exception_3 = _RANDOM[11'h1B3][5];	// rob.scala:311:28
        rob_exception_4 = _RANDOM[11'h1B3][6];	// rob.scala:311:28
        rob_exception_5 = _RANDOM[11'h1B3][7];	// rob.scala:311:28
        rob_exception_6 = _RANDOM[11'h1B3][8];	// rob.scala:311:28
        rob_exception_7 = _RANDOM[11'h1B3][9];	// rob.scala:311:28
        rob_exception_8 = _RANDOM[11'h1B3][10];	// rob.scala:311:28
        rob_exception_9 = _RANDOM[11'h1B3][11];	// rob.scala:311:28
        rob_exception_10 = _RANDOM[11'h1B3][12];	// rob.scala:311:28
        rob_exception_11 = _RANDOM[11'h1B3][13];	// rob.scala:311:28
        rob_exception_12 = _RANDOM[11'h1B3][14];	// rob.scala:311:28
        rob_exception_13 = _RANDOM[11'h1B3][15];	// rob.scala:311:28
        rob_exception_14 = _RANDOM[11'h1B3][16];	// rob.scala:311:28
        rob_exception_15 = _RANDOM[11'h1B3][17];	// rob.scala:311:28
        rob_exception_16 = _RANDOM[11'h1B3][18];	// rob.scala:311:28
        rob_exception_17 = _RANDOM[11'h1B3][19];	// rob.scala:311:28
        rob_exception_18 = _RANDOM[11'h1B3][20];	// rob.scala:311:28
        rob_exception_19 = _RANDOM[11'h1B3][21];	// rob.scala:311:28
        rob_exception_20 = _RANDOM[11'h1B3][22];	// rob.scala:311:28
        rob_exception_21 = _RANDOM[11'h1B3][23];	// rob.scala:311:28
        rob_exception_22 = _RANDOM[11'h1B3][24];	// rob.scala:311:28
        rob_exception_23 = _RANDOM[11'h1B3][25];	// rob.scala:311:28
        rob_exception_24 = _RANDOM[11'h1B3][26];	// rob.scala:311:28
        rob_exception_25 = _RANDOM[11'h1B3][27];	// rob.scala:311:28
        rob_exception_26 = _RANDOM[11'h1B3][28];	// rob.scala:311:28
        rob_exception_27 = _RANDOM[11'h1B3][29];	// rob.scala:311:28
        rob_exception_28 = _RANDOM[11'h1B3][30];	// rob.scala:311:28
        rob_exception_29 = _RANDOM[11'h1B3][31];	// rob.scala:311:28
        rob_exception_30 = _RANDOM[11'h1B4][0];	// rob.scala:311:28
        rob_exception_31 = _RANDOM[11'h1B4][1];	// rob.scala:311:28
        rob_predicated_0 = _RANDOM[11'h1B4][2];	// rob.scala:311:28, :312:29
        rob_predicated_1 = _RANDOM[11'h1B4][3];	// rob.scala:311:28, :312:29
        rob_predicated_2 = _RANDOM[11'h1B4][4];	// rob.scala:311:28, :312:29
        rob_predicated_3 = _RANDOM[11'h1B4][5];	// rob.scala:311:28, :312:29
        rob_predicated_4 = _RANDOM[11'h1B4][6];	// rob.scala:311:28, :312:29
        rob_predicated_5 = _RANDOM[11'h1B4][7];	// rob.scala:311:28, :312:29
        rob_predicated_6 = _RANDOM[11'h1B4][8];	// rob.scala:311:28, :312:29
        rob_predicated_7 = _RANDOM[11'h1B4][9];	// rob.scala:311:28, :312:29
        rob_predicated_8 = _RANDOM[11'h1B4][10];	// rob.scala:311:28, :312:29
        rob_predicated_9 = _RANDOM[11'h1B4][11];	// rob.scala:311:28, :312:29
        rob_predicated_10 = _RANDOM[11'h1B4][12];	// rob.scala:311:28, :312:29
        rob_predicated_11 = _RANDOM[11'h1B4][13];	// rob.scala:311:28, :312:29
        rob_predicated_12 = _RANDOM[11'h1B4][14];	// rob.scala:311:28, :312:29
        rob_predicated_13 = _RANDOM[11'h1B4][15];	// rob.scala:311:28, :312:29
        rob_predicated_14 = _RANDOM[11'h1B4][16];	// rob.scala:311:28, :312:29
        rob_predicated_15 = _RANDOM[11'h1B4][17];	// rob.scala:311:28, :312:29
        rob_predicated_16 = _RANDOM[11'h1B4][18];	// rob.scala:311:28, :312:29
        rob_predicated_17 = _RANDOM[11'h1B4][19];	// rob.scala:311:28, :312:29
        rob_predicated_18 = _RANDOM[11'h1B4][20];	// rob.scala:311:28, :312:29
        rob_predicated_19 = _RANDOM[11'h1B4][21];	// rob.scala:311:28, :312:29
        rob_predicated_20 = _RANDOM[11'h1B4][22];	// rob.scala:311:28, :312:29
        rob_predicated_21 = _RANDOM[11'h1B4][23];	// rob.scala:311:28, :312:29
        rob_predicated_22 = _RANDOM[11'h1B4][24];	// rob.scala:311:28, :312:29
        rob_predicated_23 = _RANDOM[11'h1B4][25];	// rob.scala:311:28, :312:29
        rob_predicated_24 = _RANDOM[11'h1B4][26];	// rob.scala:311:28, :312:29
        rob_predicated_25 = _RANDOM[11'h1B4][27];	// rob.scala:311:28, :312:29
        rob_predicated_26 = _RANDOM[11'h1B4][28];	// rob.scala:311:28, :312:29
        rob_predicated_27 = _RANDOM[11'h1B4][29];	// rob.scala:311:28, :312:29
        rob_predicated_28 = _RANDOM[11'h1B4][30];	// rob.scala:311:28, :312:29
        rob_predicated_29 = _RANDOM[11'h1B4][31];	// rob.scala:311:28, :312:29
        rob_predicated_30 = _RANDOM[11'h1B5][0];	// rob.scala:312:29
        rob_predicated_31 = _RANDOM[11'h1B5][1];	// rob.scala:312:29
        rob_val_1_0 = _RANDOM[11'h1B5][2];	// rob.scala:307:32, :312:29
        rob_val_1_1 = _RANDOM[11'h1B5][3];	// rob.scala:307:32, :312:29
        rob_val_1_2 = _RANDOM[11'h1B5][4];	// rob.scala:307:32, :312:29
        rob_val_1_3 = _RANDOM[11'h1B5][5];	// rob.scala:307:32, :312:29
        rob_val_1_4 = _RANDOM[11'h1B5][6];	// rob.scala:307:32, :312:29
        rob_val_1_5 = _RANDOM[11'h1B5][7];	// rob.scala:307:32, :312:29
        rob_val_1_6 = _RANDOM[11'h1B5][8];	// rob.scala:307:32, :312:29
        rob_val_1_7 = _RANDOM[11'h1B5][9];	// rob.scala:307:32, :312:29
        rob_val_1_8 = _RANDOM[11'h1B5][10];	// rob.scala:307:32, :312:29
        rob_val_1_9 = _RANDOM[11'h1B5][11];	// rob.scala:307:32, :312:29
        rob_val_1_10 = _RANDOM[11'h1B5][12];	// rob.scala:307:32, :312:29
        rob_val_1_11 = _RANDOM[11'h1B5][13];	// rob.scala:307:32, :312:29
        rob_val_1_12 = _RANDOM[11'h1B5][14];	// rob.scala:307:32, :312:29
        rob_val_1_13 = _RANDOM[11'h1B5][15];	// rob.scala:307:32, :312:29
        rob_val_1_14 = _RANDOM[11'h1B5][16];	// rob.scala:307:32, :312:29
        rob_val_1_15 = _RANDOM[11'h1B5][17];	// rob.scala:307:32, :312:29
        rob_val_1_16 = _RANDOM[11'h1B5][18];	// rob.scala:307:32, :312:29
        rob_val_1_17 = _RANDOM[11'h1B5][19];	// rob.scala:307:32, :312:29
        rob_val_1_18 = _RANDOM[11'h1B5][20];	// rob.scala:307:32, :312:29
        rob_val_1_19 = _RANDOM[11'h1B5][21];	// rob.scala:307:32, :312:29
        rob_val_1_20 = _RANDOM[11'h1B5][22];	// rob.scala:307:32, :312:29
        rob_val_1_21 = _RANDOM[11'h1B5][23];	// rob.scala:307:32, :312:29
        rob_val_1_22 = _RANDOM[11'h1B5][24];	// rob.scala:307:32, :312:29
        rob_val_1_23 = _RANDOM[11'h1B5][25];	// rob.scala:307:32, :312:29
        rob_val_1_24 = _RANDOM[11'h1B5][26];	// rob.scala:307:32, :312:29
        rob_val_1_25 = _RANDOM[11'h1B5][27];	// rob.scala:307:32, :312:29
        rob_val_1_26 = _RANDOM[11'h1B5][28];	// rob.scala:307:32, :312:29
        rob_val_1_27 = _RANDOM[11'h1B5][29];	// rob.scala:307:32, :312:29
        rob_val_1_28 = _RANDOM[11'h1B5][30];	// rob.scala:307:32, :312:29
        rob_val_1_29 = _RANDOM[11'h1B5][31];	// rob.scala:307:32, :312:29
        rob_val_1_30 = _RANDOM[11'h1B6][0];	// rob.scala:307:32
        rob_val_1_31 = _RANDOM[11'h1B6][1];	// rob.scala:307:32
        rob_bsy_1_0 = _RANDOM[11'h1B6][2];	// rob.scala:307:32, :308:28
        rob_bsy_1_1 = _RANDOM[11'h1B6][3];	// rob.scala:307:32, :308:28
        rob_bsy_1_2 = _RANDOM[11'h1B6][4];	// rob.scala:307:32, :308:28
        rob_bsy_1_3 = _RANDOM[11'h1B6][5];	// rob.scala:307:32, :308:28
        rob_bsy_1_4 = _RANDOM[11'h1B6][6];	// rob.scala:307:32, :308:28
        rob_bsy_1_5 = _RANDOM[11'h1B6][7];	// rob.scala:307:32, :308:28
        rob_bsy_1_6 = _RANDOM[11'h1B6][8];	// rob.scala:307:32, :308:28
        rob_bsy_1_7 = _RANDOM[11'h1B6][9];	// rob.scala:307:32, :308:28
        rob_bsy_1_8 = _RANDOM[11'h1B6][10];	// rob.scala:307:32, :308:28
        rob_bsy_1_9 = _RANDOM[11'h1B6][11];	// rob.scala:307:32, :308:28
        rob_bsy_1_10 = _RANDOM[11'h1B6][12];	// rob.scala:307:32, :308:28
        rob_bsy_1_11 = _RANDOM[11'h1B6][13];	// rob.scala:307:32, :308:28
        rob_bsy_1_12 = _RANDOM[11'h1B6][14];	// rob.scala:307:32, :308:28
        rob_bsy_1_13 = _RANDOM[11'h1B6][15];	// rob.scala:307:32, :308:28
        rob_bsy_1_14 = _RANDOM[11'h1B6][16];	// rob.scala:307:32, :308:28
        rob_bsy_1_15 = _RANDOM[11'h1B6][17];	// rob.scala:307:32, :308:28
        rob_bsy_1_16 = _RANDOM[11'h1B6][18];	// rob.scala:307:32, :308:28
        rob_bsy_1_17 = _RANDOM[11'h1B6][19];	// rob.scala:307:32, :308:28
        rob_bsy_1_18 = _RANDOM[11'h1B6][20];	// rob.scala:307:32, :308:28
        rob_bsy_1_19 = _RANDOM[11'h1B6][21];	// rob.scala:307:32, :308:28
        rob_bsy_1_20 = _RANDOM[11'h1B6][22];	// rob.scala:307:32, :308:28
        rob_bsy_1_21 = _RANDOM[11'h1B6][23];	// rob.scala:307:32, :308:28
        rob_bsy_1_22 = _RANDOM[11'h1B6][24];	// rob.scala:307:32, :308:28
        rob_bsy_1_23 = _RANDOM[11'h1B6][25];	// rob.scala:307:32, :308:28
        rob_bsy_1_24 = _RANDOM[11'h1B6][26];	// rob.scala:307:32, :308:28
        rob_bsy_1_25 = _RANDOM[11'h1B6][27];	// rob.scala:307:32, :308:28
        rob_bsy_1_26 = _RANDOM[11'h1B6][28];	// rob.scala:307:32, :308:28
        rob_bsy_1_27 = _RANDOM[11'h1B6][29];	// rob.scala:307:32, :308:28
        rob_bsy_1_28 = _RANDOM[11'h1B6][30];	// rob.scala:307:32, :308:28
        rob_bsy_1_29 = _RANDOM[11'h1B6][31];	// rob.scala:307:32, :308:28
        rob_bsy_1_30 = _RANDOM[11'h1B7][0];	// rob.scala:308:28
        rob_bsy_1_31 = _RANDOM[11'h1B7][1];	// rob.scala:308:28
        rob_unsafe_1_0 = _RANDOM[11'h1B7][2];	// rob.scala:308:28, :309:28
        rob_unsafe_1_1 = _RANDOM[11'h1B7][3];	// rob.scala:308:28, :309:28
        rob_unsafe_1_2 = _RANDOM[11'h1B7][4];	// rob.scala:308:28, :309:28
        rob_unsafe_1_3 = _RANDOM[11'h1B7][5];	// rob.scala:308:28, :309:28
        rob_unsafe_1_4 = _RANDOM[11'h1B7][6];	// rob.scala:308:28, :309:28
        rob_unsafe_1_5 = _RANDOM[11'h1B7][7];	// rob.scala:308:28, :309:28
        rob_unsafe_1_6 = _RANDOM[11'h1B7][8];	// rob.scala:308:28, :309:28
        rob_unsafe_1_7 = _RANDOM[11'h1B7][9];	// rob.scala:308:28, :309:28
        rob_unsafe_1_8 = _RANDOM[11'h1B7][10];	// rob.scala:308:28, :309:28
        rob_unsafe_1_9 = _RANDOM[11'h1B7][11];	// rob.scala:308:28, :309:28
        rob_unsafe_1_10 = _RANDOM[11'h1B7][12];	// rob.scala:308:28, :309:28
        rob_unsafe_1_11 = _RANDOM[11'h1B7][13];	// rob.scala:308:28, :309:28
        rob_unsafe_1_12 = _RANDOM[11'h1B7][14];	// rob.scala:308:28, :309:28
        rob_unsafe_1_13 = _RANDOM[11'h1B7][15];	// rob.scala:308:28, :309:28
        rob_unsafe_1_14 = _RANDOM[11'h1B7][16];	// rob.scala:308:28, :309:28
        rob_unsafe_1_15 = _RANDOM[11'h1B7][17];	// rob.scala:308:28, :309:28
        rob_unsafe_1_16 = _RANDOM[11'h1B7][18];	// rob.scala:308:28, :309:28
        rob_unsafe_1_17 = _RANDOM[11'h1B7][19];	// rob.scala:308:28, :309:28
        rob_unsafe_1_18 = _RANDOM[11'h1B7][20];	// rob.scala:308:28, :309:28
        rob_unsafe_1_19 = _RANDOM[11'h1B7][21];	// rob.scala:308:28, :309:28
        rob_unsafe_1_20 = _RANDOM[11'h1B7][22];	// rob.scala:308:28, :309:28
        rob_unsafe_1_21 = _RANDOM[11'h1B7][23];	// rob.scala:308:28, :309:28
        rob_unsafe_1_22 = _RANDOM[11'h1B7][24];	// rob.scala:308:28, :309:28
        rob_unsafe_1_23 = _RANDOM[11'h1B7][25];	// rob.scala:308:28, :309:28
        rob_unsafe_1_24 = _RANDOM[11'h1B7][26];	// rob.scala:308:28, :309:28
        rob_unsafe_1_25 = _RANDOM[11'h1B7][27];	// rob.scala:308:28, :309:28
        rob_unsafe_1_26 = _RANDOM[11'h1B7][28];	// rob.scala:308:28, :309:28
        rob_unsafe_1_27 = _RANDOM[11'h1B7][29];	// rob.scala:308:28, :309:28
        rob_unsafe_1_28 = _RANDOM[11'h1B7][30];	// rob.scala:308:28, :309:28
        rob_unsafe_1_29 = _RANDOM[11'h1B7][31];	// rob.scala:308:28, :309:28
        rob_unsafe_1_30 = _RANDOM[11'h1B8][0];	// rob.scala:309:28
        rob_unsafe_1_31 = _RANDOM[11'h1B8][1];	// rob.scala:309:28
        rob_uop_1_0_uopc = _RANDOM[11'h1B8][8:2];	// rob.scala:309:28, :310:28
        rob_uop_1_0_is_rvc = _RANDOM[11'h1BA][9];	// rob.scala:310:28
        rob_uop_1_0_br_mask = {_RANDOM[11'h1BC][31:30], _RANDOM[11'h1BD][17:0]};	// rob.scala:310:28
        rob_uop_1_0_ftq_idx = _RANDOM[11'h1BD][28:23];	// rob.scala:310:28
        rob_uop_1_0_edge_inst = _RANDOM[11'h1BD][29];	// rob.scala:310:28
        rob_uop_1_0_pc_lob = {_RANDOM[11'h1BD][31:30], _RANDOM[11'h1BE][3:0]};	// rob.scala:310:28
        rob_uop_1_0_pdst = _RANDOM[11'h1BF][30:24];	// rob.scala:310:28
        rob_uop_1_0_stale_pdst = {_RANDOM[11'h1C0][31:30], _RANDOM[11'h1C1][4:0]};	// rob.scala:310:28
        rob_uop_1_0_is_fencei = _RANDOM[11'h1C3][16];	// rob.scala:310:28
        rob_uop_1_0_uses_ldq = _RANDOM[11'h1C3][18];	// rob.scala:310:28
        rob_uop_1_0_uses_stq = _RANDOM[11'h1C3][19];	// rob.scala:310:28
        rob_uop_1_0_is_sys_pc2epc = _RANDOM[11'h1C3][20];	// rob.scala:310:28
        rob_uop_1_0_flush_on_commit = _RANDOM[11'h1C3][22];	// rob.scala:310:28
        rob_uop_1_0_ldst = _RANDOM[11'h1C3][29:24];	// rob.scala:310:28
        rob_uop_1_0_ldst_val = _RANDOM[11'h1C4][16];	// rob.scala:310:28
        rob_uop_1_0_dst_rtype = _RANDOM[11'h1C4][18:17];	// rob.scala:310:28
        rob_uop_1_0_fp_val = _RANDOM[11'h1C4][24];	// rob.scala:310:28
        rob_uop_1_1_uopc = _RANDOM[11'h1C5][9:3];	// rob.scala:310:28
        rob_uop_1_1_is_rvc = _RANDOM[11'h1C7][10];	// rob.scala:310:28
        rob_uop_1_1_br_mask = {_RANDOM[11'h1C9][31], _RANDOM[11'h1CA][18:0]};	// rob.scala:310:28
        rob_uop_1_1_ftq_idx = _RANDOM[11'h1CA][29:24];	// rob.scala:310:28
        rob_uop_1_1_edge_inst = _RANDOM[11'h1CA][30];	// rob.scala:310:28
        rob_uop_1_1_pc_lob = {_RANDOM[11'h1CA][31], _RANDOM[11'h1CB][4:0]};	// rob.scala:310:28
        rob_uop_1_1_pdst = _RANDOM[11'h1CC][31:25];	// rob.scala:310:28
        rob_uop_1_1_stale_pdst = {_RANDOM[11'h1CD][31], _RANDOM[11'h1CE][5:0]};	// rob.scala:310:28
        rob_uop_1_1_is_fencei = _RANDOM[11'h1D0][17];	// rob.scala:310:28
        rob_uop_1_1_uses_ldq = _RANDOM[11'h1D0][19];	// rob.scala:310:28
        rob_uop_1_1_uses_stq = _RANDOM[11'h1D0][20];	// rob.scala:310:28
        rob_uop_1_1_is_sys_pc2epc = _RANDOM[11'h1D0][21];	// rob.scala:310:28
        rob_uop_1_1_flush_on_commit = _RANDOM[11'h1D0][23];	// rob.scala:310:28
        rob_uop_1_1_ldst = _RANDOM[11'h1D0][30:25];	// rob.scala:310:28
        rob_uop_1_1_ldst_val = _RANDOM[11'h1D1][17];	// rob.scala:310:28
        rob_uop_1_1_dst_rtype = _RANDOM[11'h1D1][19:18];	// rob.scala:310:28
        rob_uop_1_1_fp_val = _RANDOM[11'h1D1][25];	// rob.scala:310:28
        rob_uop_1_2_uopc = _RANDOM[11'h1D2][10:4];	// rob.scala:310:28
        rob_uop_1_2_is_rvc = _RANDOM[11'h1D4][11];	// rob.scala:310:28
        rob_uop_1_2_br_mask = _RANDOM[11'h1D7][19:0];	// rob.scala:310:28
        rob_uop_1_2_ftq_idx = _RANDOM[11'h1D7][30:25];	// rob.scala:310:28
        rob_uop_1_2_edge_inst = _RANDOM[11'h1D7][31];	// rob.scala:310:28
        rob_uop_1_2_pc_lob = _RANDOM[11'h1D8][5:0];	// rob.scala:310:28
        rob_uop_1_2_pdst = {_RANDOM[11'h1D9][31:26], _RANDOM[11'h1DA][0]};	// rob.scala:310:28
        rob_uop_1_2_stale_pdst = _RANDOM[11'h1DB][6:0];	// rob.scala:310:28
        rob_uop_1_2_is_fencei = _RANDOM[11'h1DD][18];	// rob.scala:310:28
        rob_uop_1_2_uses_ldq = _RANDOM[11'h1DD][20];	// rob.scala:310:28
        rob_uop_1_2_uses_stq = _RANDOM[11'h1DD][21];	// rob.scala:310:28
        rob_uop_1_2_is_sys_pc2epc = _RANDOM[11'h1DD][22];	// rob.scala:310:28
        rob_uop_1_2_flush_on_commit = _RANDOM[11'h1DD][24];	// rob.scala:310:28
        rob_uop_1_2_ldst = _RANDOM[11'h1DD][31:26];	// rob.scala:310:28
        rob_uop_1_2_ldst_val = _RANDOM[11'h1DE][18];	// rob.scala:310:28
        rob_uop_1_2_dst_rtype = _RANDOM[11'h1DE][20:19];	// rob.scala:310:28
        rob_uop_1_2_fp_val = _RANDOM[11'h1DE][26];	// rob.scala:310:28
        rob_uop_1_3_uopc = _RANDOM[11'h1DF][11:5];	// rob.scala:310:28
        rob_uop_1_3_is_rvc = _RANDOM[11'h1E1][12];	// rob.scala:310:28
        rob_uop_1_3_br_mask = _RANDOM[11'h1E4][20:1];	// rob.scala:310:28
        rob_uop_1_3_ftq_idx = _RANDOM[11'h1E4][31:26];	// rob.scala:310:28
        rob_uop_1_3_edge_inst = _RANDOM[11'h1E5][0];	// rob.scala:310:28
        rob_uop_1_3_pc_lob = _RANDOM[11'h1E5][6:1];	// rob.scala:310:28
        rob_uop_1_3_pdst = {_RANDOM[11'h1E6][31:27], _RANDOM[11'h1E7][1:0]};	// rob.scala:310:28
        rob_uop_1_3_stale_pdst = _RANDOM[11'h1E8][7:1];	// rob.scala:310:28
        rob_uop_1_3_is_fencei = _RANDOM[11'h1EA][19];	// rob.scala:310:28
        rob_uop_1_3_uses_ldq = _RANDOM[11'h1EA][21];	// rob.scala:310:28
        rob_uop_1_3_uses_stq = _RANDOM[11'h1EA][22];	// rob.scala:310:28
        rob_uop_1_3_is_sys_pc2epc = _RANDOM[11'h1EA][23];	// rob.scala:310:28
        rob_uop_1_3_flush_on_commit = _RANDOM[11'h1EA][25];	// rob.scala:310:28
        rob_uop_1_3_ldst = {_RANDOM[11'h1EA][31:27], _RANDOM[11'h1EB][0]};	// rob.scala:310:28
        rob_uop_1_3_ldst_val = _RANDOM[11'h1EB][19];	// rob.scala:310:28
        rob_uop_1_3_dst_rtype = _RANDOM[11'h1EB][21:20];	// rob.scala:310:28
        rob_uop_1_3_fp_val = _RANDOM[11'h1EB][27];	// rob.scala:310:28
        rob_uop_1_4_uopc = _RANDOM[11'h1EC][12:6];	// rob.scala:310:28
        rob_uop_1_4_is_rvc = _RANDOM[11'h1EE][13];	// rob.scala:310:28
        rob_uop_1_4_br_mask = _RANDOM[11'h1F1][21:2];	// rob.scala:310:28
        rob_uop_1_4_ftq_idx = {_RANDOM[11'h1F1][31:27], _RANDOM[11'h1F2][0]};	// rob.scala:310:28
        rob_uop_1_4_edge_inst = _RANDOM[11'h1F2][1];	// rob.scala:310:28
        rob_uop_1_4_pc_lob = _RANDOM[11'h1F2][7:2];	// rob.scala:310:28
        rob_uop_1_4_pdst = {_RANDOM[11'h1F3][31:28], _RANDOM[11'h1F4][2:0]};	// rob.scala:310:28
        rob_uop_1_4_stale_pdst = _RANDOM[11'h1F5][8:2];	// rob.scala:310:28
        rob_uop_1_4_is_fencei = _RANDOM[11'h1F7][20];	// rob.scala:310:28
        rob_uop_1_4_uses_ldq = _RANDOM[11'h1F7][22];	// rob.scala:310:28
        rob_uop_1_4_uses_stq = _RANDOM[11'h1F7][23];	// rob.scala:310:28
        rob_uop_1_4_is_sys_pc2epc = _RANDOM[11'h1F7][24];	// rob.scala:310:28
        rob_uop_1_4_flush_on_commit = _RANDOM[11'h1F7][26];	// rob.scala:310:28
        rob_uop_1_4_ldst = {_RANDOM[11'h1F7][31:28], _RANDOM[11'h1F8][1:0]};	// rob.scala:310:28
        rob_uop_1_4_ldst_val = _RANDOM[11'h1F8][20];	// rob.scala:310:28
        rob_uop_1_4_dst_rtype = _RANDOM[11'h1F8][22:21];	// rob.scala:310:28
        rob_uop_1_4_fp_val = _RANDOM[11'h1F8][28];	// rob.scala:310:28
        rob_uop_1_5_uopc = _RANDOM[11'h1F9][13:7];	// rob.scala:310:28
        rob_uop_1_5_is_rvc = _RANDOM[11'h1FB][14];	// rob.scala:310:28
        rob_uop_1_5_br_mask = _RANDOM[11'h1FE][22:3];	// rob.scala:310:28
        rob_uop_1_5_ftq_idx = {_RANDOM[11'h1FE][31:28], _RANDOM[11'h1FF][1:0]};	// rob.scala:310:28
        rob_uop_1_5_edge_inst = _RANDOM[11'h1FF][2];	// rob.scala:310:28
        rob_uop_1_5_pc_lob = _RANDOM[11'h1FF][8:3];	// rob.scala:310:28
        rob_uop_1_5_pdst = {_RANDOM[11'h200][31:29], _RANDOM[11'h201][3:0]};	// rob.scala:310:28
        rob_uop_1_5_stale_pdst = _RANDOM[11'h202][9:3];	// rob.scala:310:28
        rob_uop_1_5_is_fencei = _RANDOM[11'h204][21];	// rob.scala:310:28
        rob_uop_1_5_uses_ldq = _RANDOM[11'h204][23];	// rob.scala:310:28
        rob_uop_1_5_uses_stq = _RANDOM[11'h204][24];	// rob.scala:310:28
        rob_uop_1_5_is_sys_pc2epc = _RANDOM[11'h204][25];	// rob.scala:310:28
        rob_uop_1_5_flush_on_commit = _RANDOM[11'h204][27];	// rob.scala:310:28
        rob_uop_1_5_ldst = {_RANDOM[11'h204][31:29], _RANDOM[11'h205][2:0]};	// rob.scala:310:28
        rob_uop_1_5_ldst_val = _RANDOM[11'h205][21];	// rob.scala:310:28
        rob_uop_1_5_dst_rtype = _RANDOM[11'h205][23:22];	// rob.scala:310:28
        rob_uop_1_5_fp_val = _RANDOM[11'h205][29];	// rob.scala:310:28
        rob_uop_1_6_uopc = _RANDOM[11'h206][14:8];	// rob.scala:310:28
        rob_uop_1_6_is_rvc = _RANDOM[11'h208][15];	// rob.scala:310:28
        rob_uop_1_6_br_mask = _RANDOM[11'h20B][23:4];	// rob.scala:310:28
        rob_uop_1_6_ftq_idx = {_RANDOM[11'h20B][31:29], _RANDOM[11'h20C][2:0]};	// rob.scala:310:28
        rob_uop_1_6_edge_inst = _RANDOM[11'h20C][3];	// rob.scala:310:28
        rob_uop_1_6_pc_lob = _RANDOM[11'h20C][9:4];	// rob.scala:310:28
        rob_uop_1_6_pdst = {_RANDOM[11'h20D][31:30], _RANDOM[11'h20E][4:0]};	// rob.scala:310:28
        rob_uop_1_6_stale_pdst = _RANDOM[11'h20F][10:4];	// rob.scala:310:28
        rob_uop_1_6_is_fencei = _RANDOM[11'h211][22];	// rob.scala:310:28
        rob_uop_1_6_uses_ldq = _RANDOM[11'h211][24];	// rob.scala:310:28
        rob_uop_1_6_uses_stq = _RANDOM[11'h211][25];	// rob.scala:310:28
        rob_uop_1_6_is_sys_pc2epc = _RANDOM[11'h211][26];	// rob.scala:310:28
        rob_uop_1_6_flush_on_commit = _RANDOM[11'h211][28];	// rob.scala:310:28
        rob_uop_1_6_ldst = {_RANDOM[11'h211][31:30], _RANDOM[11'h212][3:0]};	// rob.scala:310:28
        rob_uop_1_6_ldst_val = _RANDOM[11'h212][22];	// rob.scala:310:28
        rob_uop_1_6_dst_rtype = _RANDOM[11'h212][24:23];	// rob.scala:310:28
        rob_uop_1_6_fp_val = _RANDOM[11'h212][30];	// rob.scala:310:28
        rob_uop_1_7_uopc = _RANDOM[11'h213][15:9];	// rob.scala:310:28
        rob_uop_1_7_is_rvc = _RANDOM[11'h215][16];	// rob.scala:310:28
        rob_uop_1_7_br_mask = _RANDOM[11'h218][24:5];	// rob.scala:310:28
        rob_uop_1_7_ftq_idx = {_RANDOM[11'h218][31:30], _RANDOM[11'h219][3:0]};	// rob.scala:310:28
        rob_uop_1_7_edge_inst = _RANDOM[11'h219][4];	// rob.scala:310:28
        rob_uop_1_7_pc_lob = _RANDOM[11'h219][10:5];	// rob.scala:310:28
        rob_uop_1_7_pdst = {_RANDOM[11'h21A][31], _RANDOM[11'h21B][5:0]};	// rob.scala:310:28
        rob_uop_1_7_stale_pdst = _RANDOM[11'h21C][11:5];	// rob.scala:310:28
        rob_uop_1_7_is_fencei = _RANDOM[11'h21E][23];	// rob.scala:310:28
        rob_uop_1_7_uses_ldq = _RANDOM[11'h21E][25];	// rob.scala:310:28
        rob_uop_1_7_uses_stq = _RANDOM[11'h21E][26];	// rob.scala:310:28
        rob_uop_1_7_is_sys_pc2epc = _RANDOM[11'h21E][27];	// rob.scala:310:28
        rob_uop_1_7_flush_on_commit = _RANDOM[11'h21E][29];	// rob.scala:310:28
        rob_uop_1_7_ldst = {_RANDOM[11'h21E][31], _RANDOM[11'h21F][4:0]};	// rob.scala:310:28
        rob_uop_1_7_ldst_val = _RANDOM[11'h21F][23];	// rob.scala:310:28
        rob_uop_1_7_dst_rtype = _RANDOM[11'h21F][25:24];	// rob.scala:310:28
        rob_uop_1_7_fp_val = _RANDOM[11'h21F][31];	// rob.scala:310:28
        rob_uop_1_8_uopc = _RANDOM[11'h220][16:10];	// rob.scala:310:28
        rob_uop_1_8_is_rvc = _RANDOM[11'h222][17];	// rob.scala:310:28
        rob_uop_1_8_br_mask = _RANDOM[11'h225][25:6];	// rob.scala:310:28
        rob_uop_1_8_ftq_idx = {_RANDOM[11'h225][31], _RANDOM[11'h226][4:0]};	// rob.scala:310:28
        rob_uop_1_8_edge_inst = _RANDOM[11'h226][5];	// rob.scala:310:28
        rob_uop_1_8_pc_lob = _RANDOM[11'h226][11:6];	// rob.scala:310:28
        rob_uop_1_8_pdst = _RANDOM[11'h228][6:0];	// rob.scala:310:28
        rob_uop_1_8_stale_pdst = _RANDOM[11'h229][12:6];	// rob.scala:310:28
        rob_uop_1_8_is_fencei = _RANDOM[11'h22B][24];	// rob.scala:310:28
        rob_uop_1_8_uses_ldq = _RANDOM[11'h22B][26];	// rob.scala:310:28
        rob_uop_1_8_uses_stq = _RANDOM[11'h22B][27];	// rob.scala:310:28
        rob_uop_1_8_is_sys_pc2epc = _RANDOM[11'h22B][28];	// rob.scala:310:28
        rob_uop_1_8_flush_on_commit = _RANDOM[11'h22B][30];	// rob.scala:310:28
        rob_uop_1_8_ldst = _RANDOM[11'h22C][5:0];	// rob.scala:310:28
        rob_uop_1_8_ldst_val = _RANDOM[11'h22C][24];	// rob.scala:310:28
        rob_uop_1_8_dst_rtype = _RANDOM[11'h22C][26:25];	// rob.scala:310:28
        rob_uop_1_8_fp_val = _RANDOM[11'h22D][0];	// rob.scala:310:28
        rob_uop_1_9_uopc = _RANDOM[11'h22D][17:11];	// rob.scala:310:28
        rob_uop_1_9_is_rvc = _RANDOM[11'h22F][18];	// rob.scala:310:28
        rob_uop_1_9_br_mask = _RANDOM[11'h232][26:7];	// rob.scala:310:28
        rob_uop_1_9_ftq_idx = _RANDOM[11'h233][5:0];	// rob.scala:310:28
        rob_uop_1_9_edge_inst = _RANDOM[11'h233][6];	// rob.scala:310:28
        rob_uop_1_9_pc_lob = _RANDOM[11'h233][12:7];	// rob.scala:310:28
        rob_uop_1_9_pdst = _RANDOM[11'h235][7:1];	// rob.scala:310:28
        rob_uop_1_9_stale_pdst = _RANDOM[11'h236][13:7];	// rob.scala:310:28
        rob_uop_1_9_is_fencei = _RANDOM[11'h238][25];	// rob.scala:310:28
        rob_uop_1_9_uses_ldq = _RANDOM[11'h238][27];	// rob.scala:310:28
        rob_uop_1_9_uses_stq = _RANDOM[11'h238][28];	// rob.scala:310:28
        rob_uop_1_9_is_sys_pc2epc = _RANDOM[11'h238][29];	// rob.scala:310:28
        rob_uop_1_9_flush_on_commit = _RANDOM[11'h238][31];	// rob.scala:310:28
        rob_uop_1_9_ldst = _RANDOM[11'h239][6:1];	// rob.scala:310:28
        rob_uop_1_9_ldst_val = _RANDOM[11'h239][25];	// rob.scala:310:28
        rob_uop_1_9_dst_rtype = _RANDOM[11'h239][27:26];	// rob.scala:310:28
        rob_uop_1_9_fp_val = _RANDOM[11'h23A][1];	// rob.scala:310:28
        rob_uop_1_10_uopc = _RANDOM[11'h23A][18:12];	// rob.scala:310:28
        rob_uop_1_10_is_rvc = _RANDOM[11'h23C][19];	// rob.scala:310:28
        rob_uop_1_10_br_mask = _RANDOM[11'h23F][27:8];	// rob.scala:310:28
        rob_uop_1_10_ftq_idx = _RANDOM[11'h240][6:1];	// rob.scala:310:28
        rob_uop_1_10_edge_inst = _RANDOM[11'h240][7];	// rob.scala:310:28
        rob_uop_1_10_pc_lob = _RANDOM[11'h240][13:8];	// rob.scala:310:28
        rob_uop_1_10_pdst = _RANDOM[11'h242][8:2];	// rob.scala:310:28
        rob_uop_1_10_stale_pdst = _RANDOM[11'h243][14:8];	// rob.scala:310:28
        rob_uop_1_10_is_fencei = _RANDOM[11'h245][26];	// rob.scala:310:28
        rob_uop_1_10_uses_ldq = _RANDOM[11'h245][28];	// rob.scala:310:28
        rob_uop_1_10_uses_stq = _RANDOM[11'h245][29];	// rob.scala:310:28
        rob_uop_1_10_is_sys_pc2epc = _RANDOM[11'h245][30];	// rob.scala:310:28
        rob_uop_1_10_flush_on_commit = _RANDOM[11'h246][0];	// rob.scala:310:28
        rob_uop_1_10_ldst = _RANDOM[11'h246][7:2];	// rob.scala:310:28
        rob_uop_1_10_ldst_val = _RANDOM[11'h246][26];	// rob.scala:310:28
        rob_uop_1_10_dst_rtype = _RANDOM[11'h246][28:27];	// rob.scala:310:28
        rob_uop_1_10_fp_val = _RANDOM[11'h247][2];	// rob.scala:310:28
        rob_uop_1_11_uopc = _RANDOM[11'h247][19:13];	// rob.scala:310:28
        rob_uop_1_11_is_rvc = _RANDOM[11'h249][20];	// rob.scala:310:28
        rob_uop_1_11_br_mask = _RANDOM[11'h24C][28:9];	// rob.scala:310:28
        rob_uop_1_11_ftq_idx = _RANDOM[11'h24D][7:2];	// rob.scala:310:28
        rob_uop_1_11_edge_inst = _RANDOM[11'h24D][8];	// rob.scala:310:28
        rob_uop_1_11_pc_lob = _RANDOM[11'h24D][14:9];	// rob.scala:310:28
        rob_uop_1_11_pdst = _RANDOM[11'h24F][9:3];	// rob.scala:310:28
        rob_uop_1_11_stale_pdst = _RANDOM[11'h250][15:9];	// rob.scala:310:28
        rob_uop_1_11_is_fencei = _RANDOM[11'h252][27];	// rob.scala:310:28
        rob_uop_1_11_uses_ldq = _RANDOM[11'h252][29];	// rob.scala:310:28
        rob_uop_1_11_uses_stq = _RANDOM[11'h252][30];	// rob.scala:310:28
        rob_uop_1_11_is_sys_pc2epc = _RANDOM[11'h252][31];	// rob.scala:310:28
        rob_uop_1_11_flush_on_commit = _RANDOM[11'h253][1];	// rob.scala:310:28
        rob_uop_1_11_ldst = _RANDOM[11'h253][8:3];	// rob.scala:310:28
        rob_uop_1_11_ldst_val = _RANDOM[11'h253][27];	// rob.scala:310:28
        rob_uop_1_11_dst_rtype = _RANDOM[11'h253][29:28];	// rob.scala:310:28
        rob_uop_1_11_fp_val = _RANDOM[11'h254][3];	// rob.scala:310:28
        rob_uop_1_12_uopc = _RANDOM[11'h254][20:14];	// rob.scala:310:28
        rob_uop_1_12_is_rvc = _RANDOM[11'h256][21];	// rob.scala:310:28
        rob_uop_1_12_br_mask = _RANDOM[11'h259][29:10];	// rob.scala:310:28
        rob_uop_1_12_ftq_idx = _RANDOM[11'h25A][8:3];	// rob.scala:310:28
        rob_uop_1_12_edge_inst = _RANDOM[11'h25A][9];	// rob.scala:310:28
        rob_uop_1_12_pc_lob = _RANDOM[11'h25A][15:10];	// rob.scala:310:28
        rob_uop_1_12_pdst = _RANDOM[11'h25C][10:4];	// rob.scala:310:28
        rob_uop_1_12_stale_pdst = _RANDOM[11'h25D][16:10];	// rob.scala:310:28
        rob_uop_1_12_is_fencei = _RANDOM[11'h25F][28];	// rob.scala:310:28
        rob_uop_1_12_uses_ldq = _RANDOM[11'h25F][30];	// rob.scala:310:28
        rob_uop_1_12_uses_stq = _RANDOM[11'h25F][31];	// rob.scala:310:28
        rob_uop_1_12_is_sys_pc2epc = _RANDOM[11'h260][0];	// rob.scala:310:28
        rob_uop_1_12_flush_on_commit = _RANDOM[11'h260][2];	// rob.scala:310:28
        rob_uop_1_12_ldst = _RANDOM[11'h260][9:4];	// rob.scala:310:28
        rob_uop_1_12_ldst_val = _RANDOM[11'h260][28];	// rob.scala:310:28
        rob_uop_1_12_dst_rtype = _RANDOM[11'h260][30:29];	// rob.scala:310:28
        rob_uop_1_12_fp_val = _RANDOM[11'h261][4];	// rob.scala:310:28
        rob_uop_1_13_uopc = _RANDOM[11'h261][21:15];	// rob.scala:310:28
        rob_uop_1_13_is_rvc = _RANDOM[11'h263][22];	// rob.scala:310:28
        rob_uop_1_13_br_mask = _RANDOM[11'h266][30:11];	// rob.scala:310:28
        rob_uop_1_13_ftq_idx = _RANDOM[11'h267][9:4];	// rob.scala:310:28
        rob_uop_1_13_edge_inst = _RANDOM[11'h267][10];	// rob.scala:310:28
        rob_uop_1_13_pc_lob = _RANDOM[11'h267][16:11];	// rob.scala:310:28
        rob_uop_1_13_pdst = _RANDOM[11'h269][11:5];	// rob.scala:310:28
        rob_uop_1_13_stale_pdst = _RANDOM[11'h26A][17:11];	// rob.scala:310:28
        rob_uop_1_13_is_fencei = _RANDOM[11'h26C][29];	// rob.scala:310:28
        rob_uop_1_13_uses_ldq = _RANDOM[11'h26C][31];	// rob.scala:310:28
        rob_uop_1_13_uses_stq = _RANDOM[11'h26D][0];	// rob.scala:310:28
        rob_uop_1_13_is_sys_pc2epc = _RANDOM[11'h26D][1];	// rob.scala:310:28
        rob_uop_1_13_flush_on_commit = _RANDOM[11'h26D][3];	// rob.scala:310:28
        rob_uop_1_13_ldst = _RANDOM[11'h26D][10:5];	// rob.scala:310:28
        rob_uop_1_13_ldst_val = _RANDOM[11'h26D][29];	// rob.scala:310:28
        rob_uop_1_13_dst_rtype = _RANDOM[11'h26D][31:30];	// rob.scala:310:28
        rob_uop_1_13_fp_val = _RANDOM[11'h26E][5];	// rob.scala:310:28
        rob_uop_1_14_uopc = _RANDOM[11'h26E][22:16];	// rob.scala:310:28
        rob_uop_1_14_is_rvc = _RANDOM[11'h270][23];	// rob.scala:310:28
        rob_uop_1_14_br_mask = _RANDOM[11'h273][31:12];	// rob.scala:310:28
        rob_uop_1_14_ftq_idx = _RANDOM[11'h274][10:5];	// rob.scala:310:28
        rob_uop_1_14_edge_inst = _RANDOM[11'h274][11];	// rob.scala:310:28
        rob_uop_1_14_pc_lob = _RANDOM[11'h274][17:12];	// rob.scala:310:28
        rob_uop_1_14_pdst = _RANDOM[11'h276][12:6];	// rob.scala:310:28
        rob_uop_1_14_stale_pdst = _RANDOM[11'h277][18:12];	// rob.scala:310:28
        rob_uop_1_14_is_fencei = _RANDOM[11'h279][30];	// rob.scala:310:28
        rob_uop_1_14_uses_ldq = _RANDOM[11'h27A][0];	// rob.scala:310:28
        rob_uop_1_14_uses_stq = _RANDOM[11'h27A][1];	// rob.scala:310:28
        rob_uop_1_14_is_sys_pc2epc = _RANDOM[11'h27A][2];	// rob.scala:310:28
        rob_uop_1_14_flush_on_commit = _RANDOM[11'h27A][4];	// rob.scala:310:28
        rob_uop_1_14_ldst = _RANDOM[11'h27A][11:6];	// rob.scala:310:28
        rob_uop_1_14_ldst_val = _RANDOM[11'h27A][30];	// rob.scala:310:28
        rob_uop_1_14_dst_rtype = {_RANDOM[11'h27A][31], _RANDOM[11'h27B][0]};	// rob.scala:310:28
        rob_uop_1_14_fp_val = _RANDOM[11'h27B][6];	// rob.scala:310:28
        rob_uop_1_15_uopc = _RANDOM[11'h27B][23:17];	// rob.scala:310:28
        rob_uop_1_15_is_rvc = _RANDOM[11'h27D][24];	// rob.scala:310:28
        rob_uop_1_15_br_mask = {_RANDOM[11'h280][31:13], _RANDOM[11'h281][0]};	// rob.scala:310:28
        rob_uop_1_15_ftq_idx = _RANDOM[11'h281][11:6];	// rob.scala:310:28
        rob_uop_1_15_edge_inst = _RANDOM[11'h281][12];	// rob.scala:310:28
        rob_uop_1_15_pc_lob = _RANDOM[11'h281][18:13];	// rob.scala:310:28
        rob_uop_1_15_pdst = _RANDOM[11'h283][13:7];	// rob.scala:310:28
        rob_uop_1_15_stale_pdst = _RANDOM[11'h284][19:13];	// rob.scala:310:28
        rob_uop_1_15_is_fencei = _RANDOM[11'h286][31];	// rob.scala:310:28
        rob_uop_1_15_uses_ldq = _RANDOM[11'h287][1];	// rob.scala:310:28
        rob_uop_1_15_uses_stq = _RANDOM[11'h287][2];	// rob.scala:310:28
        rob_uop_1_15_is_sys_pc2epc = _RANDOM[11'h287][3];	// rob.scala:310:28
        rob_uop_1_15_flush_on_commit = _RANDOM[11'h287][5];	// rob.scala:310:28
        rob_uop_1_15_ldst = _RANDOM[11'h287][12:7];	// rob.scala:310:28
        rob_uop_1_15_ldst_val = _RANDOM[11'h287][31];	// rob.scala:310:28
        rob_uop_1_15_dst_rtype = _RANDOM[11'h288][1:0];	// rob.scala:310:28
        rob_uop_1_15_fp_val = _RANDOM[11'h288][7];	// rob.scala:310:28
        rob_uop_1_16_uopc = _RANDOM[11'h288][24:18];	// rob.scala:310:28
        rob_uop_1_16_is_rvc = _RANDOM[11'h28A][25];	// rob.scala:310:28
        rob_uop_1_16_br_mask = {_RANDOM[11'h28D][31:14], _RANDOM[11'h28E][1:0]};	// rob.scala:310:28
        rob_uop_1_16_ftq_idx = _RANDOM[11'h28E][12:7];	// rob.scala:310:28
        rob_uop_1_16_edge_inst = _RANDOM[11'h28E][13];	// rob.scala:310:28
        rob_uop_1_16_pc_lob = _RANDOM[11'h28E][19:14];	// rob.scala:310:28
        rob_uop_1_16_pdst = _RANDOM[11'h290][14:8];	// rob.scala:310:28
        rob_uop_1_16_stale_pdst = _RANDOM[11'h291][20:14];	// rob.scala:310:28
        rob_uop_1_16_is_fencei = _RANDOM[11'h294][0];	// rob.scala:310:28
        rob_uop_1_16_uses_ldq = _RANDOM[11'h294][2];	// rob.scala:310:28
        rob_uop_1_16_uses_stq = _RANDOM[11'h294][3];	// rob.scala:310:28
        rob_uop_1_16_is_sys_pc2epc = _RANDOM[11'h294][4];	// rob.scala:310:28
        rob_uop_1_16_flush_on_commit = _RANDOM[11'h294][6];	// rob.scala:310:28
        rob_uop_1_16_ldst = _RANDOM[11'h294][13:8];	// rob.scala:310:28
        rob_uop_1_16_ldst_val = _RANDOM[11'h295][0];	// rob.scala:310:28
        rob_uop_1_16_dst_rtype = _RANDOM[11'h295][2:1];	// rob.scala:310:28
        rob_uop_1_16_fp_val = _RANDOM[11'h295][8];	// rob.scala:310:28
        rob_uop_1_17_uopc = _RANDOM[11'h295][25:19];	// rob.scala:310:28
        rob_uop_1_17_is_rvc = _RANDOM[11'h297][26];	// rob.scala:310:28
        rob_uop_1_17_br_mask = {_RANDOM[11'h29A][31:15], _RANDOM[11'h29B][2:0]};	// rob.scala:310:28
        rob_uop_1_17_ftq_idx = _RANDOM[11'h29B][13:8];	// rob.scala:310:28
        rob_uop_1_17_edge_inst = _RANDOM[11'h29B][14];	// rob.scala:310:28
        rob_uop_1_17_pc_lob = _RANDOM[11'h29B][20:15];	// rob.scala:310:28
        rob_uop_1_17_pdst = _RANDOM[11'h29D][15:9];	// rob.scala:310:28
        rob_uop_1_17_stale_pdst = _RANDOM[11'h29E][21:15];	// rob.scala:310:28
        rob_uop_1_17_is_fencei = _RANDOM[11'h2A1][1];	// rob.scala:310:28
        rob_uop_1_17_uses_ldq = _RANDOM[11'h2A1][3];	// rob.scala:310:28
        rob_uop_1_17_uses_stq = _RANDOM[11'h2A1][4];	// rob.scala:310:28
        rob_uop_1_17_is_sys_pc2epc = _RANDOM[11'h2A1][5];	// rob.scala:310:28
        rob_uop_1_17_flush_on_commit = _RANDOM[11'h2A1][7];	// rob.scala:310:28
        rob_uop_1_17_ldst = _RANDOM[11'h2A1][14:9];	// rob.scala:310:28
        rob_uop_1_17_ldst_val = _RANDOM[11'h2A2][1];	// rob.scala:310:28
        rob_uop_1_17_dst_rtype = _RANDOM[11'h2A2][3:2];	// rob.scala:310:28
        rob_uop_1_17_fp_val = _RANDOM[11'h2A2][9];	// rob.scala:310:28
        rob_uop_1_18_uopc = _RANDOM[11'h2A2][26:20];	// rob.scala:310:28
        rob_uop_1_18_is_rvc = _RANDOM[11'h2A4][27];	// rob.scala:310:28
        rob_uop_1_18_br_mask = {_RANDOM[11'h2A7][31:16], _RANDOM[11'h2A8][3:0]};	// rob.scala:310:28
        rob_uop_1_18_ftq_idx = _RANDOM[11'h2A8][14:9];	// rob.scala:310:28
        rob_uop_1_18_edge_inst = _RANDOM[11'h2A8][15];	// rob.scala:310:28
        rob_uop_1_18_pc_lob = _RANDOM[11'h2A8][21:16];	// rob.scala:310:28
        rob_uop_1_18_pdst = _RANDOM[11'h2AA][16:10];	// rob.scala:310:28
        rob_uop_1_18_stale_pdst = _RANDOM[11'h2AB][22:16];	// rob.scala:310:28
        rob_uop_1_18_is_fencei = _RANDOM[11'h2AE][2];	// rob.scala:310:28
        rob_uop_1_18_uses_ldq = _RANDOM[11'h2AE][4];	// rob.scala:310:28
        rob_uop_1_18_uses_stq = _RANDOM[11'h2AE][5];	// rob.scala:310:28
        rob_uop_1_18_is_sys_pc2epc = _RANDOM[11'h2AE][6];	// rob.scala:310:28
        rob_uop_1_18_flush_on_commit = _RANDOM[11'h2AE][8];	// rob.scala:310:28
        rob_uop_1_18_ldst = _RANDOM[11'h2AE][15:10];	// rob.scala:310:28
        rob_uop_1_18_ldst_val = _RANDOM[11'h2AF][2];	// rob.scala:310:28
        rob_uop_1_18_dst_rtype = _RANDOM[11'h2AF][4:3];	// rob.scala:310:28
        rob_uop_1_18_fp_val = _RANDOM[11'h2AF][10];	// rob.scala:310:28
        rob_uop_1_19_uopc = _RANDOM[11'h2AF][27:21];	// rob.scala:310:28
        rob_uop_1_19_is_rvc = _RANDOM[11'h2B1][28];	// rob.scala:310:28
        rob_uop_1_19_br_mask = {_RANDOM[11'h2B4][31:17], _RANDOM[11'h2B5][4:0]};	// rob.scala:310:28
        rob_uop_1_19_ftq_idx = _RANDOM[11'h2B5][15:10];	// rob.scala:310:28
        rob_uop_1_19_edge_inst = _RANDOM[11'h2B5][16];	// rob.scala:310:28
        rob_uop_1_19_pc_lob = _RANDOM[11'h2B5][22:17];	// rob.scala:310:28
        rob_uop_1_19_pdst = _RANDOM[11'h2B7][17:11];	// rob.scala:310:28
        rob_uop_1_19_stale_pdst = _RANDOM[11'h2B8][23:17];	// rob.scala:310:28
        rob_uop_1_19_is_fencei = _RANDOM[11'h2BB][3];	// rob.scala:310:28
        rob_uop_1_19_uses_ldq = _RANDOM[11'h2BB][5];	// rob.scala:310:28
        rob_uop_1_19_uses_stq = _RANDOM[11'h2BB][6];	// rob.scala:310:28
        rob_uop_1_19_is_sys_pc2epc = _RANDOM[11'h2BB][7];	// rob.scala:310:28
        rob_uop_1_19_flush_on_commit = _RANDOM[11'h2BB][9];	// rob.scala:310:28
        rob_uop_1_19_ldst = _RANDOM[11'h2BB][16:11];	// rob.scala:310:28
        rob_uop_1_19_ldst_val = _RANDOM[11'h2BC][3];	// rob.scala:310:28
        rob_uop_1_19_dst_rtype = _RANDOM[11'h2BC][5:4];	// rob.scala:310:28
        rob_uop_1_19_fp_val = _RANDOM[11'h2BC][11];	// rob.scala:310:28
        rob_uop_1_20_uopc = _RANDOM[11'h2BC][28:22];	// rob.scala:310:28
        rob_uop_1_20_is_rvc = _RANDOM[11'h2BE][29];	// rob.scala:310:28
        rob_uop_1_20_br_mask = {_RANDOM[11'h2C1][31:18], _RANDOM[11'h2C2][5:0]};	// rob.scala:310:28
        rob_uop_1_20_ftq_idx = _RANDOM[11'h2C2][16:11];	// rob.scala:310:28
        rob_uop_1_20_edge_inst = _RANDOM[11'h2C2][17];	// rob.scala:310:28
        rob_uop_1_20_pc_lob = _RANDOM[11'h2C2][23:18];	// rob.scala:310:28
        rob_uop_1_20_pdst = _RANDOM[11'h2C4][18:12];	// rob.scala:310:28
        rob_uop_1_20_stale_pdst = _RANDOM[11'h2C5][24:18];	// rob.scala:310:28
        rob_uop_1_20_is_fencei = _RANDOM[11'h2C8][4];	// rob.scala:310:28
        rob_uop_1_20_uses_ldq = _RANDOM[11'h2C8][6];	// rob.scala:310:28
        rob_uop_1_20_uses_stq = _RANDOM[11'h2C8][7];	// rob.scala:310:28
        rob_uop_1_20_is_sys_pc2epc = _RANDOM[11'h2C8][8];	// rob.scala:310:28
        rob_uop_1_20_flush_on_commit = _RANDOM[11'h2C8][10];	// rob.scala:310:28
        rob_uop_1_20_ldst = _RANDOM[11'h2C8][17:12];	// rob.scala:310:28
        rob_uop_1_20_ldst_val = _RANDOM[11'h2C9][4];	// rob.scala:310:28
        rob_uop_1_20_dst_rtype = _RANDOM[11'h2C9][6:5];	// rob.scala:310:28
        rob_uop_1_20_fp_val = _RANDOM[11'h2C9][12];	// rob.scala:310:28
        rob_uop_1_21_uopc = _RANDOM[11'h2C9][29:23];	// rob.scala:310:28
        rob_uop_1_21_is_rvc = _RANDOM[11'h2CB][30];	// rob.scala:310:28
        rob_uop_1_21_br_mask = {_RANDOM[11'h2CE][31:19], _RANDOM[11'h2CF][6:0]};	// rob.scala:310:28
        rob_uop_1_21_ftq_idx = _RANDOM[11'h2CF][17:12];	// rob.scala:310:28
        rob_uop_1_21_edge_inst = _RANDOM[11'h2CF][18];	// rob.scala:310:28
        rob_uop_1_21_pc_lob = _RANDOM[11'h2CF][24:19];	// rob.scala:310:28
        rob_uop_1_21_pdst = _RANDOM[11'h2D1][19:13];	// rob.scala:310:28
        rob_uop_1_21_stale_pdst = _RANDOM[11'h2D2][25:19];	// rob.scala:310:28
        rob_uop_1_21_is_fencei = _RANDOM[11'h2D5][5];	// rob.scala:310:28
        rob_uop_1_21_uses_ldq = _RANDOM[11'h2D5][7];	// rob.scala:310:28
        rob_uop_1_21_uses_stq = _RANDOM[11'h2D5][8];	// rob.scala:310:28
        rob_uop_1_21_is_sys_pc2epc = _RANDOM[11'h2D5][9];	// rob.scala:310:28
        rob_uop_1_21_flush_on_commit = _RANDOM[11'h2D5][11];	// rob.scala:310:28
        rob_uop_1_21_ldst = _RANDOM[11'h2D5][18:13];	// rob.scala:310:28
        rob_uop_1_21_ldst_val = _RANDOM[11'h2D6][5];	// rob.scala:310:28
        rob_uop_1_21_dst_rtype = _RANDOM[11'h2D6][7:6];	// rob.scala:310:28
        rob_uop_1_21_fp_val = _RANDOM[11'h2D6][13];	// rob.scala:310:28
        rob_uop_1_22_uopc = _RANDOM[11'h2D6][30:24];	// rob.scala:310:28
        rob_uop_1_22_is_rvc = _RANDOM[11'h2D8][31];	// rob.scala:310:28
        rob_uop_1_22_br_mask = {_RANDOM[11'h2DB][31:20], _RANDOM[11'h2DC][7:0]};	// rob.scala:310:28
        rob_uop_1_22_ftq_idx = _RANDOM[11'h2DC][18:13];	// rob.scala:310:28
        rob_uop_1_22_edge_inst = _RANDOM[11'h2DC][19];	// rob.scala:310:28
        rob_uop_1_22_pc_lob = _RANDOM[11'h2DC][25:20];	// rob.scala:310:28
        rob_uop_1_22_pdst = _RANDOM[11'h2DE][20:14];	// rob.scala:310:28
        rob_uop_1_22_stale_pdst = _RANDOM[11'h2DF][26:20];	// rob.scala:310:28
        rob_uop_1_22_is_fencei = _RANDOM[11'h2E2][6];	// rob.scala:310:28
        rob_uop_1_22_uses_ldq = _RANDOM[11'h2E2][8];	// rob.scala:310:28
        rob_uop_1_22_uses_stq = _RANDOM[11'h2E2][9];	// rob.scala:310:28
        rob_uop_1_22_is_sys_pc2epc = _RANDOM[11'h2E2][10];	// rob.scala:310:28
        rob_uop_1_22_flush_on_commit = _RANDOM[11'h2E2][12];	// rob.scala:310:28
        rob_uop_1_22_ldst = _RANDOM[11'h2E2][19:14];	// rob.scala:310:28
        rob_uop_1_22_ldst_val = _RANDOM[11'h2E3][6];	// rob.scala:310:28
        rob_uop_1_22_dst_rtype = _RANDOM[11'h2E3][8:7];	// rob.scala:310:28
        rob_uop_1_22_fp_val = _RANDOM[11'h2E3][14];	// rob.scala:310:28
        rob_uop_1_23_uopc = _RANDOM[11'h2E3][31:25];	// rob.scala:310:28
        rob_uop_1_23_is_rvc = _RANDOM[11'h2E6][0];	// rob.scala:310:28
        rob_uop_1_23_br_mask = {_RANDOM[11'h2E8][31:21], _RANDOM[11'h2E9][8:0]};	// rob.scala:310:28
        rob_uop_1_23_ftq_idx = _RANDOM[11'h2E9][19:14];	// rob.scala:310:28
        rob_uop_1_23_edge_inst = _RANDOM[11'h2E9][20];	// rob.scala:310:28
        rob_uop_1_23_pc_lob = _RANDOM[11'h2E9][26:21];	// rob.scala:310:28
        rob_uop_1_23_pdst = _RANDOM[11'h2EB][21:15];	// rob.scala:310:28
        rob_uop_1_23_stale_pdst = _RANDOM[11'h2EC][27:21];	// rob.scala:310:28
        rob_uop_1_23_is_fencei = _RANDOM[11'h2EF][7];	// rob.scala:310:28
        rob_uop_1_23_uses_ldq = _RANDOM[11'h2EF][9];	// rob.scala:310:28
        rob_uop_1_23_uses_stq = _RANDOM[11'h2EF][10];	// rob.scala:310:28
        rob_uop_1_23_is_sys_pc2epc = _RANDOM[11'h2EF][11];	// rob.scala:310:28
        rob_uop_1_23_flush_on_commit = _RANDOM[11'h2EF][13];	// rob.scala:310:28
        rob_uop_1_23_ldst = _RANDOM[11'h2EF][20:15];	// rob.scala:310:28
        rob_uop_1_23_ldst_val = _RANDOM[11'h2F0][7];	// rob.scala:310:28
        rob_uop_1_23_dst_rtype = _RANDOM[11'h2F0][9:8];	// rob.scala:310:28
        rob_uop_1_23_fp_val = _RANDOM[11'h2F0][15];	// rob.scala:310:28
        rob_uop_1_24_uopc = {_RANDOM[11'h2F0][31:26], _RANDOM[11'h2F1][0]};	// rob.scala:310:28
        rob_uop_1_24_is_rvc = _RANDOM[11'h2F3][1];	// rob.scala:310:28
        rob_uop_1_24_br_mask = {_RANDOM[11'h2F5][31:22], _RANDOM[11'h2F6][9:0]};	// rob.scala:310:28
        rob_uop_1_24_ftq_idx = _RANDOM[11'h2F6][20:15];	// rob.scala:310:28
        rob_uop_1_24_edge_inst = _RANDOM[11'h2F6][21];	// rob.scala:310:28
        rob_uop_1_24_pc_lob = _RANDOM[11'h2F6][27:22];	// rob.scala:310:28
        rob_uop_1_24_pdst = _RANDOM[11'h2F8][22:16];	// rob.scala:310:28
        rob_uop_1_24_stale_pdst = _RANDOM[11'h2F9][28:22];	// rob.scala:310:28
        rob_uop_1_24_is_fencei = _RANDOM[11'h2FC][8];	// rob.scala:310:28
        rob_uop_1_24_uses_ldq = _RANDOM[11'h2FC][10];	// rob.scala:310:28
        rob_uop_1_24_uses_stq = _RANDOM[11'h2FC][11];	// rob.scala:310:28
        rob_uop_1_24_is_sys_pc2epc = _RANDOM[11'h2FC][12];	// rob.scala:310:28
        rob_uop_1_24_flush_on_commit = _RANDOM[11'h2FC][14];	// rob.scala:310:28
        rob_uop_1_24_ldst = _RANDOM[11'h2FC][21:16];	// rob.scala:310:28
        rob_uop_1_24_ldst_val = _RANDOM[11'h2FD][8];	// rob.scala:310:28
        rob_uop_1_24_dst_rtype = _RANDOM[11'h2FD][10:9];	// rob.scala:310:28
        rob_uop_1_24_fp_val = _RANDOM[11'h2FD][16];	// rob.scala:310:28
        rob_uop_1_25_uopc = {_RANDOM[11'h2FD][31:27], _RANDOM[11'h2FE][1:0]};	// rob.scala:310:28
        rob_uop_1_25_is_rvc = _RANDOM[11'h300][2];	// rob.scala:310:28
        rob_uop_1_25_br_mask = {_RANDOM[11'h302][31:23], _RANDOM[11'h303][10:0]};	// rob.scala:310:28
        rob_uop_1_25_ftq_idx = _RANDOM[11'h303][21:16];	// rob.scala:310:28
        rob_uop_1_25_edge_inst = _RANDOM[11'h303][22];	// rob.scala:310:28
        rob_uop_1_25_pc_lob = _RANDOM[11'h303][28:23];	// rob.scala:310:28
        rob_uop_1_25_pdst = _RANDOM[11'h305][23:17];	// rob.scala:310:28
        rob_uop_1_25_stale_pdst = _RANDOM[11'h306][29:23];	// rob.scala:310:28
        rob_uop_1_25_is_fencei = _RANDOM[11'h309][9];	// rob.scala:310:28
        rob_uop_1_25_uses_ldq = _RANDOM[11'h309][11];	// rob.scala:310:28
        rob_uop_1_25_uses_stq = _RANDOM[11'h309][12];	// rob.scala:310:28
        rob_uop_1_25_is_sys_pc2epc = _RANDOM[11'h309][13];	// rob.scala:310:28
        rob_uop_1_25_flush_on_commit = _RANDOM[11'h309][15];	// rob.scala:310:28
        rob_uop_1_25_ldst = _RANDOM[11'h309][22:17];	// rob.scala:310:28
        rob_uop_1_25_ldst_val = _RANDOM[11'h30A][9];	// rob.scala:310:28
        rob_uop_1_25_dst_rtype = _RANDOM[11'h30A][11:10];	// rob.scala:310:28
        rob_uop_1_25_fp_val = _RANDOM[11'h30A][17];	// rob.scala:310:28
        rob_uop_1_26_uopc = {_RANDOM[11'h30A][31:28], _RANDOM[11'h30B][2:0]};	// rob.scala:310:28
        rob_uop_1_26_is_rvc = _RANDOM[11'h30D][3];	// rob.scala:310:28
        rob_uop_1_26_br_mask = {_RANDOM[11'h30F][31:24], _RANDOM[11'h310][11:0]};	// rob.scala:310:28
        rob_uop_1_26_ftq_idx = _RANDOM[11'h310][22:17];	// rob.scala:310:28
        rob_uop_1_26_edge_inst = _RANDOM[11'h310][23];	// rob.scala:310:28
        rob_uop_1_26_pc_lob = _RANDOM[11'h310][29:24];	// rob.scala:310:28
        rob_uop_1_26_pdst = _RANDOM[11'h312][24:18];	// rob.scala:310:28
        rob_uop_1_26_stale_pdst = _RANDOM[11'h313][30:24];	// rob.scala:310:28
        rob_uop_1_26_is_fencei = _RANDOM[11'h316][10];	// rob.scala:310:28
        rob_uop_1_26_uses_ldq = _RANDOM[11'h316][12];	// rob.scala:310:28
        rob_uop_1_26_uses_stq = _RANDOM[11'h316][13];	// rob.scala:310:28
        rob_uop_1_26_is_sys_pc2epc = _RANDOM[11'h316][14];	// rob.scala:310:28
        rob_uop_1_26_flush_on_commit = _RANDOM[11'h316][16];	// rob.scala:310:28
        rob_uop_1_26_ldst = _RANDOM[11'h316][23:18];	// rob.scala:310:28
        rob_uop_1_26_ldst_val = _RANDOM[11'h317][10];	// rob.scala:310:28
        rob_uop_1_26_dst_rtype = _RANDOM[11'h317][12:11];	// rob.scala:310:28
        rob_uop_1_26_fp_val = _RANDOM[11'h317][18];	// rob.scala:310:28
        rob_uop_1_27_uopc = {_RANDOM[11'h317][31:29], _RANDOM[11'h318][3:0]};	// rob.scala:310:28
        rob_uop_1_27_is_rvc = _RANDOM[11'h31A][4];	// rob.scala:310:28
        rob_uop_1_27_br_mask = {_RANDOM[11'h31C][31:25], _RANDOM[11'h31D][12:0]};	// rob.scala:310:28
        rob_uop_1_27_ftq_idx = _RANDOM[11'h31D][23:18];	// rob.scala:310:28
        rob_uop_1_27_edge_inst = _RANDOM[11'h31D][24];	// rob.scala:310:28
        rob_uop_1_27_pc_lob = _RANDOM[11'h31D][30:25];	// rob.scala:310:28
        rob_uop_1_27_pdst = _RANDOM[11'h31F][25:19];	// rob.scala:310:28
        rob_uop_1_27_stale_pdst = _RANDOM[11'h320][31:25];	// rob.scala:310:28
        rob_uop_1_27_is_fencei = _RANDOM[11'h323][11];	// rob.scala:310:28
        rob_uop_1_27_uses_ldq = _RANDOM[11'h323][13];	// rob.scala:310:28
        rob_uop_1_27_uses_stq = _RANDOM[11'h323][14];	// rob.scala:310:28
        rob_uop_1_27_is_sys_pc2epc = _RANDOM[11'h323][15];	// rob.scala:310:28
        rob_uop_1_27_flush_on_commit = _RANDOM[11'h323][17];	// rob.scala:310:28
        rob_uop_1_27_ldst = _RANDOM[11'h323][24:19];	// rob.scala:310:28
        rob_uop_1_27_ldst_val = _RANDOM[11'h324][11];	// rob.scala:310:28
        rob_uop_1_27_dst_rtype = _RANDOM[11'h324][13:12];	// rob.scala:310:28
        rob_uop_1_27_fp_val = _RANDOM[11'h324][19];	// rob.scala:310:28
        rob_uop_1_28_uopc = {_RANDOM[11'h324][31:30], _RANDOM[11'h325][4:0]};	// rob.scala:310:28
        rob_uop_1_28_is_rvc = _RANDOM[11'h327][5];	// rob.scala:310:28
        rob_uop_1_28_br_mask = {_RANDOM[11'h329][31:26], _RANDOM[11'h32A][13:0]};	// rob.scala:310:28
        rob_uop_1_28_ftq_idx = _RANDOM[11'h32A][24:19];	// rob.scala:310:28
        rob_uop_1_28_edge_inst = _RANDOM[11'h32A][25];	// rob.scala:310:28
        rob_uop_1_28_pc_lob = _RANDOM[11'h32A][31:26];	// rob.scala:310:28
        rob_uop_1_28_pdst = _RANDOM[11'h32C][26:20];	// rob.scala:310:28
        rob_uop_1_28_stale_pdst = {_RANDOM[11'h32D][31:26], _RANDOM[11'h32E][0]};	// rob.scala:310:28
        rob_uop_1_28_is_fencei = _RANDOM[11'h330][12];	// rob.scala:310:28
        rob_uop_1_28_uses_ldq = _RANDOM[11'h330][14];	// rob.scala:310:28
        rob_uop_1_28_uses_stq = _RANDOM[11'h330][15];	// rob.scala:310:28
        rob_uop_1_28_is_sys_pc2epc = _RANDOM[11'h330][16];	// rob.scala:310:28
        rob_uop_1_28_flush_on_commit = _RANDOM[11'h330][18];	// rob.scala:310:28
        rob_uop_1_28_ldst = _RANDOM[11'h330][25:20];	// rob.scala:310:28
        rob_uop_1_28_ldst_val = _RANDOM[11'h331][12];	// rob.scala:310:28
        rob_uop_1_28_dst_rtype = _RANDOM[11'h331][14:13];	// rob.scala:310:28
        rob_uop_1_28_fp_val = _RANDOM[11'h331][20];	// rob.scala:310:28
        rob_uop_1_29_uopc = {_RANDOM[11'h331][31], _RANDOM[11'h332][5:0]};	// rob.scala:310:28
        rob_uop_1_29_is_rvc = _RANDOM[11'h334][6];	// rob.scala:310:28
        rob_uop_1_29_br_mask = {_RANDOM[11'h336][31:27], _RANDOM[11'h337][14:0]};	// rob.scala:310:28
        rob_uop_1_29_ftq_idx = _RANDOM[11'h337][25:20];	// rob.scala:310:28
        rob_uop_1_29_edge_inst = _RANDOM[11'h337][26];	// rob.scala:310:28
        rob_uop_1_29_pc_lob = {_RANDOM[11'h337][31:27], _RANDOM[11'h338][0]};	// rob.scala:310:28
        rob_uop_1_29_pdst = _RANDOM[11'h339][27:21];	// rob.scala:310:28
        rob_uop_1_29_stale_pdst = {_RANDOM[11'h33A][31:27], _RANDOM[11'h33B][1:0]};	// rob.scala:310:28
        rob_uop_1_29_is_fencei = _RANDOM[11'h33D][13];	// rob.scala:310:28
        rob_uop_1_29_uses_ldq = _RANDOM[11'h33D][15];	// rob.scala:310:28
        rob_uop_1_29_uses_stq = _RANDOM[11'h33D][16];	// rob.scala:310:28
        rob_uop_1_29_is_sys_pc2epc = _RANDOM[11'h33D][17];	// rob.scala:310:28
        rob_uop_1_29_flush_on_commit = _RANDOM[11'h33D][19];	// rob.scala:310:28
        rob_uop_1_29_ldst = _RANDOM[11'h33D][26:21];	// rob.scala:310:28
        rob_uop_1_29_ldst_val = _RANDOM[11'h33E][13];	// rob.scala:310:28
        rob_uop_1_29_dst_rtype = _RANDOM[11'h33E][15:14];	// rob.scala:310:28
        rob_uop_1_29_fp_val = _RANDOM[11'h33E][21];	// rob.scala:310:28
        rob_uop_1_30_uopc = _RANDOM[11'h33F][6:0];	// rob.scala:310:28
        rob_uop_1_30_is_rvc = _RANDOM[11'h341][7];	// rob.scala:310:28
        rob_uop_1_30_br_mask = {_RANDOM[11'h343][31:28], _RANDOM[11'h344][15:0]};	// rob.scala:310:28
        rob_uop_1_30_ftq_idx = _RANDOM[11'h344][26:21];	// rob.scala:310:28
        rob_uop_1_30_edge_inst = _RANDOM[11'h344][27];	// rob.scala:310:28
        rob_uop_1_30_pc_lob = {_RANDOM[11'h344][31:28], _RANDOM[11'h345][1:0]};	// rob.scala:310:28
        rob_uop_1_30_pdst = _RANDOM[11'h346][28:22];	// rob.scala:310:28
        rob_uop_1_30_stale_pdst = {_RANDOM[11'h347][31:28], _RANDOM[11'h348][2:0]};	// rob.scala:310:28
        rob_uop_1_30_is_fencei = _RANDOM[11'h34A][14];	// rob.scala:310:28
        rob_uop_1_30_uses_ldq = _RANDOM[11'h34A][16];	// rob.scala:310:28
        rob_uop_1_30_uses_stq = _RANDOM[11'h34A][17];	// rob.scala:310:28
        rob_uop_1_30_is_sys_pc2epc = _RANDOM[11'h34A][18];	// rob.scala:310:28
        rob_uop_1_30_flush_on_commit = _RANDOM[11'h34A][20];	// rob.scala:310:28
        rob_uop_1_30_ldst = _RANDOM[11'h34A][27:22];	// rob.scala:310:28
        rob_uop_1_30_ldst_val = _RANDOM[11'h34B][14];	// rob.scala:310:28
        rob_uop_1_30_dst_rtype = _RANDOM[11'h34B][16:15];	// rob.scala:310:28
        rob_uop_1_30_fp_val = _RANDOM[11'h34B][22];	// rob.scala:310:28
        rob_uop_1_31_uopc = _RANDOM[11'h34C][7:1];	// rob.scala:310:28
        rob_uop_1_31_is_rvc = _RANDOM[11'h34E][8];	// rob.scala:310:28
        rob_uop_1_31_br_mask = {_RANDOM[11'h350][31:29], _RANDOM[11'h351][16:0]};	// rob.scala:310:28
        rob_uop_1_31_ftq_idx = _RANDOM[11'h351][27:22];	// rob.scala:310:28
        rob_uop_1_31_edge_inst = _RANDOM[11'h351][28];	// rob.scala:310:28
        rob_uop_1_31_pc_lob = {_RANDOM[11'h351][31:29], _RANDOM[11'h352][2:0]};	// rob.scala:310:28
        rob_uop_1_31_pdst = _RANDOM[11'h353][29:23];	// rob.scala:310:28
        rob_uop_1_31_stale_pdst = {_RANDOM[11'h354][31:29], _RANDOM[11'h355][3:0]};	// rob.scala:310:28
        rob_uop_1_31_is_fencei = _RANDOM[11'h357][15];	// rob.scala:310:28
        rob_uop_1_31_uses_ldq = _RANDOM[11'h357][17];	// rob.scala:310:28
        rob_uop_1_31_uses_stq = _RANDOM[11'h357][18];	// rob.scala:310:28
        rob_uop_1_31_is_sys_pc2epc = _RANDOM[11'h357][19];	// rob.scala:310:28
        rob_uop_1_31_flush_on_commit = _RANDOM[11'h357][21];	// rob.scala:310:28
        rob_uop_1_31_ldst = _RANDOM[11'h357][28:23];	// rob.scala:310:28
        rob_uop_1_31_ldst_val = _RANDOM[11'h358][15];	// rob.scala:310:28
        rob_uop_1_31_dst_rtype = _RANDOM[11'h358][17:16];	// rob.scala:310:28
        rob_uop_1_31_fp_val = _RANDOM[11'h358][23];	// rob.scala:310:28
        rob_exception_1_0 = _RANDOM[11'h359][2];	// rob.scala:311:28
        rob_exception_1_1 = _RANDOM[11'h359][3];	// rob.scala:311:28
        rob_exception_1_2 = _RANDOM[11'h359][4];	// rob.scala:311:28
        rob_exception_1_3 = _RANDOM[11'h359][5];	// rob.scala:311:28
        rob_exception_1_4 = _RANDOM[11'h359][6];	// rob.scala:311:28
        rob_exception_1_5 = _RANDOM[11'h359][7];	// rob.scala:311:28
        rob_exception_1_6 = _RANDOM[11'h359][8];	// rob.scala:311:28
        rob_exception_1_7 = _RANDOM[11'h359][9];	// rob.scala:311:28
        rob_exception_1_8 = _RANDOM[11'h359][10];	// rob.scala:311:28
        rob_exception_1_9 = _RANDOM[11'h359][11];	// rob.scala:311:28
        rob_exception_1_10 = _RANDOM[11'h359][12];	// rob.scala:311:28
        rob_exception_1_11 = _RANDOM[11'h359][13];	// rob.scala:311:28
        rob_exception_1_12 = _RANDOM[11'h359][14];	// rob.scala:311:28
        rob_exception_1_13 = _RANDOM[11'h359][15];	// rob.scala:311:28
        rob_exception_1_14 = _RANDOM[11'h359][16];	// rob.scala:311:28
        rob_exception_1_15 = _RANDOM[11'h359][17];	// rob.scala:311:28
        rob_exception_1_16 = _RANDOM[11'h359][18];	// rob.scala:311:28
        rob_exception_1_17 = _RANDOM[11'h359][19];	// rob.scala:311:28
        rob_exception_1_18 = _RANDOM[11'h359][20];	// rob.scala:311:28
        rob_exception_1_19 = _RANDOM[11'h359][21];	// rob.scala:311:28
        rob_exception_1_20 = _RANDOM[11'h359][22];	// rob.scala:311:28
        rob_exception_1_21 = _RANDOM[11'h359][23];	// rob.scala:311:28
        rob_exception_1_22 = _RANDOM[11'h359][24];	// rob.scala:311:28
        rob_exception_1_23 = _RANDOM[11'h359][25];	// rob.scala:311:28
        rob_exception_1_24 = _RANDOM[11'h359][26];	// rob.scala:311:28
        rob_exception_1_25 = _RANDOM[11'h359][27];	// rob.scala:311:28
        rob_exception_1_26 = _RANDOM[11'h359][28];	// rob.scala:311:28
        rob_exception_1_27 = _RANDOM[11'h359][29];	// rob.scala:311:28
        rob_exception_1_28 = _RANDOM[11'h359][30];	// rob.scala:311:28
        rob_exception_1_29 = _RANDOM[11'h359][31];	// rob.scala:311:28
        rob_exception_1_30 = _RANDOM[11'h35A][0];	// rob.scala:311:28
        rob_exception_1_31 = _RANDOM[11'h35A][1];	// rob.scala:311:28
        rob_predicated_1_0 = _RANDOM[11'h35A][2];	// rob.scala:311:28, :312:29
        rob_predicated_1_1 = _RANDOM[11'h35A][3];	// rob.scala:311:28, :312:29
        rob_predicated_1_2 = _RANDOM[11'h35A][4];	// rob.scala:311:28, :312:29
        rob_predicated_1_3 = _RANDOM[11'h35A][5];	// rob.scala:311:28, :312:29
        rob_predicated_1_4 = _RANDOM[11'h35A][6];	// rob.scala:311:28, :312:29
        rob_predicated_1_5 = _RANDOM[11'h35A][7];	// rob.scala:311:28, :312:29
        rob_predicated_1_6 = _RANDOM[11'h35A][8];	// rob.scala:311:28, :312:29
        rob_predicated_1_7 = _RANDOM[11'h35A][9];	// rob.scala:311:28, :312:29
        rob_predicated_1_8 = _RANDOM[11'h35A][10];	// rob.scala:311:28, :312:29
        rob_predicated_1_9 = _RANDOM[11'h35A][11];	// rob.scala:311:28, :312:29
        rob_predicated_1_10 = _RANDOM[11'h35A][12];	// rob.scala:311:28, :312:29
        rob_predicated_1_11 = _RANDOM[11'h35A][13];	// rob.scala:311:28, :312:29
        rob_predicated_1_12 = _RANDOM[11'h35A][14];	// rob.scala:311:28, :312:29
        rob_predicated_1_13 = _RANDOM[11'h35A][15];	// rob.scala:311:28, :312:29
        rob_predicated_1_14 = _RANDOM[11'h35A][16];	// rob.scala:311:28, :312:29
        rob_predicated_1_15 = _RANDOM[11'h35A][17];	// rob.scala:311:28, :312:29
        rob_predicated_1_16 = _RANDOM[11'h35A][18];	// rob.scala:311:28, :312:29
        rob_predicated_1_17 = _RANDOM[11'h35A][19];	// rob.scala:311:28, :312:29
        rob_predicated_1_18 = _RANDOM[11'h35A][20];	// rob.scala:311:28, :312:29
        rob_predicated_1_19 = _RANDOM[11'h35A][21];	// rob.scala:311:28, :312:29
        rob_predicated_1_20 = _RANDOM[11'h35A][22];	// rob.scala:311:28, :312:29
        rob_predicated_1_21 = _RANDOM[11'h35A][23];	// rob.scala:311:28, :312:29
        rob_predicated_1_22 = _RANDOM[11'h35A][24];	// rob.scala:311:28, :312:29
        rob_predicated_1_23 = _RANDOM[11'h35A][25];	// rob.scala:311:28, :312:29
        rob_predicated_1_24 = _RANDOM[11'h35A][26];	// rob.scala:311:28, :312:29
        rob_predicated_1_25 = _RANDOM[11'h35A][27];	// rob.scala:311:28, :312:29
        rob_predicated_1_26 = _RANDOM[11'h35A][28];	// rob.scala:311:28, :312:29
        rob_predicated_1_27 = _RANDOM[11'h35A][29];	// rob.scala:311:28, :312:29
        rob_predicated_1_28 = _RANDOM[11'h35A][30];	// rob.scala:311:28, :312:29
        rob_predicated_1_29 = _RANDOM[11'h35A][31];	// rob.scala:311:28, :312:29
        rob_predicated_1_30 = _RANDOM[11'h35B][0];	// rob.scala:312:29
        rob_predicated_1_31 = _RANDOM[11'h35B][1];	// rob.scala:312:29
        rob_val_2_0 = _RANDOM[11'h35B][2];	// rob.scala:307:32, :312:29
        rob_val_2_1 = _RANDOM[11'h35B][3];	// rob.scala:307:32, :312:29
        rob_val_2_2 = _RANDOM[11'h35B][4];	// rob.scala:307:32, :312:29
        rob_val_2_3 = _RANDOM[11'h35B][5];	// rob.scala:307:32, :312:29
        rob_val_2_4 = _RANDOM[11'h35B][6];	// rob.scala:307:32, :312:29
        rob_val_2_5 = _RANDOM[11'h35B][7];	// rob.scala:307:32, :312:29
        rob_val_2_6 = _RANDOM[11'h35B][8];	// rob.scala:307:32, :312:29
        rob_val_2_7 = _RANDOM[11'h35B][9];	// rob.scala:307:32, :312:29
        rob_val_2_8 = _RANDOM[11'h35B][10];	// rob.scala:307:32, :312:29
        rob_val_2_9 = _RANDOM[11'h35B][11];	// rob.scala:307:32, :312:29
        rob_val_2_10 = _RANDOM[11'h35B][12];	// rob.scala:307:32, :312:29
        rob_val_2_11 = _RANDOM[11'h35B][13];	// rob.scala:307:32, :312:29
        rob_val_2_12 = _RANDOM[11'h35B][14];	// rob.scala:307:32, :312:29
        rob_val_2_13 = _RANDOM[11'h35B][15];	// rob.scala:307:32, :312:29
        rob_val_2_14 = _RANDOM[11'h35B][16];	// rob.scala:307:32, :312:29
        rob_val_2_15 = _RANDOM[11'h35B][17];	// rob.scala:307:32, :312:29
        rob_val_2_16 = _RANDOM[11'h35B][18];	// rob.scala:307:32, :312:29
        rob_val_2_17 = _RANDOM[11'h35B][19];	// rob.scala:307:32, :312:29
        rob_val_2_18 = _RANDOM[11'h35B][20];	// rob.scala:307:32, :312:29
        rob_val_2_19 = _RANDOM[11'h35B][21];	// rob.scala:307:32, :312:29
        rob_val_2_20 = _RANDOM[11'h35B][22];	// rob.scala:307:32, :312:29
        rob_val_2_21 = _RANDOM[11'h35B][23];	// rob.scala:307:32, :312:29
        rob_val_2_22 = _RANDOM[11'h35B][24];	// rob.scala:307:32, :312:29
        rob_val_2_23 = _RANDOM[11'h35B][25];	// rob.scala:307:32, :312:29
        rob_val_2_24 = _RANDOM[11'h35B][26];	// rob.scala:307:32, :312:29
        rob_val_2_25 = _RANDOM[11'h35B][27];	// rob.scala:307:32, :312:29
        rob_val_2_26 = _RANDOM[11'h35B][28];	// rob.scala:307:32, :312:29
        rob_val_2_27 = _RANDOM[11'h35B][29];	// rob.scala:307:32, :312:29
        rob_val_2_28 = _RANDOM[11'h35B][30];	// rob.scala:307:32, :312:29
        rob_val_2_29 = _RANDOM[11'h35B][31];	// rob.scala:307:32, :312:29
        rob_val_2_30 = _RANDOM[11'h35C][0];	// rob.scala:307:32
        rob_val_2_31 = _RANDOM[11'h35C][1];	// rob.scala:307:32
        rob_bsy_2_0 = _RANDOM[11'h35C][2];	// rob.scala:307:32, :308:28
        rob_bsy_2_1 = _RANDOM[11'h35C][3];	// rob.scala:307:32, :308:28
        rob_bsy_2_2 = _RANDOM[11'h35C][4];	// rob.scala:307:32, :308:28
        rob_bsy_2_3 = _RANDOM[11'h35C][5];	// rob.scala:307:32, :308:28
        rob_bsy_2_4 = _RANDOM[11'h35C][6];	// rob.scala:307:32, :308:28
        rob_bsy_2_5 = _RANDOM[11'h35C][7];	// rob.scala:307:32, :308:28
        rob_bsy_2_6 = _RANDOM[11'h35C][8];	// rob.scala:307:32, :308:28
        rob_bsy_2_7 = _RANDOM[11'h35C][9];	// rob.scala:307:32, :308:28
        rob_bsy_2_8 = _RANDOM[11'h35C][10];	// rob.scala:307:32, :308:28
        rob_bsy_2_9 = _RANDOM[11'h35C][11];	// rob.scala:307:32, :308:28
        rob_bsy_2_10 = _RANDOM[11'h35C][12];	// rob.scala:307:32, :308:28
        rob_bsy_2_11 = _RANDOM[11'h35C][13];	// rob.scala:307:32, :308:28
        rob_bsy_2_12 = _RANDOM[11'h35C][14];	// rob.scala:307:32, :308:28
        rob_bsy_2_13 = _RANDOM[11'h35C][15];	// rob.scala:307:32, :308:28
        rob_bsy_2_14 = _RANDOM[11'h35C][16];	// rob.scala:307:32, :308:28
        rob_bsy_2_15 = _RANDOM[11'h35C][17];	// rob.scala:307:32, :308:28
        rob_bsy_2_16 = _RANDOM[11'h35C][18];	// rob.scala:307:32, :308:28
        rob_bsy_2_17 = _RANDOM[11'h35C][19];	// rob.scala:307:32, :308:28
        rob_bsy_2_18 = _RANDOM[11'h35C][20];	// rob.scala:307:32, :308:28
        rob_bsy_2_19 = _RANDOM[11'h35C][21];	// rob.scala:307:32, :308:28
        rob_bsy_2_20 = _RANDOM[11'h35C][22];	// rob.scala:307:32, :308:28
        rob_bsy_2_21 = _RANDOM[11'h35C][23];	// rob.scala:307:32, :308:28
        rob_bsy_2_22 = _RANDOM[11'h35C][24];	// rob.scala:307:32, :308:28
        rob_bsy_2_23 = _RANDOM[11'h35C][25];	// rob.scala:307:32, :308:28
        rob_bsy_2_24 = _RANDOM[11'h35C][26];	// rob.scala:307:32, :308:28
        rob_bsy_2_25 = _RANDOM[11'h35C][27];	// rob.scala:307:32, :308:28
        rob_bsy_2_26 = _RANDOM[11'h35C][28];	// rob.scala:307:32, :308:28
        rob_bsy_2_27 = _RANDOM[11'h35C][29];	// rob.scala:307:32, :308:28
        rob_bsy_2_28 = _RANDOM[11'h35C][30];	// rob.scala:307:32, :308:28
        rob_bsy_2_29 = _RANDOM[11'h35C][31];	// rob.scala:307:32, :308:28
        rob_bsy_2_30 = _RANDOM[11'h35D][0];	// rob.scala:308:28
        rob_bsy_2_31 = _RANDOM[11'h35D][1];	// rob.scala:308:28
        rob_unsafe_2_0 = _RANDOM[11'h35D][2];	// rob.scala:308:28, :309:28
        rob_unsafe_2_1 = _RANDOM[11'h35D][3];	// rob.scala:308:28, :309:28
        rob_unsafe_2_2 = _RANDOM[11'h35D][4];	// rob.scala:308:28, :309:28
        rob_unsafe_2_3 = _RANDOM[11'h35D][5];	// rob.scala:308:28, :309:28
        rob_unsafe_2_4 = _RANDOM[11'h35D][6];	// rob.scala:308:28, :309:28
        rob_unsafe_2_5 = _RANDOM[11'h35D][7];	// rob.scala:308:28, :309:28
        rob_unsafe_2_6 = _RANDOM[11'h35D][8];	// rob.scala:308:28, :309:28
        rob_unsafe_2_7 = _RANDOM[11'h35D][9];	// rob.scala:308:28, :309:28
        rob_unsafe_2_8 = _RANDOM[11'h35D][10];	// rob.scala:308:28, :309:28
        rob_unsafe_2_9 = _RANDOM[11'h35D][11];	// rob.scala:308:28, :309:28
        rob_unsafe_2_10 = _RANDOM[11'h35D][12];	// rob.scala:308:28, :309:28
        rob_unsafe_2_11 = _RANDOM[11'h35D][13];	// rob.scala:308:28, :309:28
        rob_unsafe_2_12 = _RANDOM[11'h35D][14];	// rob.scala:308:28, :309:28
        rob_unsafe_2_13 = _RANDOM[11'h35D][15];	// rob.scala:308:28, :309:28
        rob_unsafe_2_14 = _RANDOM[11'h35D][16];	// rob.scala:308:28, :309:28
        rob_unsafe_2_15 = _RANDOM[11'h35D][17];	// rob.scala:308:28, :309:28
        rob_unsafe_2_16 = _RANDOM[11'h35D][18];	// rob.scala:308:28, :309:28
        rob_unsafe_2_17 = _RANDOM[11'h35D][19];	// rob.scala:308:28, :309:28
        rob_unsafe_2_18 = _RANDOM[11'h35D][20];	// rob.scala:308:28, :309:28
        rob_unsafe_2_19 = _RANDOM[11'h35D][21];	// rob.scala:308:28, :309:28
        rob_unsafe_2_20 = _RANDOM[11'h35D][22];	// rob.scala:308:28, :309:28
        rob_unsafe_2_21 = _RANDOM[11'h35D][23];	// rob.scala:308:28, :309:28
        rob_unsafe_2_22 = _RANDOM[11'h35D][24];	// rob.scala:308:28, :309:28
        rob_unsafe_2_23 = _RANDOM[11'h35D][25];	// rob.scala:308:28, :309:28
        rob_unsafe_2_24 = _RANDOM[11'h35D][26];	// rob.scala:308:28, :309:28
        rob_unsafe_2_25 = _RANDOM[11'h35D][27];	// rob.scala:308:28, :309:28
        rob_unsafe_2_26 = _RANDOM[11'h35D][28];	// rob.scala:308:28, :309:28
        rob_unsafe_2_27 = _RANDOM[11'h35D][29];	// rob.scala:308:28, :309:28
        rob_unsafe_2_28 = _RANDOM[11'h35D][30];	// rob.scala:308:28, :309:28
        rob_unsafe_2_29 = _RANDOM[11'h35D][31];	// rob.scala:308:28, :309:28
        rob_unsafe_2_30 = _RANDOM[11'h35E][0];	// rob.scala:309:28
        rob_unsafe_2_31 = _RANDOM[11'h35E][1];	// rob.scala:309:28
        rob_uop_2_0_uopc = _RANDOM[11'h35E][8:2];	// rob.scala:309:28, :310:28
        rob_uop_2_0_is_rvc = _RANDOM[11'h360][9];	// rob.scala:310:28
        rob_uop_2_0_br_mask = {_RANDOM[11'h362][31:30], _RANDOM[11'h363][17:0]};	// rob.scala:310:28
        rob_uop_2_0_ftq_idx = _RANDOM[11'h363][28:23];	// rob.scala:310:28
        rob_uop_2_0_edge_inst = _RANDOM[11'h363][29];	// rob.scala:310:28
        rob_uop_2_0_pc_lob = {_RANDOM[11'h363][31:30], _RANDOM[11'h364][3:0]};	// rob.scala:310:28
        rob_uop_2_0_pdst = _RANDOM[11'h365][30:24];	// rob.scala:310:28
        rob_uop_2_0_stale_pdst = {_RANDOM[11'h366][31:30], _RANDOM[11'h367][4:0]};	// rob.scala:310:28
        rob_uop_2_0_is_fencei = _RANDOM[11'h369][16];	// rob.scala:310:28
        rob_uop_2_0_uses_ldq = _RANDOM[11'h369][18];	// rob.scala:310:28
        rob_uop_2_0_uses_stq = _RANDOM[11'h369][19];	// rob.scala:310:28
        rob_uop_2_0_is_sys_pc2epc = _RANDOM[11'h369][20];	// rob.scala:310:28
        rob_uop_2_0_flush_on_commit = _RANDOM[11'h369][22];	// rob.scala:310:28
        rob_uop_2_0_ldst = _RANDOM[11'h369][29:24];	// rob.scala:310:28
        rob_uop_2_0_ldst_val = _RANDOM[11'h36A][16];	// rob.scala:310:28
        rob_uop_2_0_dst_rtype = _RANDOM[11'h36A][18:17];	// rob.scala:310:28
        rob_uop_2_0_fp_val = _RANDOM[11'h36A][24];	// rob.scala:310:28
        rob_uop_2_1_uopc = _RANDOM[11'h36B][9:3];	// rob.scala:310:28
        rob_uop_2_1_is_rvc = _RANDOM[11'h36D][10];	// rob.scala:310:28
        rob_uop_2_1_br_mask = {_RANDOM[11'h36F][31], _RANDOM[11'h370][18:0]};	// rob.scala:310:28
        rob_uop_2_1_ftq_idx = _RANDOM[11'h370][29:24];	// rob.scala:310:28
        rob_uop_2_1_edge_inst = _RANDOM[11'h370][30];	// rob.scala:310:28
        rob_uop_2_1_pc_lob = {_RANDOM[11'h370][31], _RANDOM[11'h371][4:0]};	// rob.scala:310:28
        rob_uop_2_1_pdst = _RANDOM[11'h372][31:25];	// rob.scala:310:28
        rob_uop_2_1_stale_pdst = {_RANDOM[11'h373][31], _RANDOM[11'h374][5:0]};	// rob.scala:310:28
        rob_uop_2_1_is_fencei = _RANDOM[11'h376][17];	// rob.scala:310:28
        rob_uop_2_1_uses_ldq = _RANDOM[11'h376][19];	// rob.scala:310:28
        rob_uop_2_1_uses_stq = _RANDOM[11'h376][20];	// rob.scala:310:28
        rob_uop_2_1_is_sys_pc2epc = _RANDOM[11'h376][21];	// rob.scala:310:28
        rob_uop_2_1_flush_on_commit = _RANDOM[11'h376][23];	// rob.scala:310:28
        rob_uop_2_1_ldst = _RANDOM[11'h376][30:25];	// rob.scala:310:28
        rob_uop_2_1_ldst_val = _RANDOM[11'h377][17];	// rob.scala:310:28
        rob_uop_2_1_dst_rtype = _RANDOM[11'h377][19:18];	// rob.scala:310:28
        rob_uop_2_1_fp_val = _RANDOM[11'h377][25];	// rob.scala:310:28
        rob_uop_2_2_uopc = _RANDOM[11'h378][10:4];	// rob.scala:310:28
        rob_uop_2_2_is_rvc = _RANDOM[11'h37A][11];	// rob.scala:310:28
        rob_uop_2_2_br_mask = _RANDOM[11'h37D][19:0];	// rob.scala:310:28
        rob_uop_2_2_ftq_idx = _RANDOM[11'h37D][30:25];	// rob.scala:310:28
        rob_uop_2_2_edge_inst = _RANDOM[11'h37D][31];	// rob.scala:310:28
        rob_uop_2_2_pc_lob = _RANDOM[11'h37E][5:0];	// rob.scala:310:28
        rob_uop_2_2_pdst = {_RANDOM[11'h37F][31:26], _RANDOM[11'h380][0]};	// rob.scala:310:28
        rob_uop_2_2_stale_pdst = _RANDOM[11'h381][6:0];	// rob.scala:310:28
        rob_uop_2_2_is_fencei = _RANDOM[11'h383][18];	// rob.scala:310:28
        rob_uop_2_2_uses_ldq = _RANDOM[11'h383][20];	// rob.scala:310:28
        rob_uop_2_2_uses_stq = _RANDOM[11'h383][21];	// rob.scala:310:28
        rob_uop_2_2_is_sys_pc2epc = _RANDOM[11'h383][22];	// rob.scala:310:28
        rob_uop_2_2_flush_on_commit = _RANDOM[11'h383][24];	// rob.scala:310:28
        rob_uop_2_2_ldst = _RANDOM[11'h383][31:26];	// rob.scala:310:28
        rob_uop_2_2_ldst_val = _RANDOM[11'h384][18];	// rob.scala:310:28
        rob_uop_2_2_dst_rtype = _RANDOM[11'h384][20:19];	// rob.scala:310:28
        rob_uop_2_2_fp_val = _RANDOM[11'h384][26];	// rob.scala:310:28
        rob_uop_2_3_uopc = _RANDOM[11'h385][11:5];	// rob.scala:310:28
        rob_uop_2_3_is_rvc = _RANDOM[11'h387][12];	// rob.scala:310:28
        rob_uop_2_3_br_mask = _RANDOM[11'h38A][20:1];	// rob.scala:310:28
        rob_uop_2_3_ftq_idx = _RANDOM[11'h38A][31:26];	// rob.scala:310:28
        rob_uop_2_3_edge_inst = _RANDOM[11'h38B][0];	// rob.scala:310:28
        rob_uop_2_3_pc_lob = _RANDOM[11'h38B][6:1];	// rob.scala:310:28
        rob_uop_2_3_pdst = {_RANDOM[11'h38C][31:27], _RANDOM[11'h38D][1:0]};	// rob.scala:310:28
        rob_uop_2_3_stale_pdst = _RANDOM[11'h38E][7:1];	// rob.scala:310:28
        rob_uop_2_3_is_fencei = _RANDOM[11'h390][19];	// rob.scala:310:28
        rob_uop_2_3_uses_ldq = _RANDOM[11'h390][21];	// rob.scala:310:28
        rob_uop_2_3_uses_stq = _RANDOM[11'h390][22];	// rob.scala:310:28
        rob_uop_2_3_is_sys_pc2epc = _RANDOM[11'h390][23];	// rob.scala:310:28
        rob_uop_2_3_flush_on_commit = _RANDOM[11'h390][25];	// rob.scala:310:28
        rob_uop_2_3_ldst = {_RANDOM[11'h390][31:27], _RANDOM[11'h391][0]};	// rob.scala:310:28
        rob_uop_2_3_ldst_val = _RANDOM[11'h391][19];	// rob.scala:310:28
        rob_uop_2_3_dst_rtype = _RANDOM[11'h391][21:20];	// rob.scala:310:28
        rob_uop_2_3_fp_val = _RANDOM[11'h391][27];	// rob.scala:310:28
        rob_uop_2_4_uopc = _RANDOM[11'h392][12:6];	// rob.scala:310:28
        rob_uop_2_4_is_rvc = _RANDOM[11'h394][13];	// rob.scala:310:28
        rob_uop_2_4_br_mask = _RANDOM[11'h397][21:2];	// rob.scala:310:28
        rob_uop_2_4_ftq_idx = {_RANDOM[11'h397][31:27], _RANDOM[11'h398][0]};	// rob.scala:310:28
        rob_uop_2_4_edge_inst = _RANDOM[11'h398][1];	// rob.scala:310:28
        rob_uop_2_4_pc_lob = _RANDOM[11'h398][7:2];	// rob.scala:310:28
        rob_uop_2_4_pdst = {_RANDOM[11'h399][31:28], _RANDOM[11'h39A][2:0]};	// rob.scala:310:28
        rob_uop_2_4_stale_pdst = _RANDOM[11'h39B][8:2];	// rob.scala:310:28
        rob_uop_2_4_is_fencei = _RANDOM[11'h39D][20];	// rob.scala:310:28
        rob_uop_2_4_uses_ldq = _RANDOM[11'h39D][22];	// rob.scala:310:28
        rob_uop_2_4_uses_stq = _RANDOM[11'h39D][23];	// rob.scala:310:28
        rob_uop_2_4_is_sys_pc2epc = _RANDOM[11'h39D][24];	// rob.scala:310:28
        rob_uop_2_4_flush_on_commit = _RANDOM[11'h39D][26];	// rob.scala:310:28
        rob_uop_2_4_ldst = {_RANDOM[11'h39D][31:28], _RANDOM[11'h39E][1:0]};	// rob.scala:310:28
        rob_uop_2_4_ldst_val = _RANDOM[11'h39E][20];	// rob.scala:310:28
        rob_uop_2_4_dst_rtype = _RANDOM[11'h39E][22:21];	// rob.scala:310:28
        rob_uop_2_4_fp_val = _RANDOM[11'h39E][28];	// rob.scala:310:28
        rob_uop_2_5_uopc = _RANDOM[11'h39F][13:7];	// rob.scala:310:28
        rob_uop_2_5_is_rvc = _RANDOM[11'h3A1][14];	// rob.scala:310:28
        rob_uop_2_5_br_mask = _RANDOM[11'h3A4][22:3];	// rob.scala:310:28
        rob_uop_2_5_ftq_idx = {_RANDOM[11'h3A4][31:28], _RANDOM[11'h3A5][1:0]};	// rob.scala:310:28
        rob_uop_2_5_edge_inst = _RANDOM[11'h3A5][2];	// rob.scala:310:28
        rob_uop_2_5_pc_lob = _RANDOM[11'h3A5][8:3];	// rob.scala:310:28
        rob_uop_2_5_pdst = {_RANDOM[11'h3A6][31:29], _RANDOM[11'h3A7][3:0]};	// rob.scala:310:28
        rob_uop_2_5_stale_pdst = _RANDOM[11'h3A8][9:3];	// rob.scala:310:28
        rob_uop_2_5_is_fencei = _RANDOM[11'h3AA][21];	// rob.scala:310:28
        rob_uop_2_5_uses_ldq = _RANDOM[11'h3AA][23];	// rob.scala:310:28
        rob_uop_2_5_uses_stq = _RANDOM[11'h3AA][24];	// rob.scala:310:28
        rob_uop_2_5_is_sys_pc2epc = _RANDOM[11'h3AA][25];	// rob.scala:310:28
        rob_uop_2_5_flush_on_commit = _RANDOM[11'h3AA][27];	// rob.scala:310:28
        rob_uop_2_5_ldst = {_RANDOM[11'h3AA][31:29], _RANDOM[11'h3AB][2:0]};	// rob.scala:310:28
        rob_uop_2_5_ldst_val = _RANDOM[11'h3AB][21];	// rob.scala:310:28
        rob_uop_2_5_dst_rtype = _RANDOM[11'h3AB][23:22];	// rob.scala:310:28
        rob_uop_2_5_fp_val = _RANDOM[11'h3AB][29];	// rob.scala:310:28
        rob_uop_2_6_uopc = _RANDOM[11'h3AC][14:8];	// rob.scala:310:28
        rob_uop_2_6_is_rvc = _RANDOM[11'h3AE][15];	// rob.scala:310:28
        rob_uop_2_6_br_mask = _RANDOM[11'h3B1][23:4];	// rob.scala:310:28
        rob_uop_2_6_ftq_idx = {_RANDOM[11'h3B1][31:29], _RANDOM[11'h3B2][2:0]};	// rob.scala:310:28
        rob_uop_2_6_edge_inst = _RANDOM[11'h3B2][3];	// rob.scala:310:28
        rob_uop_2_6_pc_lob = _RANDOM[11'h3B2][9:4];	// rob.scala:310:28
        rob_uop_2_6_pdst = {_RANDOM[11'h3B3][31:30], _RANDOM[11'h3B4][4:0]};	// rob.scala:310:28
        rob_uop_2_6_stale_pdst = _RANDOM[11'h3B5][10:4];	// rob.scala:310:28
        rob_uop_2_6_is_fencei = _RANDOM[11'h3B7][22];	// rob.scala:310:28
        rob_uop_2_6_uses_ldq = _RANDOM[11'h3B7][24];	// rob.scala:310:28
        rob_uop_2_6_uses_stq = _RANDOM[11'h3B7][25];	// rob.scala:310:28
        rob_uop_2_6_is_sys_pc2epc = _RANDOM[11'h3B7][26];	// rob.scala:310:28
        rob_uop_2_6_flush_on_commit = _RANDOM[11'h3B7][28];	// rob.scala:310:28
        rob_uop_2_6_ldst = {_RANDOM[11'h3B7][31:30], _RANDOM[11'h3B8][3:0]};	// rob.scala:310:28
        rob_uop_2_6_ldst_val = _RANDOM[11'h3B8][22];	// rob.scala:310:28
        rob_uop_2_6_dst_rtype = _RANDOM[11'h3B8][24:23];	// rob.scala:310:28
        rob_uop_2_6_fp_val = _RANDOM[11'h3B8][30];	// rob.scala:310:28
        rob_uop_2_7_uopc = _RANDOM[11'h3B9][15:9];	// rob.scala:310:28
        rob_uop_2_7_is_rvc = _RANDOM[11'h3BB][16];	// rob.scala:310:28
        rob_uop_2_7_br_mask = _RANDOM[11'h3BE][24:5];	// rob.scala:310:28
        rob_uop_2_7_ftq_idx = {_RANDOM[11'h3BE][31:30], _RANDOM[11'h3BF][3:0]};	// rob.scala:310:28
        rob_uop_2_7_edge_inst = _RANDOM[11'h3BF][4];	// rob.scala:310:28
        rob_uop_2_7_pc_lob = _RANDOM[11'h3BF][10:5];	// rob.scala:310:28
        rob_uop_2_7_pdst = {_RANDOM[11'h3C0][31], _RANDOM[11'h3C1][5:0]};	// rob.scala:310:28
        rob_uop_2_7_stale_pdst = _RANDOM[11'h3C2][11:5];	// rob.scala:310:28
        rob_uop_2_7_is_fencei = _RANDOM[11'h3C4][23];	// rob.scala:310:28
        rob_uop_2_7_uses_ldq = _RANDOM[11'h3C4][25];	// rob.scala:310:28
        rob_uop_2_7_uses_stq = _RANDOM[11'h3C4][26];	// rob.scala:310:28
        rob_uop_2_7_is_sys_pc2epc = _RANDOM[11'h3C4][27];	// rob.scala:310:28
        rob_uop_2_7_flush_on_commit = _RANDOM[11'h3C4][29];	// rob.scala:310:28
        rob_uop_2_7_ldst = {_RANDOM[11'h3C4][31], _RANDOM[11'h3C5][4:0]};	// rob.scala:310:28
        rob_uop_2_7_ldst_val = _RANDOM[11'h3C5][23];	// rob.scala:310:28
        rob_uop_2_7_dst_rtype = _RANDOM[11'h3C5][25:24];	// rob.scala:310:28
        rob_uop_2_7_fp_val = _RANDOM[11'h3C5][31];	// rob.scala:310:28
        rob_uop_2_8_uopc = _RANDOM[11'h3C6][16:10];	// rob.scala:310:28
        rob_uop_2_8_is_rvc = _RANDOM[11'h3C8][17];	// rob.scala:310:28
        rob_uop_2_8_br_mask = _RANDOM[11'h3CB][25:6];	// rob.scala:310:28
        rob_uop_2_8_ftq_idx = {_RANDOM[11'h3CB][31], _RANDOM[11'h3CC][4:0]};	// rob.scala:310:28
        rob_uop_2_8_edge_inst = _RANDOM[11'h3CC][5];	// rob.scala:310:28
        rob_uop_2_8_pc_lob = _RANDOM[11'h3CC][11:6];	// rob.scala:310:28
        rob_uop_2_8_pdst = _RANDOM[11'h3CE][6:0];	// rob.scala:310:28
        rob_uop_2_8_stale_pdst = _RANDOM[11'h3CF][12:6];	// rob.scala:310:28
        rob_uop_2_8_is_fencei = _RANDOM[11'h3D1][24];	// rob.scala:310:28
        rob_uop_2_8_uses_ldq = _RANDOM[11'h3D1][26];	// rob.scala:310:28
        rob_uop_2_8_uses_stq = _RANDOM[11'h3D1][27];	// rob.scala:310:28
        rob_uop_2_8_is_sys_pc2epc = _RANDOM[11'h3D1][28];	// rob.scala:310:28
        rob_uop_2_8_flush_on_commit = _RANDOM[11'h3D1][30];	// rob.scala:310:28
        rob_uop_2_8_ldst = _RANDOM[11'h3D2][5:0];	// rob.scala:310:28
        rob_uop_2_8_ldst_val = _RANDOM[11'h3D2][24];	// rob.scala:310:28
        rob_uop_2_8_dst_rtype = _RANDOM[11'h3D2][26:25];	// rob.scala:310:28
        rob_uop_2_8_fp_val = _RANDOM[11'h3D3][0];	// rob.scala:310:28
        rob_uop_2_9_uopc = _RANDOM[11'h3D3][17:11];	// rob.scala:310:28
        rob_uop_2_9_is_rvc = _RANDOM[11'h3D5][18];	// rob.scala:310:28
        rob_uop_2_9_br_mask = _RANDOM[11'h3D8][26:7];	// rob.scala:310:28
        rob_uop_2_9_ftq_idx = _RANDOM[11'h3D9][5:0];	// rob.scala:310:28
        rob_uop_2_9_edge_inst = _RANDOM[11'h3D9][6];	// rob.scala:310:28
        rob_uop_2_9_pc_lob = _RANDOM[11'h3D9][12:7];	// rob.scala:310:28
        rob_uop_2_9_pdst = _RANDOM[11'h3DB][7:1];	// rob.scala:310:28
        rob_uop_2_9_stale_pdst = _RANDOM[11'h3DC][13:7];	// rob.scala:310:28
        rob_uop_2_9_is_fencei = _RANDOM[11'h3DE][25];	// rob.scala:310:28
        rob_uop_2_9_uses_ldq = _RANDOM[11'h3DE][27];	// rob.scala:310:28
        rob_uop_2_9_uses_stq = _RANDOM[11'h3DE][28];	// rob.scala:310:28
        rob_uop_2_9_is_sys_pc2epc = _RANDOM[11'h3DE][29];	// rob.scala:310:28
        rob_uop_2_9_flush_on_commit = _RANDOM[11'h3DE][31];	// rob.scala:310:28
        rob_uop_2_9_ldst = _RANDOM[11'h3DF][6:1];	// rob.scala:310:28
        rob_uop_2_9_ldst_val = _RANDOM[11'h3DF][25];	// rob.scala:310:28
        rob_uop_2_9_dst_rtype = _RANDOM[11'h3DF][27:26];	// rob.scala:310:28
        rob_uop_2_9_fp_val = _RANDOM[11'h3E0][1];	// rob.scala:310:28
        rob_uop_2_10_uopc = _RANDOM[11'h3E0][18:12];	// rob.scala:310:28
        rob_uop_2_10_is_rvc = _RANDOM[11'h3E2][19];	// rob.scala:310:28
        rob_uop_2_10_br_mask = _RANDOM[11'h3E5][27:8];	// rob.scala:310:28
        rob_uop_2_10_ftq_idx = _RANDOM[11'h3E6][6:1];	// rob.scala:310:28
        rob_uop_2_10_edge_inst = _RANDOM[11'h3E6][7];	// rob.scala:310:28
        rob_uop_2_10_pc_lob = _RANDOM[11'h3E6][13:8];	// rob.scala:310:28
        rob_uop_2_10_pdst = _RANDOM[11'h3E8][8:2];	// rob.scala:310:28
        rob_uop_2_10_stale_pdst = _RANDOM[11'h3E9][14:8];	// rob.scala:310:28
        rob_uop_2_10_is_fencei = _RANDOM[11'h3EB][26];	// rob.scala:310:28
        rob_uop_2_10_uses_ldq = _RANDOM[11'h3EB][28];	// rob.scala:310:28
        rob_uop_2_10_uses_stq = _RANDOM[11'h3EB][29];	// rob.scala:310:28
        rob_uop_2_10_is_sys_pc2epc = _RANDOM[11'h3EB][30];	// rob.scala:310:28
        rob_uop_2_10_flush_on_commit = _RANDOM[11'h3EC][0];	// rob.scala:310:28
        rob_uop_2_10_ldst = _RANDOM[11'h3EC][7:2];	// rob.scala:310:28
        rob_uop_2_10_ldst_val = _RANDOM[11'h3EC][26];	// rob.scala:310:28
        rob_uop_2_10_dst_rtype = _RANDOM[11'h3EC][28:27];	// rob.scala:310:28
        rob_uop_2_10_fp_val = _RANDOM[11'h3ED][2];	// rob.scala:310:28
        rob_uop_2_11_uopc = _RANDOM[11'h3ED][19:13];	// rob.scala:310:28
        rob_uop_2_11_is_rvc = _RANDOM[11'h3EF][20];	// rob.scala:310:28
        rob_uop_2_11_br_mask = _RANDOM[11'h3F2][28:9];	// rob.scala:310:28
        rob_uop_2_11_ftq_idx = _RANDOM[11'h3F3][7:2];	// rob.scala:310:28
        rob_uop_2_11_edge_inst = _RANDOM[11'h3F3][8];	// rob.scala:310:28
        rob_uop_2_11_pc_lob = _RANDOM[11'h3F3][14:9];	// rob.scala:310:28
        rob_uop_2_11_pdst = _RANDOM[11'h3F5][9:3];	// rob.scala:310:28
        rob_uop_2_11_stale_pdst = _RANDOM[11'h3F6][15:9];	// rob.scala:310:28
        rob_uop_2_11_is_fencei = _RANDOM[11'h3F8][27];	// rob.scala:310:28
        rob_uop_2_11_uses_ldq = _RANDOM[11'h3F8][29];	// rob.scala:310:28
        rob_uop_2_11_uses_stq = _RANDOM[11'h3F8][30];	// rob.scala:310:28
        rob_uop_2_11_is_sys_pc2epc = _RANDOM[11'h3F8][31];	// rob.scala:310:28
        rob_uop_2_11_flush_on_commit = _RANDOM[11'h3F9][1];	// rob.scala:310:28
        rob_uop_2_11_ldst = _RANDOM[11'h3F9][8:3];	// rob.scala:310:28
        rob_uop_2_11_ldst_val = _RANDOM[11'h3F9][27];	// rob.scala:310:28
        rob_uop_2_11_dst_rtype = _RANDOM[11'h3F9][29:28];	// rob.scala:310:28
        rob_uop_2_11_fp_val = _RANDOM[11'h3FA][3];	// rob.scala:310:28
        rob_uop_2_12_uopc = _RANDOM[11'h3FA][20:14];	// rob.scala:310:28
        rob_uop_2_12_is_rvc = _RANDOM[11'h3FC][21];	// rob.scala:310:28
        rob_uop_2_12_br_mask = _RANDOM[11'h3FF][29:10];	// rob.scala:310:28
        rob_uop_2_12_ftq_idx = _RANDOM[11'h400][8:3];	// rob.scala:310:28
        rob_uop_2_12_edge_inst = _RANDOM[11'h400][9];	// rob.scala:310:28
        rob_uop_2_12_pc_lob = _RANDOM[11'h400][15:10];	// rob.scala:310:28
        rob_uop_2_12_pdst = _RANDOM[11'h402][10:4];	// rob.scala:310:28
        rob_uop_2_12_stale_pdst = _RANDOM[11'h403][16:10];	// rob.scala:310:28
        rob_uop_2_12_is_fencei = _RANDOM[11'h405][28];	// rob.scala:310:28
        rob_uop_2_12_uses_ldq = _RANDOM[11'h405][30];	// rob.scala:310:28
        rob_uop_2_12_uses_stq = _RANDOM[11'h405][31];	// rob.scala:310:28
        rob_uop_2_12_is_sys_pc2epc = _RANDOM[11'h406][0];	// rob.scala:310:28
        rob_uop_2_12_flush_on_commit = _RANDOM[11'h406][2];	// rob.scala:310:28
        rob_uop_2_12_ldst = _RANDOM[11'h406][9:4];	// rob.scala:310:28
        rob_uop_2_12_ldst_val = _RANDOM[11'h406][28];	// rob.scala:310:28
        rob_uop_2_12_dst_rtype = _RANDOM[11'h406][30:29];	// rob.scala:310:28
        rob_uop_2_12_fp_val = _RANDOM[11'h407][4];	// rob.scala:310:28
        rob_uop_2_13_uopc = _RANDOM[11'h407][21:15];	// rob.scala:310:28
        rob_uop_2_13_is_rvc = _RANDOM[11'h409][22];	// rob.scala:310:28
        rob_uop_2_13_br_mask = _RANDOM[11'h40C][30:11];	// rob.scala:310:28
        rob_uop_2_13_ftq_idx = _RANDOM[11'h40D][9:4];	// rob.scala:310:28
        rob_uop_2_13_edge_inst = _RANDOM[11'h40D][10];	// rob.scala:310:28
        rob_uop_2_13_pc_lob = _RANDOM[11'h40D][16:11];	// rob.scala:310:28
        rob_uop_2_13_pdst = _RANDOM[11'h40F][11:5];	// rob.scala:310:28
        rob_uop_2_13_stale_pdst = _RANDOM[11'h410][17:11];	// rob.scala:310:28
        rob_uop_2_13_is_fencei = _RANDOM[11'h412][29];	// rob.scala:310:28
        rob_uop_2_13_uses_ldq = _RANDOM[11'h412][31];	// rob.scala:310:28
        rob_uop_2_13_uses_stq = _RANDOM[11'h413][0];	// rob.scala:310:28
        rob_uop_2_13_is_sys_pc2epc = _RANDOM[11'h413][1];	// rob.scala:310:28
        rob_uop_2_13_flush_on_commit = _RANDOM[11'h413][3];	// rob.scala:310:28
        rob_uop_2_13_ldst = _RANDOM[11'h413][10:5];	// rob.scala:310:28
        rob_uop_2_13_ldst_val = _RANDOM[11'h413][29];	// rob.scala:310:28
        rob_uop_2_13_dst_rtype = _RANDOM[11'h413][31:30];	// rob.scala:310:28
        rob_uop_2_13_fp_val = _RANDOM[11'h414][5];	// rob.scala:310:28
        rob_uop_2_14_uopc = _RANDOM[11'h414][22:16];	// rob.scala:310:28
        rob_uop_2_14_is_rvc = _RANDOM[11'h416][23];	// rob.scala:310:28
        rob_uop_2_14_br_mask = _RANDOM[11'h419][31:12];	// rob.scala:310:28
        rob_uop_2_14_ftq_idx = _RANDOM[11'h41A][10:5];	// rob.scala:310:28
        rob_uop_2_14_edge_inst = _RANDOM[11'h41A][11];	// rob.scala:310:28
        rob_uop_2_14_pc_lob = _RANDOM[11'h41A][17:12];	// rob.scala:310:28
        rob_uop_2_14_pdst = _RANDOM[11'h41C][12:6];	// rob.scala:310:28
        rob_uop_2_14_stale_pdst = _RANDOM[11'h41D][18:12];	// rob.scala:310:28
        rob_uop_2_14_is_fencei = _RANDOM[11'h41F][30];	// rob.scala:310:28
        rob_uop_2_14_uses_ldq = _RANDOM[11'h420][0];	// rob.scala:310:28
        rob_uop_2_14_uses_stq = _RANDOM[11'h420][1];	// rob.scala:310:28
        rob_uop_2_14_is_sys_pc2epc = _RANDOM[11'h420][2];	// rob.scala:310:28
        rob_uop_2_14_flush_on_commit = _RANDOM[11'h420][4];	// rob.scala:310:28
        rob_uop_2_14_ldst = _RANDOM[11'h420][11:6];	// rob.scala:310:28
        rob_uop_2_14_ldst_val = _RANDOM[11'h420][30];	// rob.scala:310:28
        rob_uop_2_14_dst_rtype = {_RANDOM[11'h420][31], _RANDOM[11'h421][0]};	// rob.scala:310:28
        rob_uop_2_14_fp_val = _RANDOM[11'h421][6];	// rob.scala:310:28
        rob_uop_2_15_uopc = _RANDOM[11'h421][23:17];	// rob.scala:310:28
        rob_uop_2_15_is_rvc = _RANDOM[11'h423][24];	// rob.scala:310:28
        rob_uop_2_15_br_mask = {_RANDOM[11'h426][31:13], _RANDOM[11'h427][0]};	// rob.scala:310:28
        rob_uop_2_15_ftq_idx = _RANDOM[11'h427][11:6];	// rob.scala:310:28
        rob_uop_2_15_edge_inst = _RANDOM[11'h427][12];	// rob.scala:310:28
        rob_uop_2_15_pc_lob = _RANDOM[11'h427][18:13];	// rob.scala:310:28
        rob_uop_2_15_pdst = _RANDOM[11'h429][13:7];	// rob.scala:310:28
        rob_uop_2_15_stale_pdst = _RANDOM[11'h42A][19:13];	// rob.scala:310:28
        rob_uop_2_15_is_fencei = _RANDOM[11'h42C][31];	// rob.scala:310:28
        rob_uop_2_15_uses_ldq = _RANDOM[11'h42D][1];	// rob.scala:310:28
        rob_uop_2_15_uses_stq = _RANDOM[11'h42D][2];	// rob.scala:310:28
        rob_uop_2_15_is_sys_pc2epc = _RANDOM[11'h42D][3];	// rob.scala:310:28
        rob_uop_2_15_flush_on_commit = _RANDOM[11'h42D][5];	// rob.scala:310:28
        rob_uop_2_15_ldst = _RANDOM[11'h42D][12:7];	// rob.scala:310:28
        rob_uop_2_15_ldst_val = _RANDOM[11'h42D][31];	// rob.scala:310:28
        rob_uop_2_15_dst_rtype = _RANDOM[11'h42E][1:0];	// rob.scala:310:28
        rob_uop_2_15_fp_val = _RANDOM[11'h42E][7];	// rob.scala:310:28
        rob_uop_2_16_uopc = _RANDOM[11'h42E][24:18];	// rob.scala:310:28
        rob_uop_2_16_is_rvc = _RANDOM[11'h430][25];	// rob.scala:310:28
        rob_uop_2_16_br_mask = {_RANDOM[11'h433][31:14], _RANDOM[11'h434][1:0]};	// rob.scala:310:28
        rob_uop_2_16_ftq_idx = _RANDOM[11'h434][12:7];	// rob.scala:310:28
        rob_uop_2_16_edge_inst = _RANDOM[11'h434][13];	// rob.scala:310:28
        rob_uop_2_16_pc_lob = _RANDOM[11'h434][19:14];	// rob.scala:310:28
        rob_uop_2_16_pdst = _RANDOM[11'h436][14:8];	// rob.scala:310:28
        rob_uop_2_16_stale_pdst = _RANDOM[11'h437][20:14];	// rob.scala:310:28
        rob_uop_2_16_is_fencei = _RANDOM[11'h43A][0];	// rob.scala:310:28
        rob_uop_2_16_uses_ldq = _RANDOM[11'h43A][2];	// rob.scala:310:28
        rob_uop_2_16_uses_stq = _RANDOM[11'h43A][3];	// rob.scala:310:28
        rob_uop_2_16_is_sys_pc2epc = _RANDOM[11'h43A][4];	// rob.scala:310:28
        rob_uop_2_16_flush_on_commit = _RANDOM[11'h43A][6];	// rob.scala:310:28
        rob_uop_2_16_ldst = _RANDOM[11'h43A][13:8];	// rob.scala:310:28
        rob_uop_2_16_ldst_val = _RANDOM[11'h43B][0];	// rob.scala:310:28
        rob_uop_2_16_dst_rtype = _RANDOM[11'h43B][2:1];	// rob.scala:310:28
        rob_uop_2_16_fp_val = _RANDOM[11'h43B][8];	// rob.scala:310:28
        rob_uop_2_17_uopc = _RANDOM[11'h43B][25:19];	// rob.scala:310:28
        rob_uop_2_17_is_rvc = _RANDOM[11'h43D][26];	// rob.scala:310:28
        rob_uop_2_17_br_mask = {_RANDOM[11'h440][31:15], _RANDOM[11'h441][2:0]};	// rob.scala:310:28
        rob_uop_2_17_ftq_idx = _RANDOM[11'h441][13:8];	// rob.scala:310:28
        rob_uop_2_17_edge_inst = _RANDOM[11'h441][14];	// rob.scala:310:28
        rob_uop_2_17_pc_lob = _RANDOM[11'h441][20:15];	// rob.scala:310:28
        rob_uop_2_17_pdst = _RANDOM[11'h443][15:9];	// rob.scala:310:28
        rob_uop_2_17_stale_pdst = _RANDOM[11'h444][21:15];	// rob.scala:310:28
        rob_uop_2_17_is_fencei = _RANDOM[11'h447][1];	// rob.scala:310:28
        rob_uop_2_17_uses_ldq = _RANDOM[11'h447][3];	// rob.scala:310:28
        rob_uop_2_17_uses_stq = _RANDOM[11'h447][4];	// rob.scala:310:28
        rob_uop_2_17_is_sys_pc2epc = _RANDOM[11'h447][5];	// rob.scala:310:28
        rob_uop_2_17_flush_on_commit = _RANDOM[11'h447][7];	// rob.scala:310:28
        rob_uop_2_17_ldst = _RANDOM[11'h447][14:9];	// rob.scala:310:28
        rob_uop_2_17_ldst_val = _RANDOM[11'h448][1];	// rob.scala:310:28
        rob_uop_2_17_dst_rtype = _RANDOM[11'h448][3:2];	// rob.scala:310:28
        rob_uop_2_17_fp_val = _RANDOM[11'h448][9];	// rob.scala:310:28
        rob_uop_2_18_uopc = _RANDOM[11'h448][26:20];	// rob.scala:310:28
        rob_uop_2_18_is_rvc = _RANDOM[11'h44A][27];	// rob.scala:310:28
        rob_uop_2_18_br_mask = {_RANDOM[11'h44D][31:16], _RANDOM[11'h44E][3:0]};	// rob.scala:310:28
        rob_uop_2_18_ftq_idx = _RANDOM[11'h44E][14:9];	// rob.scala:310:28
        rob_uop_2_18_edge_inst = _RANDOM[11'h44E][15];	// rob.scala:310:28
        rob_uop_2_18_pc_lob = _RANDOM[11'h44E][21:16];	// rob.scala:310:28
        rob_uop_2_18_pdst = _RANDOM[11'h450][16:10];	// rob.scala:310:28
        rob_uop_2_18_stale_pdst = _RANDOM[11'h451][22:16];	// rob.scala:310:28
        rob_uop_2_18_is_fencei = _RANDOM[11'h454][2];	// rob.scala:310:28
        rob_uop_2_18_uses_ldq = _RANDOM[11'h454][4];	// rob.scala:310:28
        rob_uop_2_18_uses_stq = _RANDOM[11'h454][5];	// rob.scala:310:28
        rob_uop_2_18_is_sys_pc2epc = _RANDOM[11'h454][6];	// rob.scala:310:28
        rob_uop_2_18_flush_on_commit = _RANDOM[11'h454][8];	// rob.scala:310:28
        rob_uop_2_18_ldst = _RANDOM[11'h454][15:10];	// rob.scala:310:28
        rob_uop_2_18_ldst_val = _RANDOM[11'h455][2];	// rob.scala:310:28
        rob_uop_2_18_dst_rtype = _RANDOM[11'h455][4:3];	// rob.scala:310:28
        rob_uop_2_18_fp_val = _RANDOM[11'h455][10];	// rob.scala:310:28
        rob_uop_2_19_uopc = _RANDOM[11'h455][27:21];	// rob.scala:310:28
        rob_uop_2_19_is_rvc = _RANDOM[11'h457][28];	// rob.scala:310:28
        rob_uop_2_19_br_mask = {_RANDOM[11'h45A][31:17], _RANDOM[11'h45B][4:0]};	// rob.scala:310:28
        rob_uop_2_19_ftq_idx = _RANDOM[11'h45B][15:10];	// rob.scala:310:28
        rob_uop_2_19_edge_inst = _RANDOM[11'h45B][16];	// rob.scala:310:28
        rob_uop_2_19_pc_lob = _RANDOM[11'h45B][22:17];	// rob.scala:310:28
        rob_uop_2_19_pdst = _RANDOM[11'h45D][17:11];	// rob.scala:310:28
        rob_uop_2_19_stale_pdst = _RANDOM[11'h45E][23:17];	// rob.scala:310:28
        rob_uop_2_19_is_fencei = _RANDOM[11'h461][3];	// rob.scala:310:28
        rob_uop_2_19_uses_ldq = _RANDOM[11'h461][5];	// rob.scala:310:28
        rob_uop_2_19_uses_stq = _RANDOM[11'h461][6];	// rob.scala:310:28
        rob_uop_2_19_is_sys_pc2epc = _RANDOM[11'h461][7];	// rob.scala:310:28
        rob_uop_2_19_flush_on_commit = _RANDOM[11'h461][9];	// rob.scala:310:28
        rob_uop_2_19_ldst = _RANDOM[11'h461][16:11];	// rob.scala:310:28
        rob_uop_2_19_ldst_val = _RANDOM[11'h462][3];	// rob.scala:310:28
        rob_uop_2_19_dst_rtype = _RANDOM[11'h462][5:4];	// rob.scala:310:28
        rob_uop_2_19_fp_val = _RANDOM[11'h462][11];	// rob.scala:310:28
        rob_uop_2_20_uopc = _RANDOM[11'h462][28:22];	// rob.scala:310:28
        rob_uop_2_20_is_rvc = _RANDOM[11'h464][29];	// rob.scala:310:28
        rob_uop_2_20_br_mask = {_RANDOM[11'h467][31:18], _RANDOM[11'h468][5:0]};	// rob.scala:310:28
        rob_uop_2_20_ftq_idx = _RANDOM[11'h468][16:11];	// rob.scala:310:28
        rob_uop_2_20_edge_inst = _RANDOM[11'h468][17];	// rob.scala:310:28
        rob_uop_2_20_pc_lob = _RANDOM[11'h468][23:18];	// rob.scala:310:28
        rob_uop_2_20_pdst = _RANDOM[11'h46A][18:12];	// rob.scala:310:28
        rob_uop_2_20_stale_pdst = _RANDOM[11'h46B][24:18];	// rob.scala:310:28
        rob_uop_2_20_is_fencei = _RANDOM[11'h46E][4];	// rob.scala:310:28
        rob_uop_2_20_uses_ldq = _RANDOM[11'h46E][6];	// rob.scala:310:28
        rob_uop_2_20_uses_stq = _RANDOM[11'h46E][7];	// rob.scala:310:28
        rob_uop_2_20_is_sys_pc2epc = _RANDOM[11'h46E][8];	// rob.scala:310:28
        rob_uop_2_20_flush_on_commit = _RANDOM[11'h46E][10];	// rob.scala:310:28
        rob_uop_2_20_ldst = _RANDOM[11'h46E][17:12];	// rob.scala:310:28
        rob_uop_2_20_ldst_val = _RANDOM[11'h46F][4];	// rob.scala:310:28
        rob_uop_2_20_dst_rtype = _RANDOM[11'h46F][6:5];	// rob.scala:310:28
        rob_uop_2_20_fp_val = _RANDOM[11'h46F][12];	// rob.scala:310:28
        rob_uop_2_21_uopc = _RANDOM[11'h46F][29:23];	// rob.scala:310:28
        rob_uop_2_21_is_rvc = _RANDOM[11'h471][30];	// rob.scala:310:28
        rob_uop_2_21_br_mask = {_RANDOM[11'h474][31:19], _RANDOM[11'h475][6:0]};	// rob.scala:310:28
        rob_uop_2_21_ftq_idx = _RANDOM[11'h475][17:12];	// rob.scala:310:28
        rob_uop_2_21_edge_inst = _RANDOM[11'h475][18];	// rob.scala:310:28
        rob_uop_2_21_pc_lob = _RANDOM[11'h475][24:19];	// rob.scala:310:28
        rob_uop_2_21_pdst = _RANDOM[11'h477][19:13];	// rob.scala:310:28
        rob_uop_2_21_stale_pdst = _RANDOM[11'h478][25:19];	// rob.scala:310:28
        rob_uop_2_21_is_fencei = _RANDOM[11'h47B][5];	// rob.scala:310:28
        rob_uop_2_21_uses_ldq = _RANDOM[11'h47B][7];	// rob.scala:310:28
        rob_uop_2_21_uses_stq = _RANDOM[11'h47B][8];	// rob.scala:310:28
        rob_uop_2_21_is_sys_pc2epc = _RANDOM[11'h47B][9];	// rob.scala:310:28
        rob_uop_2_21_flush_on_commit = _RANDOM[11'h47B][11];	// rob.scala:310:28
        rob_uop_2_21_ldst = _RANDOM[11'h47B][18:13];	// rob.scala:310:28
        rob_uop_2_21_ldst_val = _RANDOM[11'h47C][5];	// rob.scala:310:28
        rob_uop_2_21_dst_rtype = _RANDOM[11'h47C][7:6];	// rob.scala:310:28
        rob_uop_2_21_fp_val = _RANDOM[11'h47C][13];	// rob.scala:310:28
        rob_uop_2_22_uopc = _RANDOM[11'h47C][30:24];	// rob.scala:310:28
        rob_uop_2_22_is_rvc = _RANDOM[11'h47E][31];	// rob.scala:310:28
        rob_uop_2_22_br_mask = {_RANDOM[11'h481][31:20], _RANDOM[11'h482][7:0]};	// rob.scala:310:28
        rob_uop_2_22_ftq_idx = _RANDOM[11'h482][18:13];	// rob.scala:310:28
        rob_uop_2_22_edge_inst = _RANDOM[11'h482][19];	// rob.scala:310:28
        rob_uop_2_22_pc_lob = _RANDOM[11'h482][25:20];	// rob.scala:310:28
        rob_uop_2_22_pdst = _RANDOM[11'h484][20:14];	// rob.scala:310:28
        rob_uop_2_22_stale_pdst = _RANDOM[11'h485][26:20];	// rob.scala:310:28
        rob_uop_2_22_is_fencei = _RANDOM[11'h488][6];	// rob.scala:310:28
        rob_uop_2_22_uses_ldq = _RANDOM[11'h488][8];	// rob.scala:310:28
        rob_uop_2_22_uses_stq = _RANDOM[11'h488][9];	// rob.scala:310:28
        rob_uop_2_22_is_sys_pc2epc = _RANDOM[11'h488][10];	// rob.scala:310:28
        rob_uop_2_22_flush_on_commit = _RANDOM[11'h488][12];	// rob.scala:310:28
        rob_uop_2_22_ldst = _RANDOM[11'h488][19:14];	// rob.scala:310:28
        rob_uop_2_22_ldst_val = _RANDOM[11'h489][6];	// rob.scala:310:28
        rob_uop_2_22_dst_rtype = _RANDOM[11'h489][8:7];	// rob.scala:310:28
        rob_uop_2_22_fp_val = _RANDOM[11'h489][14];	// rob.scala:310:28
        rob_uop_2_23_uopc = _RANDOM[11'h489][31:25];	// rob.scala:310:28
        rob_uop_2_23_is_rvc = _RANDOM[11'h48C][0];	// rob.scala:310:28
        rob_uop_2_23_br_mask = {_RANDOM[11'h48E][31:21], _RANDOM[11'h48F][8:0]};	// rob.scala:310:28
        rob_uop_2_23_ftq_idx = _RANDOM[11'h48F][19:14];	// rob.scala:310:28
        rob_uop_2_23_edge_inst = _RANDOM[11'h48F][20];	// rob.scala:310:28
        rob_uop_2_23_pc_lob = _RANDOM[11'h48F][26:21];	// rob.scala:310:28
        rob_uop_2_23_pdst = _RANDOM[11'h491][21:15];	// rob.scala:310:28
        rob_uop_2_23_stale_pdst = _RANDOM[11'h492][27:21];	// rob.scala:310:28
        rob_uop_2_23_is_fencei = _RANDOM[11'h495][7];	// rob.scala:310:28
        rob_uop_2_23_uses_ldq = _RANDOM[11'h495][9];	// rob.scala:310:28
        rob_uop_2_23_uses_stq = _RANDOM[11'h495][10];	// rob.scala:310:28
        rob_uop_2_23_is_sys_pc2epc = _RANDOM[11'h495][11];	// rob.scala:310:28
        rob_uop_2_23_flush_on_commit = _RANDOM[11'h495][13];	// rob.scala:310:28
        rob_uop_2_23_ldst = _RANDOM[11'h495][20:15];	// rob.scala:310:28
        rob_uop_2_23_ldst_val = _RANDOM[11'h496][7];	// rob.scala:310:28
        rob_uop_2_23_dst_rtype = _RANDOM[11'h496][9:8];	// rob.scala:310:28
        rob_uop_2_23_fp_val = _RANDOM[11'h496][15];	// rob.scala:310:28
        rob_uop_2_24_uopc = {_RANDOM[11'h496][31:26], _RANDOM[11'h497][0]};	// rob.scala:310:28
        rob_uop_2_24_is_rvc = _RANDOM[11'h499][1];	// rob.scala:310:28
        rob_uop_2_24_br_mask = {_RANDOM[11'h49B][31:22], _RANDOM[11'h49C][9:0]};	// rob.scala:310:28
        rob_uop_2_24_ftq_idx = _RANDOM[11'h49C][20:15];	// rob.scala:310:28
        rob_uop_2_24_edge_inst = _RANDOM[11'h49C][21];	// rob.scala:310:28
        rob_uop_2_24_pc_lob = _RANDOM[11'h49C][27:22];	// rob.scala:310:28
        rob_uop_2_24_pdst = _RANDOM[11'h49E][22:16];	// rob.scala:310:28
        rob_uop_2_24_stale_pdst = _RANDOM[11'h49F][28:22];	// rob.scala:310:28
        rob_uop_2_24_is_fencei = _RANDOM[11'h4A2][8];	// rob.scala:310:28
        rob_uop_2_24_uses_ldq = _RANDOM[11'h4A2][10];	// rob.scala:310:28
        rob_uop_2_24_uses_stq = _RANDOM[11'h4A2][11];	// rob.scala:310:28
        rob_uop_2_24_is_sys_pc2epc = _RANDOM[11'h4A2][12];	// rob.scala:310:28
        rob_uop_2_24_flush_on_commit = _RANDOM[11'h4A2][14];	// rob.scala:310:28
        rob_uop_2_24_ldst = _RANDOM[11'h4A2][21:16];	// rob.scala:310:28
        rob_uop_2_24_ldst_val = _RANDOM[11'h4A3][8];	// rob.scala:310:28
        rob_uop_2_24_dst_rtype = _RANDOM[11'h4A3][10:9];	// rob.scala:310:28
        rob_uop_2_24_fp_val = _RANDOM[11'h4A3][16];	// rob.scala:310:28
        rob_uop_2_25_uopc = {_RANDOM[11'h4A3][31:27], _RANDOM[11'h4A4][1:0]};	// rob.scala:310:28
        rob_uop_2_25_is_rvc = _RANDOM[11'h4A6][2];	// rob.scala:310:28
        rob_uop_2_25_br_mask = {_RANDOM[11'h4A8][31:23], _RANDOM[11'h4A9][10:0]};	// rob.scala:310:28
        rob_uop_2_25_ftq_idx = _RANDOM[11'h4A9][21:16];	// rob.scala:310:28
        rob_uop_2_25_edge_inst = _RANDOM[11'h4A9][22];	// rob.scala:310:28
        rob_uop_2_25_pc_lob = _RANDOM[11'h4A9][28:23];	// rob.scala:310:28
        rob_uop_2_25_pdst = _RANDOM[11'h4AB][23:17];	// rob.scala:310:28
        rob_uop_2_25_stale_pdst = _RANDOM[11'h4AC][29:23];	// rob.scala:310:28
        rob_uop_2_25_is_fencei = _RANDOM[11'h4AF][9];	// rob.scala:310:28
        rob_uop_2_25_uses_ldq = _RANDOM[11'h4AF][11];	// rob.scala:310:28
        rob_uop_2_25_uses_stq = _RANDOM[11'h4AF][12];	// rob.scala:310:28
        rob_uop_2_25_is_sys_pc2epc = _RANDOM[11'h4AF][13];	// rob.scala:310:28
        rob_uop_2_25_flush_on_commit = _RANDOM[11'h4AF][15];	// rob.scala:310:28
        rob_uop_2_25_ldst = _RANDOM[11'h4AF][22:17];	// rob.scala:310:28
        rob_uop_2_25_ldst_val = _RANDOM[11'h4B0][9];	// rob.scala:310:28
        rob_uop_2_25_dst_rtype = _RANDOM[11'h4B0][11:10];	// rob.scala:310:28
        rob_uop_2_25_fp_val = _RANDOM[11'h4B0][17];	// rob.scala:310:28
        rob_uop_2_26_uopc = {_RANDOM[11'h4B0][31:28], _RANDOM[11'h4B1][2:0]};	// rob.scala:310:28
        rob_uop_2_26_is_rvc = _RANDOM[11'h4B3][3];	// rob.scala:310:28
        rob_uop_2_26_br_mask = {_RANDOM[11'h4B5][31:24], _RANDOM[11'h4B6][11:0]};	// rob.scala:310:28
        rob_uop_2_26_ftq_idx = _RANDOM[11'h4B6][22:17];	// rob.scala:310:28
        rob_uop_2_26_edge_inst = _RANDOM[11'h4B6][23];	// rob.scala:310:28
        rob_uop_2_26_pc_lob = _RANDOM[11'h4B6][29:24];	// rob.scala:310:28
        rob_uop_2_26_pdst = _RANDOM[11'h4B8][24:18];	// rob.scala:310:28
        rob_uop_2_26_stale_pdst = _RANDOM[11'h4B9][30:24];	// rob.scala:310:28
        rob_uop_2_26_is_fencei = _RANDOM[11'h4BC][10];	// rob.scala:310:28
        rob_uop_2_26_uses_ldq = _RANDOM[11'h4BC][12];	// rob.scala:310:28
        rob_uop_2_26_uses_stq = _RANDOM[11'h4BC][13];	// rob.scala:310:28
        rob_uop_2_26_is_sys_pc2epc = _RANDOM[11'h4BC][14];	// rob.scala:310:28
        rob_uop_2_26_flush_on_commit = _RANDOM[11'h4BC][16];	// rob.scala:310:28
        rob_uop_2_26_ldst = _RANDOM[11'h4BC][23:18];	// rob.scala:310:28
        rob_uop_2_26_ldst_val = _RANDOM[11'h4BD][10];	// rob.scala:310:28
        rob_uop_2_26_dst_rtype = _RANDOM[11'h4BD][12:11];	// rob.scala:310:28
        rob_uop_2_26_fp_val = _RANDOM[11'h4BD][18];	// rob.scala:310:28
        rob_uop_2_27_uopc = {_RANDOM[11'h4BD][31:29], _RANDOM[11'h4BE][3:0]};	// rob.scala:310:28
        rob_uop_2_27_is_rvc = _RANDOM[11'h4C0][4];	// rob.scala:310:28
        rob_uop_2_27_br_mask = {_RANDOM[11'h4C2][31:25], _RANDOM[11'h4C3][12:0]};	// rob.scala:310:28
        rob_uop_2_27_ftq_idx = _RANDOM[11'h4C3][23:18];	// rob.scala:310:28
        rob_uop_2_27_edge_inst = _RANDOM[11'h4C3][24];	// rob.scala:310:28
        rob_uop_2_27_pc_lob = _RANDOM[11'h4C3][30:25];	// rob.scala:310:28
        rob_uop_2_27_pdst = _RANDOM[11'h4C5][25:19];	// rob.scala:310:28
        rob_uop_2_27_stale_pdst = _RANDOM[11'h4C6][31:25];	// rob.scala:310:28
        rob_uop_2_27_is_fencei = _RANDOM[11'h4C9][11];	// rob.scala:310:28
        rob_uop_2_27_uses_ldq = _RANDOM[11'h4C9][13];	// rob.scala:310:28
        rob_uop_2_27_uses_stq = _RANDOM[11'h4C9][14];	// rob.scala:310:28
        rob_uop_2_27_is_sys_pc2epc = _RANDOM[11'h4C9][15];	// rob.scala:310:28
        rob_uop_2_27_flush_on_commit = _RANDOM[11'h4C9][17];	// rob.scala:310:28
        rob_uop_2_27_ldst = _RANDOM[11'h4C9][24:19];	// rob.scala:310:28
        rob_uop_2_27_ldst_val = _RANDOM[11'h4CA][11];	// rob.scala:310:28
        rob_uop_2_27_dst_rtype = _RANDOM[11'h4CA][13:12];	// rob.scala:310:28
        rob_uop_2_27_fp_val = _RANDOM[11'h4CA][19];	// rob.scala:310:28
        rob_uop_2_28_uopc = {_RANDOM[11'h4CA][31:30], _RANDOM[11'h4CB][4:0]};	// rob.scala:310:28
        rob_uop_2_28_is_rvc = _RANDOM[11'h4CD][5];	// rob.scala:310:28
        rob_uop_2_28_br_mask = {_RANDOM[11'h4CF][31:26], _RANDOM[11'h4D0][13:0]};	// rob.scala:310:28
        rob_uop_2_28_ftq_idx = _RANDOM[11'h4D0][24:19];	// rob.scala:310:28
        rob_uop_2_28_edge_inst = _RANDOM[11'h4D0][25];	// rob.scala:310:28
        rob_uop_2_28_pc_lob = _RANDOM[11'h4D0][31:26];	// rob.scala:310:28
        rob_uop_2_28_pdst = _RANDOM[11'h4D2][26:20];	// rob.scala:310:28
        rob_uop_2_28_stale_pdst = {_RANDOM[11'h4D3][31:26], _RANDOM[11'h4D4][0]};	// rob.scala:310:28
        rob_uop_2_28_is_fencei = _RANDOM[11'h4D6][12];	// rob.scala:310:28
        rob_uop_2_28_uses_ldq = _RANDOM[11'h4D6][14];	// rob.scala:310:28
        rob_uop_2_28_uses_stq = _RANDOM[11'h4D6][15];	// rob.scala:310:28
        rob_uop_2_28_is_sys_pc2epc = _RANDOM[11'h4D6][16];	// rob.scala:310:28
        rob_uop_2_28_flush_on_commit = _RANDOM[11'h4D6][18];	// rob.scala:310:28
        rob_uop_2_28_ldst = _RANDOM[11'h4D6][25:20];	// rob.scala:310:28
        rob_uop_2_28_ldst_val = _RANDOM[11'h4D7][12];	// rob.scala:310:28
        rob_uop_2_28_dst_rtype = _RANDOM[11'h4D7][14:13];	// rob.scala:310:28
        rob_uop_2_28_fp_val = _RANDOM[11'h4D7][20];	// rob.scala:310:28
        rob_uop_2_29_uopc = {_RANDOM[11'h4D7][31], _RANDOM[11'h4D8][5:0]};	// rob.scala:310:28
        rob_uop_2_29_is_rvc = _RANDOM[11'h4DA][6];	// rob.scala:310:28
        rob_uop_2_29_br_mask = {_RANDOM[11'h4DC][31:27], _RANDOM[11'h4DD][14:0]};	// rob.scala:310:28
        rob_uop_2_29_ftq_idx = _RANDOM[11'h4DD][25:20];	// rob.scala:310:28
        rob_uop_2_29_edge_inst = _RANDOM[11'h4DD][26];	// rob.scala:310:28
        rob_uop_2_29_pc_lob = {_RANDOM[11'h4DD][31:27], _RANDOM[11'h4DE][0]};	// rob.scala:310:28
        rob_uop_2_29_pdst = _RANDOM[11'h4DF][27:21];	// rob.scala:310:28
        rob_uop_2_29_stale_pdst = {_RANDOM[11'h4E0][31:27], _RANDOM[11'h4E1][1:0]};	// rob.scala:310:28
        rob_uop_2_29_is_fencei = _RANDOM[11'h4E3][13];	// rob.scala:310:28
        rob_uop_2_29_uses_ldq = _RANDOM[11'h4E3][15];	// rob.scala:310:28
        rob_uop_2_29_uses_stq = _RANDOM[11'h4E3][16];	// rob.scala:310:28
        rob_uop_2_29_is_sys_pc2epc = _RANDOM[11'h4E3][17];	// rob.scala:310:28
        rob_uop_2_29_flush_on_commit = _RANDOM[11'h4E3][19];	// rob.scala:310:28
        rob_uop_2_29_ldst = _RANDOM[11'h4E3][26:21];	// rob.scala:310:28
        rob_uop_2_29_ldst_val = _RANDOM[11'h4E4][13];	// rob.scala:310:28
        rob_uop_2_29_dst_rtype = _RANDOM[11'h4E4][15:14];	// rob.scala:310:28
        rob_uop_2_29_fp_val = _RANDOM[11'h4E4][21];	// rob.scala:310:28
        rob_uop_2_30_uopc = _RANDOM[11'h4E5][6:0];	// rob.scala:310:28
        rob_uop_2_30_is_rvc = _RANDOM[11'h4E7][7];	// rob.scala:310:28
        rob_uop_2_30_br_mask = {_RANDOM[11'h4E9][31:28], _RANDOM[11'h4EA][15:0]};	// rob.scala:310:28
        rob_uop_2_30_ftq_idx = _RANDOM[11'h4EA][26:21];	// rob.scala:310:28
        rob_uop_2_30_edge_inst = _RANDOM[11'h4EA][27];	// rob.scala:310:28
        rob_uop_2_30_pc_lob = {_RANDOM[11'h4EA][31:28], _RANDOM[11'h4EB][1:0]};	// rob.scala:310:28
        rob_uop_2_30_pdst = _RANDOM[11'h4EC][28:22];	// rob.scala:310:28
        rob_uop_2_30_stale_pdst = {_RANDOM[11'h4ED][31:28], _RANDOM[11'h4EE][2:0]};	// rob.scala:310:28
        rob_uop_2_30_is_fencei = _RANDOM[11'h4F0][14];	// rob.scala:310:28
        rob_uop_2_30_uses_ldq = _RANDOM[11'h4F0][16];	// rob.scala:310:28
        rob_uop_2_30_uses_stq = _RANDOM[11'h4F0][17];	// rob.scala:310:28
        rob_uop_2_30_is_sys_pc2epc = _RANDOM[11'h4F0][18];	// rob.scala:310:28
        rob_uop_2_30_flush_on_commit = _RANDOM[11'h4F0][20];	// rob.scala:310:28
        rob_uop_2_30_ldst = _RANDOM[11'h4F0][27:22];	// rob.scala:310:28
        rob_uop_2_30_ldst_val = _RANDOM[11'h4F1][14];	// rob.scala:310:28
        rob_uop_2_30_dst_rtype = _RANDOM[11'h4F1][16:15];	// rob.scala:310:28
        rob_uop_2_30_fp_val = _RANDOM[11'h4F1][22];	// rob.scala:310:28
        rob_uop_2_31_uopc = _RANDOM[11'h4F2][7:1];	// rob.scala:310:28
        rob_uop_2_31_is_rvc = _RANDOM[11'h4F4][8];	// rob.scala:310:28
        rob_uop_2_31_br_mask = {_RANDOM[11'h4F6][31:29], _RANDOM[11'h4F7][16:0]};	// rob.scala:310:28
        rob_uop_2_31_ftq_idx = _RANDOM[11'h4F7][27:22];	// rob.scala:310:28
        rob_uop_2_31_edge_inst = _RANDOM[11'h4F7][28];	// rob.scala:310:28
        rob_uop_2_31_pc_lob = {_RANDOM[11'h4F7][31:29], _RANDOM[11'h4F8][2:0]};	// rob.scala:310:28
        rob_uop_2_31_pdst = _RANDOM[11'h4F9][29:23];	// rob.scala:310:28
        rob_uop_2_31_stale_pdst = {_RANDOM[11'h4FA][31:29], _RANDOM[11'h4FB][3:0]};	// rob.scala:310:28
        rob_uop_2_31_is_fencei = _RANDOM[11'h4FD][15];	// rob.scala:310:28
        rob_uop_2_31_uses_ldq = _RANDOM[11'h4FD][17];	// rob.scala:310:28
        rob_uop_2_31_uses_stq = _RANDOM[11'h4FD][18];	// rob.scala:310:28
        rob_uop_2_31_is_sys_pc2epc = _RANDOM[11'h4FD][19];	// rob.scala:310:28
        rob_uop_2_31_flush_on_commit = _RANDOM[11'h4FD][21];	// rob.scala:310:28
        rob_uop_2_31_ldst = _RANDOM[11'h4FD][28:23];	// rob.scala:310:28
        rob_uop_2_31_ldst_val = _RANDOM[11'h4FE][15];	// rob.scala:310:28
        rob_uop_2_31_dst_rtype = _RANDOM[11'h4FE][17:16];	// rob.scala:310:28
        rob_uop_2_31_fp_val = _RANDOM[11'h4FE][23];	// rob.scala:310:28
        rob_exception_2_0 = _RANDOM[11'h4FF][2];	// rob.scala:311:28
        rob_exception_2_1 = _RANDOM[11'h4FF][3];	// rob.scala:311:28
        rob_exception_2_2 = _RANDOM[11'h4FF][4];	// rob.scala:311:28
        rob_exception_2_3 = _RANDOM[11'h4FF][5];	// rob.scala:311:28
        rob_exception_2_4 = _RANDOM[11'h4FF][6];	// rob.scala:311:28
        rob_exception_2_5 = _RANDOM[11'h4FF][7];	// rob.scala:311:28
        rob_exception_2_6 = _RANDOM[11'h4FF][8];	// rob.scala:311:28
        rob_exception_2_7 = _RANDOM[11'h4FF][9];	// rob.scala:311:28
        rob_exception_2_8 = _RANDOM[11'h4FF][10];	// rob.scala:311:28
        rob_exception_2_9 = _RANDOM[11'h4FF][11];	// rob.scala:311:28
        rob_exception_2_10 = _RANDOM[11'h4FF][12];	// rob.scala:311:28
        rob_exception_2_11 = _RANDOM[11'h4FF][13];	// rob.scala:311:28
        rob_exception_2_12 = _RANDOM[11'h4FF][14];	// rob.scala:311:28
        rob_exception_2_13 = _RANDOM[11'h4FF][15];	// rob.scala:311:28
        rob_exception_2_14 = _RANDOM[11'h4FF][16];	// rob.scala:311:28
        rob_exception_2_15 = _RANDOM[11'h4FF][17];	// rob.scala:311:28
        rob_exception_2_16 = _RANDOM[11'h4FF][18];	// rob.scala:311:28
        rob_exception_2_17 = _RANDOM[11'h4FF][19];	// rob.scala:311:28
        rob_exception_2_18 = _RANDOM[11'h4FF][20];	// rob.scala:311:28
        rob_exception_2_19 = _RANDOM[11'h4FF][21];	// rob.scala:311:28
        rob_exception_2_20 = _RANDOM[11'h4FF][22];	// rob.scala:311:28
        rob_exception_2_21 = _RANDOM[11'h4FF][23];	// rob.scala:311:28
        rob_exception_2_22 = _RANDOM[11'h4FF][24];	// rob.scala:311:28
        rob_exception_2_23 = _RANDOM[11'h4FF][25];	// rob.scala:311:28
        rob_exception_2_24 = _RANDOM[11'h4FF][26];	// rob.scala:311:28
        rob_exception_2_25 = _RANDOM[11'h4FF][27];	// rob.scala:311:28
        rob_exception_2_26 = _RANDOM[11'h4FF][28];	// rob.scala:311:28
        rob_exception_2_27 = _RANDOM[11'h4FF][29];	// rob.scala:311:28
        rob_exception_2_28 = _RANDOM[11'h4FF][30];	// rob.scala:311:28
        rob_exception_2_29 = _RANDOM[11'h4FF][31];	// rob.scala:311:28
        rob_exception_2_30 = _RANDOM[11'h500][0];	// rob.scala:311:28
        rob_exception_2_31 = _RANDOM[11'h500][1];	// rob.scala:311:28
        rob_predicated_2_0 = _RANDOM[11'h500][2];	// rob.scala:311:28, :312:29
        rob_predicated_2_1 = _RANDOM[11'h500][3];	// rob.scala:311:28, :312:29
        rob_predicated_2_2 = _RANDOM[11'h500][4];	// rob.scala:311:28, :312:29
        rob_predicated_2_3 = _RANDOM[11'h500][5];	// rob.scala:311:28, :312:29
        rob_predicated_2_4 = _RANDOM[11'h500][6];	// rob.scala:311:28, :312:29
        rob_predicated_2_5 = _RANDOM[11'h500][7];	// rob.scala:311:28, :312:29
        rob_predicated_2_6 = _RANDOM[11'h500][8];	// rob.scala:311:28, :312:29
        rob_predicated_2_7 = _RANDOM[11'h500][9];	// rob.scala:311:28, :312:29
        rob_predicated_2_8 = _RANDOM[11'h500][10];	// rob.scala:311:28, :312:29
        rob_predicated_2_9 = _RANDOM[11'h500][11];	// rob.scala:311:28, :312:29
        rob_predicated_2_10 = _RANDOM[11'h500][12];	// rob.scala:311:28, :312:29
        rob_predicated_2_11 = _RANDOM[11'h500][13];	// rob.scala:311:28, :312:29
        rob_predicated_2_12 = _RANDOM[11'h500][14];	// rob.scala:311:28, :312:29
        rob_predicated_2_13 = _RANDOM[11'h500][15];	// rob.scala:311:28, :312:29
        rob_predicated_2_14 = _RANDOM[11'h500][16];	// rob.scala:311:28, :312:29
        rob_predicated_2_15 = _RANDOM[11'h500][17];	// rob.scala:311:28, :312:29
        rob_predicated_2_16 = _RANDOM[11'h500][18];	// rob.scala:311:28, :312:29
        rob_predicated_2_17 = _RANDOM[11'h500][19];	// rob.scala:311:28, :312:29
        rob_predicated_2_18 = _RANDOM[11'h500][20];	// rob.scala:311:28, :312:29
        rob_predicated_2_19 = _RANDOM[11'h500][21];	// rob.scala:311:28, :312:29
        rob_predicated_2_20 = _RANDOM[11'h500][22];	// rob.scala:311:28, :312:29
        rob_predicated_2_21 = _RANDOM[11'h500][23];	// rob.scala:311:28, :312:29
        rob_predicated_2_22 = _RANDOM[11'h500][24];	// rob.scala:311:28, :312:29
        rob_predicated_2_23 = _RANDOM[11'h500][25];	// rob.scala:311:28, :312:29
        rob_predicated_2_24 = _RANDOM[11'h500][26];	// rob.scala:311:28, :312:29
        rob_predicated_2_25 = _RANDOM[11'h500][27];	// rob.scala:311:28, :312:29
        rob_predicated_2_26 = _RANDOM[11'h500][28];	// rob.scala:311:28, :312:29
        rob_predicated_2_27 = _RANDOM[11'h500][29];	// rob.scala:311:28, :312:29
        rob_predicated_2_28 = _RANDOM[11'h500][30];	// rob.scala:311:28, :312:29
        rob_predicated_2_29 = _RANDOM[11'h500][31];	// rob.scala:311:28, :312:29
        rob_predicated_2_30 = _RANDOM[11'h501][0];	// rob.scala:312:29
        rob_predicated_2_31 = _RANDOM[11'h501][1];	// rob.scala:312:29
        rob_val_3_0 = _RANDOM[11'h501][2];	// rob.scala:307:32, :312:29
        rob_val_3_1 = _RANDOM[11'h501][3];	// rob.scala:307:32, :312:29
        rob_val_3_2 = _RANDOM[11'h501][4];	// rob.scala:307:32, :312:29
        rob_val_3_3 = _RANDOM[11'h501][5];	// rob.scala:307:32, :312:29
        rob_val_3_4 = _RANDOM[11'h501][6];	// rob.scala:307:32, :312:29
        rob_val_3_5 = _RANDOM[11'h501][7];	// rob.scala:307:32, :312:29
        rob_val_3_6 = _RANDOM[11'h501][8];	// rob.scala:307:32, :312:29
        rob_val_3_7 = _RANDOM[11'h501][9];	// rob.scala:307:32, :312:29
        rob_val_3_8 = _RANDOM[11'h501][10];	// rob.scala:307:32, :312:29
        rob_val_3_9 = _RANDOM[11'h501][11];	// rob.scala:307:32, :312:29
        rob_val_3_10 = _RANDOM[11'h501][12];	// rob.scala:307:32, :312:29
        rob_val_3_11 = _RANDOM[11'h501][13];	// rob.scala:307:32, :312:29
        rob_val_3_12 = _RANDOM[11'h501][14];	// rob.scala:307:32, :312:29
        rob_val_3_13 = _RANDOM[11'h501][15];	// rob.scala:307:32, :312:29
        rob_val_3_14 = _RANDOM[11'h501][16];	// rob.scala:307:32, :312:29
        rob_val_3_15 = _RANDOM[11'h501][17];	// rob.scala:307:32, :312:29
        rob_val_3_16 = _RANDOM[11'h501][18];	// rob.scala:307:32, :312:29
        rob_val_3_17 = _RANDOM[11'h501][19];	// rob.scala:307:32, :312:29
        rob_val_3_18 = _RANDOM[11'h501][20];	// rob.scala:307:32, :312:29
        rob_val_3_19 = _RANDOM[11'h501][21];	// rob.scala:307:32, :312:29
        rob_val_3_20 = _RANDOM[11'h501][22];	// rob.scala:307:32, :312:29
        rob_val_3_21 = _RANDOM[11'h501][23];	// rob.scala:307:32, :312:29
        rob_val_3_22 = _RANDOM[11'h501][24];	// rob.scala:307:32, :312:29
        rob_val_3_23 = _RANDOM[11'h501][25];	// rob.scala:307:32, :312:29
        rob_val_3_24 = _RANDOM[11'h501][26];	// rob.scala:307:32, :312:29
        rob_val_3_25 = _RANDOM[11'h501][27];	// rob.scala:307:32, :312:29
        rob_val_3_26 = _RANDOM[11'h501][28];	// rob.scala:307:32, :312:29
        rob_val_3_27 = _RANDOM[11'h501][29];	// rob.scala:307:32, :312:29
        rob_val_3_28 = _RANDOM[11'h501][30];	// rob.scala:307:32, :312:29
        rob_val_3_29 = _RANDOM[11'h501][31];	// rob.scala:307:32, :312:29
        rob_val_3_30 = _RANDOM[11'h502][0];	// rob.scala:307:32
        rob_val_3_31 = _RANDOM[11'h502][1];	// rob.scala:307:32
        rob_bsy_3_0 = _RANDOM[11'h502][2];	// rob.scala:307:32, :308:28
        rob_bsy_3_1 = _RANDOM[11'h502][3];	// rob.scala:307:32, :308:28
        rob_bsy_3_2 = _RANDOM[11'h502][4];	// rob.scala:307:32, :308:28
        rob_bsy_3_3 = _RANDOM[11'h502][5];	// rob.scala:307:32, :308:28
        rob_bsy_3_4 = _RANDOM[11'h502][6];	// rob.scala:307:32, :308:28
        rob_bsy_3_5 = _RANDOM[11'h502][7];	// rob.scala:307:32, :308:28
        rob_bsy_3_6 = _RANDOM[11'h502][8];	// rob.scala:307:32, :308:28
        rob_bsy_3_7 = _RANDOM[11'h502][9];	// rob.scala:307:32, :308:28
        rob_bsy_3_8 = _RANDOM[11'h502][10];	// rob.scala:307:32, :308:28
        rob_bsy_3_9 = _RANDOM[11'h502][11];	// rob.scala:307:32, :308:28
        rob_bsy_3_10 = _RANDOM[11'h502][12];	// rob.scala:307:32, :308:28
        rob_bsy_3_11 = _RANDOM[11'h502][13];	// rob.scala:307:32, :308:28
        rob_bsy_3_12 = _RANDOM[11'h502][14];	// rob.scala:307:32, :308:28
        rob_bsy_3_13 = _RANDOM[11'h502][15];	// rob.scala:307:32, :308:28
        rob_bsy_3_14 = _RANDOM[11'h502][16];	// rob.scala:307:32, :308:28
        rob_bsy_3_15 = _RANDOM[11'h502][17];	// rob.scala:307:32, :308:28
        rob_bsy_3_16 = _RANDOM[11'h502][18];	// rob.scala:307:32, :308:28
        rob_bsy_3_17 = _RANDOM[11'h502][19];	// rob.scala:307:32, :308:28
        rob_bsy_3_18 = _RANDOM[11'h502][20];	// rob.scala:307:32, :308:28
        rob_bsy_3_19 = _RANDOM[11'h502][21];	// rob.scala:307:32, :308:28
        rob_bsy_3_20 = _RANDOM[11'h502][22];	// rob.scala:307:32, :308:28
        rob_bsy_3_21 = _RANDOM[11'h502][23];	// rob.scala:307:32, :308:28
        rob_bsy_3_22 = _RANDOM[11'h502][24];	// rob.scala:307:32, :308:28
        rob_bsy_3_23 = _RANDOM[11'h502][25];	// rob.scala:307:32, :308:28
        rob_bsy_3_24 = _RANDOM[11'h502][26];	// rob.scala:307:32, :308:28
        rob_bsy_3_25 = _RANDOM[11'h502][27];	// rob.scala:307:32, :308:28
        rob_bsy_3_26 = _RANDOM[11'h502][28];	// rob.scala:307:32, :308:28
        rob_bsy_3_27 = _RANDOM[11'h502][29];	// rob.scala:307:32, :308:28
        rob_bsy_3_28 = _RANDOM[11'h502][30];	// rob.scala:307:32, :308:28
        rob_bsy_3_29 = _RANDOM[11'h502][31];	// rob.scala:307:32, :308:28
        rob_bsy_3_30 = _RANDOM[11'h503][0];	// rob.scala:308:28
        rob_bsy_3_31 = _RANDOM[11'h503][1];	// rob.scala:308:28
        rob_unsafe_3_0 = _RANDOM[11'h503][2];	// rob.scala:308:28, :309:28
        rob_unsafe_3_1 = _RANDOM[11'h503][3];	// rob.scala:308:28, :309:28
        rob_unsafe_3_2 = _RANDOM[11'h503][4];	// rob.scala:308:28, :309:28
        rob_unsafe_3_3 = _RANDOM[11'h503][5];	// rob.scala:308:28, :309:28
        rob_unsafe_3_4 = _RANDOM[11'h503][6];	// rob.scala:308:28, :309:28
        rob_unsafe_3_5 = _RANDOM[11'h503][7];	// rob.scala:308:28, :309:28
        rob_unsafe_3_6 = _RANDOM[11'h503][8];	// rob.scala:308:28, :309:28
        rob_unsafe_3_7 = _RANDOM[11'h503][9];	// rob.scala:308:28, :309:28
        rob_unsafe_3_8 = _RANDOM[11'h503][10];	// rob.scala:308:28, :309:28
        rob_unsafe_3_9 = _RANDOM[11'h503][11];	// rob.scala:308:28, :309:28
        rob_unsafe_3_10 = _RANDOM[11'h503][12];	// rob.scala:308:28, :309:28
        rob_unsafe_3_11 = _RANDOM[11'h503][13];	// rob.scala:308:28, :309:28
        rob_unsafe_3_12 = _RANDOM[11'h503][14];	// rob.scala:308:28, :309:28
        rob_unsafe_3_13 = _RANDOM[11'h503][15];	// rob.scala:308:28, :309:28
        rob_unsafe_3_14 = _RANDOM[11'h503][16];	// rob.scala:308:28, :309:28
        rob_unsafe_3_15 = _RANDOM[11'h503][17];	// rob.scala:308:28, :309:28
        rob_unsafe_3_16 = _RANDOM[11'h503][18];	// rob.scala:308:28, :309:28
        rob_unsafe_3_17 = _RANDOM[11'h503][19];	// rob.scala:308:28, :309:28
        rob_unsafe_3_18 = _RANDOM[11'h503][20];	// rob.scala:308:28, :309:28
        rob_unsafe_3_19 = _RANDOM[11'h503][21];	// rob.scala:308:28, :309:28
        rob_unsafe_3_20 = _RANDOM[11'h503][22];	// rob.scala:308:28, :309:28
        rob_unsafe_3_21 = _RANDOM[11'h503][23];	// rob.scala:308:28, :309:28
        rob_unsafe_3_22 = _RANDOM[11'h503][24];	// rob.scala:308:28, :309:28
        rob_unsafe_3_23 = _RANDOM[11'h503][25];	// rob.scala:308:28, :309:28
        rob_unsafe_3_24 = _RANDOM[11'h503][26];	// rob.scala:308:28, :309:28
        rob_unsafe_3_25 = _RANDOM[11'h503][27];	// rob.scala:308:28, :309:28
        rob_unsafe_3_26 = _RANDOM[11'h503][28];	// rob.scala:308:28, :309:28
        rob_unsafe_3_27 = _RANDOM[11'h503][29];	// rob.scala:308:28, :309:28
        rob_unsafe_3_28 = _RANDOM[11'h503][30];	// rob.scala:308:28, :309:28
        rob_unsafe_3_29 = _RANDOM[11'h503][31];	// rob.scala:308:28, :309:28
        rob_unsafe_3_30 = _RANDOM[11'h504][0];	// rob.scala:309:28
        rob_unsafe_3_31 = _RANDOM[11'h504][1];	// rob.scala:309:28
        rob_uop_3_0_uopc = _RANDOM[11'h504][8:2];	// rob.scala:309:28, :310:28
        rob_uop_3_0_is_rvc = _RANDOM[11'h506][9];	// rob.scala:310:28
        rob_uop_3_0_br_mask = {_RANDOM[11'h508][31:30], _RANDOM[11'h509][17:0]};	// rob.scala:310:28
        rob_uop_3_0_ftq_idx = _RANDOM[11'h509][28:23];	// rob.scala:310:28
        rob_uop_3_0_edge_inst = _RANDOM[11'h509][29];	// rob.scala:310:28
        rob_uop_3_0_pc_lob = {_RANDOM[11'h509][31:30], _RANDOM[11'h50A][3:0]};	// rob.scala:310:28
        rob_uop_3_0_pdst = _RANDOM[11'h50B][30:24];	// rob.scala:310:28
        rob_uop_3_0_stale_pdst = {_RANDOM[11'h50C][31:30], _RANDOM[11'h50D][4:0]};	// rob.scala:310:28
        rob_uop_3_0_is_fencei = _RANDOM[11'h50F][16];	// rob.scala:310:28
        rob_uop_3_0_uses_ldq = _RANDOM[11'h50F][18];	// rob.scala:310:28
        rob_uop_3_0_uses_stq = _RANDOM[11'h50F][19];	// rob.scala:310:28
        rob_uop_3_0_is_sys_pc2epc = _RANDOM[11'h50F][20];	// rob.scala:310:28
        rob_uop_3_0_flush_on_commit = _RANDOM[11'h50F][22];	// rob.scala:310:28
        rob_uop_3_0_ldst = _RANDOM[11'h50F][29:24];	// rob.scala:310:28
        rob_uop_3_0_ldst_val = _RANDOM[11'h510][16];	// rob.scala:310:28
        rob_uop_3_0_dst_rtype = _RANDOM[11'h510][18:17];	// rob.scala:310:28
        rob_uop_3_0_fp_val = _RANDOM[11'h510][24];	// rob.scala:310:28
        rob_uop_3_1_uopc = _RANDOM[11'h511][9:3];	// rob.scala:310:28
        rob_uop_3_1_is_rvc = _RANDOM[11'h513][10];	// rob.scala:310:28
        rob_uop_3_1_br_mask = {_RANDOM[11'h515][31], _RANDOM[11'h516][18:0]};	// rob.scala:310:28
        rob_uop_3_1_ftq_idx = _RANDOM[11'h516][29:24];	// rob.scala:310:28
        rob_uop_3_1_edge_inst = _RANDOM[11'h516][30];	// rob.scala:310:28
        rob_uop_3_1_pc_lob = {_RANDOM[11'h516][31], _RANDOM[11'h517][4:0]};	// rob.scala:310:28
        rob_uop_3_1_pdst = _RANDOM[11'h518][31:25];	// rob.scala:310:28
        rob_uop_3_1_stale_pdst = {_RANDOM[11'h519][31], _RANDOM[11'h51A][5:0]};	// rob.scala:310:28
        rob_uop_3_1_is_fencei = _RANDOM[11'h51C][17];	// rob.scala:310:28
        rob_uop_3_1_uses_ldq = _RANDOM[11'h51C][19];	// rob.scala:310:28
        rob_uop_3_1_uses_stq = _RANDOM[11'h51C][20];	// rob.scala:310:28
        rob_uop_3_1_is_sys_pc2epc = _RANDOM[11'h51C][21];	// rob.scala:310:28
        rob_uop_3_1_flush_on_commit = _RANDOM[11'h51C][23];	// rob.scala:310:28
        rob_uop_3_1_ldst = _RANDOM[11'h51C][30:25];	// rob.scala:310:28
        rob_uop_3_1_ldst_val = _RANDOM[11'h51D][17];	// rob.scala:310:28
        rob_uop_3_1_dst_rtype = _RANDOM[11'h51D][19:18];	// rob.scala:310:28
        rob_uop_3_1_fp_val = _RANDOM[11'h51D][25];	// rob.scala:310:28
        rob_uop_3_2_uopc = _RANDOM[11'h51E][10:4];	// rob.scala:310:28
        rob_uop_3_2_is_rvc = _RANDOM[11'h520][11];	// rob.scala:310:28
        rob_uop_3_2_br_mask = _RANDOM[11'h523][19:0];	// rob.scala:310:28
        rob_uop_3_2_ftq_idx = _RANDOM[11'h523][30:25];	// rob.scala:310:28
        rob_uop_3_2_edge_inst = _RANDOM[11'h523][31];	// rob.scala:310:28
        rob_uop_3_2_pc_lob = _RANDOM[11'h524][5:0];	// rob.scala:310:28
        rob_uop_3_2_pdst = {_RANDOM[11'h525][31:26], _RANDOM[11'h526][0]};	// rob.scala:310:28
        rob_uop_3_2_stale_pdst = _RANDOM[11'h527][6:0];	// rob.scala:310:28
        rob_uop_3_2_is_fencei = _RANDOM[11'h529][18];	// rob.scala:310:28
        rob_uop_3_2_uses_ldq = _RANDOM[11'h529][20];	// rob.scala:310:28
        rob_uop_3_2_uses_stq = _RANDOM[11'h529][21];	// rob.scala:310:28
        rob_uop_3_2_is_sys_pc2epc = _RANDOM[11'h529][22];	// rob.scala:310:28
        rob_uop_3_2_flush_on_commit = _RANDOM[11'h529][24];	// rob.scala:310:28
        rob_uop_3_2_ldst = _RANDOM[11'h529][31:26];	// rob.scala:310:28
        rob_uop_3_2_ldst_val = _RANDOM[11'h52A][18];	// rob.scala:310:28
        rob_uop_3_2_dst_rtype = _RANDOM[11'h52A][20:19];	// rob.scala:310:28
        rob_uop_3_2_fp_val = _RANDOM[11'h52A][26];	// rob.scala:310:28
        rob_uop_3_3_uopc = _RANDOM[11'h52B][11:5];	// rob.scala:310:28
        rob_uop_3_3_is_rvc = _RANDOM[11'h52D][12];	// rob.scala:310:28
        rob_uop_3_3_br_mask = _RANDOM[11'h530][20:1];	// rob.scala:310:28
        rob_uop_3_3_ftq_idx = _RANDOM[11'h530][31:26];	// rob.scala:310:28
        rob_uop_3_3_edge_inst = _RANDOM[11'h531][0];	// rob.scala:310:28
        rob_uop_3_3_pc_lob = _RANDOM[11'h531][6:1];	// rob.scala:310:28
        rob_uop_3_3_pdst = {_RANDOM[11'h532][31:27], _RANDOM[11'h533][1:0]};	// rob.scala:310:28
        rob_uop_3_3_stale_pdst = _RANDOM[11'h534][7:1];	// rob.scala:310:28
        rob_uop_3_3_is_fencei = _RANDOM[11'h536][19];	// rob.scala:310:28
        rob_uop_3_3_uses_ldq = _RANDOM[11'h536][21];	// rob.scala:310:28
        rob_uop_3_3_uses_stq = _RANDOM[11'h536][22];	// rob.scala:310:28
        rob_uop_3_3_is_sys_pc2epc = _RANDOM[11'h536][23];	// rob.scala:310:28
        rob_uop_3_3_flush_on_commit = _RANDOM[11'h536][25];	// rob.scala:310:28
        rob_uop_3_3_ldst = {_RANDOM[11'h536][31:27], _RANDOM[11'h537][0]};	// rob.scala:310:28
        rob_uop_3_3_ldst_val = _RANDOM[11'h537][19];	// rob.scala:310:28
        rob_uop_3_3_dst_rtype = _RANDOM[11'h537][21:20];	// rob.scala:310:28
        rob_uop_3_3_fp_val = _RANDOM[11'h537][27];	// rob.scala:310:28
        rob_uop_3_4_uopc = _RANDOM[11'h538][12:6];	// rob.scala:310:28
        rob_uop_3_4_is_rvc = _RANDOM[11'h53A][13];	// rob.scala:310:28
        rob_uop_3_4_br_mask = _RANDOM[11'h53D][21:2];	// rob.scala:310:28
        rob_uop_3_4_ftq_idx = {_RANDOM[11'h53D][31:27], _RANDOM[11'h53E][0]};	// rob.scala:310:28
        rob_uop_3_4_edge_inst = _RANDOM[11'h53E][1];	// rob.scala:310:28
        rob_uop_3_4_pc_lob = _RANDOM[11'h53E][7:2];	// rob.scala:310:28
        rob_uop_3_4_pdst = {_RANDOM[11'h53F][31:28], _RANDOM[11'h540][2:0]};	// rob.scala:310:28
        rob_uop_3_4_stale_pdst = _RANDOM[11'h541][8:2];	// rob.scala:310:28
        rob_uop_3_4_is_fencei = _RANDOM[11'h543][20];	// rob.scala:310:28
        rob_uop_3_4_uses_ldq = _RANDOM[11'h543][22];	// rob.scala:310:28
        rob_uop_3_4_uses_stq = _RANDOM[11'h543][23];	// rob.scala:310:28
        rob_uop_3_4_is_sys_pc2epc = _RANDOM[11'h543][24];	// rob.scala:310:28
        rob_uop_3_4_flush_on_commit = _RANDOM[11'h543][26];	// rob.scala:310:28
        rob_uop_3_4_ldst = {_RANDOM[11'h543][31:28], _RANDOM[11'h544][1:0]};	// rob.scala:310:28
        rob_uop_3_4_ldst_val = _RANDOM[11'h544][20];	// rob.scala:310:28
        rob_uop_3_4_dst_rtype = _RANDOM[11'h544][22:21];	// rob.scala:310:28
        rob_uop_3_4_fp_val = _RANDOM[11'h544][28];	// rob.scala:310:28
        rob_uop_3_5_uopc = _RANDOM[11'h545][13:7];	// rob.scala:310:28
        rob_uop_3_5_is_rvc = _RANDOM[11'h547][14];	// rob.scala:310:28
        rob_uop_3_5_br_mask = _RANDOM[11'h54A][22:3];	// rob.scala:310:28
        rob_uop_3_5_ftq_idx = {_RANDOM[11'h54A][31:28], _RANDOM[11'h54B][1:0]};	// rob.scala:310:28
        rob_uop_3_5_edge_inst = _RANDOM[11'h54B][2];	// rob.scala:310:28
        rob_uop_3_5_pc_lob = _RANDOM[11'h54B][8:3];	// rob.scala:310:28
        rob_uop_3_5_pdst = {_RANDOM[11'h54C][31:29], _RANDOM[11'h54D][3:0]};	// rob.scala:310:28
        rob_uop_3_5_stale_pdst = _RANDOM[11'h54E][9:3];	// rob.scala:310:28
        rob_uop_3_5_is_fencei = _RANDOM[11'h550][21];	// rob.scala:310:28
        rob_uop_3_5_uses_ldq = _RANDOM[11'h550][23];	// rob.scala:310:28
        rob_uop_3_5_uses_stq = _RANDOM[11'h550][24];	// rob.scala:310:28
        rob_uop_3_5_is_sys_pc2epc = _RANDOM[11'h550][25];	// rob.scala:310:28
        rob_uop_3_5_flush_on_commit = _RANDOM[11'h550][27];	// rob.scala:310:28
        rob_uop_3_5_ldst = {_RANDOM[11'h550][31:29], _RANDOM[11'h551][2:0]};	// rob.scala:310:28
        rob_uop_3_5_ldst_val = _RANDOM[11'h551][21];	// rob.scala:310:28
        rob_uop_3_5_dst_rtype = _RANDOM[11'h551][23:22];	// rob.scala:310:28
        rob_uop_3_5_fp_val = _RANDOM[11'h551][29];	// rob.scala:310:28
        rob_uop_3_6_uopc = _RANDOM[11'h552][14:8];	// rob.scala:310:28
        rob_uop_3_6_is_rvc = _RANDOM[11'h554][15];	// rob.scala:310:28
        rob_uop_3_6_br_mask = _RANDOM[11'h557][23:4];	// rob.scala:310:28
        rob_uop_3_6_ftq_idx = {_RANDOM[11'h557][31:29], _RANDOM[11'h558][2:0]};	// rob.scala:310:28
        rob_uop_3_6_edge_inst = _RANDOM[11'h558][3];	// rob.scala:310:28
        rob_uop_3_6_pc_lob = _RANDOM[11'h558][9:4];	// rob.scala:310:28
        rob_uop_3_6_pdst = {_RANDOM[11'h559][31:30], _RANDOM[11'h55A][4:0]};	// rob.scala:310:28
        rob_uop_3_6_stale_pdst = _RANDOM[11'h55B][10:4];	// rob.scala:310:28
        rob_uop_3_6_is_fencei = _RANDOM[11'h55D][22];	// rob.scala:310:28
        rob_uop_3_6_uses_ldq = _RANDOM[11'h55D][24];	// rob.scala:310:28
        rob_uop_3_6_uses_stq = _RANDOM[11'h55D][25];	// rob.scala:310:28
        rob_uop_3_6_is_sys_pc2epc = _RANDOM[11'h55D][26];	// rob.scala:310:28
        rob_uop_3_6_flush_on_commit = _RANDOM[11'h55D][28];	// rob.scala:310:28
        rob_uop_3_6_ldst = {_RANDOM[11'h55D][31:30], _RANDOM[11'h55E][3:0]};	// rob.scala:310:28
        rob_uop_3_6_ldst_val = _RANDOM[11'h55E][22];	// rob.scala:310:28
        rob_uop_3_6_dst_rtype = _RANDOM[11'h55E][24:23];	// rob.scala:310:28
        rob_uop_3_6_fp_val = _RANDOM[11'h55E][30];	// rob.scala:310:28
        rob_uop_3_7_uopc = _RANDOM[11'h55F][15:9];	// rob.scala:310:28
        rob_uop_3_7_is_rvc = _RANDOM[11'h561][16];	// rob.scala:310:28
        rob_uop_3_7_br_mask = _RANDOM[11'h564][24:5];	// rob.scala:310:28
        rob_uop_3_7_ftq_idx = {_RANDOM[11'h564][31:30], _RANDOM[11'h565][3:0]};	// rob.scala:310:28
        rob_uop_3_7_edge_inst = _RANDOM[11'h565][4];	// rob.scala:310:28
        rob_uop_3_7_pc_lob = _RANDOM[11'h565][10:5];	// rob.scala:310:28
        rob_uop_3_7_pdst = {_RANDOM[11'h566][31], _RANDOM[11'h567][5:0]};	// rob.scala:310:28
        rob_uop_3_7_stale_pdst = _RANDOM[11'h568][11:5];	// rob.scala:310:28
        rob_uop_3_7_is_fencei = _RANDOM[11'h56A][23];	// rob.scala:310:28
        rob_uop_3_7_uses_ldq = _RANDOM[11'h56A][25];	// rob.scala:310:28
        rob_uop_3_7_uses_stq = _RANDOM[11'h56A][26];	// rob.scala:310:28
        rob_uop_3_7_is_sys_pc2epc = _RANDOM[11'h56A][27];	// rob.scala:310:28
        rob_uop_3_7_flush_on_commit = _RANDOM[11'h56A][29];	// rob.scala:310:28
        rob_uop_3_7_ldst = {_RANDOM[11'h56A][31], _RANDOM[11'h56B][4:0]};	// rob.scala:310:28
        rob_uop_3_7_ldst_val = _RANDOM[11'h56B][23];	// rob.scala:310:28
        rob_uop_3_7_dst_rtype = _RANDOM[11'h56B][25:24];	// rob.scala:310:28
        rob_uop_3_7_fp_val = _RANDOM[11'h56B][31];	// rob.scala:310:28
        rob_uop_3_8_uopc = _RANDOM[11'h56C][16:10];	// rob.scala:310:28
        rob_uop_3_8_is_rvc = _RANDOM[11'h56E][17];	// rob.scala:310:28
        rob_uop_3_8_br_mask = _RANDOM[11'h571][25:6];	// rob.scala:310:28
        rob_uop_3_8_ftq_idx = {_RANDOM[11'h571][31], _RANDOM[11'h572][4:0]};	// rob.scala:310:28
        rob_uop_3_8_edge_inst = _RANDOM[11'h572][5];	// rob.scala:310:28
        rob_uop_3_8_pc_lob = _RANDOM[11'h572][11:6];	// rob.scala:310:28
        rob_uop_3_8_pdst = _RANDOM[11'h574][6:0];	// rob.scala:310:28
        rob_uop_3_8_stale_pdst = _RANDOM[11'h575][12:6];	// rob.scala:310:28
        rob_uop_3_8_is_fencei = _RANDOM[11'h577][24];	// rob.scala:310:28
        rob_uop_3_8_uses_ldq = _RANDOM[11'h577][26];	// rob.scala:310:28
        rob_uop_3_8_uses_stq = _RANDOM[11'h577][27];	// rob.scala:310:28
        rob_uop_3_8_is_sys_pc2epc = _RANDOM[11'h577][28];	// rob.scala:310:28
        rob_uop_3_8_flush_on_commit = _RANDOM[11'h577][30];	// rob.scala:310:28
        rob_uop_3_8_ldst = _RANDOM[11'h578][5:0];	// rob.scala:310:28
        rob_uop_3_8_ldst_val = _RANDOM[11'h578][24];	// rob.scala:310:28
        rob_uop_3_8_dst_rtype = _RANDOM[11'h578][26:25];	// rob.scala:310:28
        rob_uop_3_8_fp_val = _RANDOM[11'h579][0];	// rob.scala:310:28
        rob_uop_3_9_uopc = _RANDOM[11'h579][17:11];	// rob.scala:310:28
        rob_uop_3_9_is_rvc = _RANDOM[11'h57B][18];	// rob.scala:310:28
        rob_uop_3_9_br_mask = _RANDOM[11'h57E][26:7];	// rob.scala:310:28
        rob_uop_3_9_ftq_idx = _RANDOM[11'h57F][5:0];	// rob.scala:310:28
        rob_uop_3_9_edge_inst = _RANDOM[11'h57F][6];	// rob.scala:310:28
        rob_uop_3_9_pc_lob = _RANDOM[11'h57F][12:7];	// rob.scala:310:28
        rob_uop_3_9_pdst = _RANDOM[11'h581][7:1];	// rob.scala:310:28
        rob_uop_3_9_stale_pdst = _RANDOM[11'h582][13:7];	// rob.scala:310:28
        rob_uop_3_9_is_fencei = _RANDOM[11'h584][25];	// rob.scala:310:28
        rob_uop_3_9_uses_ldq = _RANDOM[11'h584][27];	// rob.scala:310:28
        rob_uop_3_9_uses_stq = _RANDOM[11'h584][28];	// rob.scala:310:28
        rob_uop_3_9_is_sys_pc2epc = _RANDOM[11'h584][29];	// rob.scala:310:28
        rob_uop_3_9_flush_on_commit = _RANDOM[11'h584][31];	// rob.scala:310:28
        rob_uop_3_9_ldst = _RANDOM[11'h585][6:1];	// rob.scala:310:28
        rob_uop_3_9_ldst_val = _RANDOM[11'h585][25];	// rob.scala:310:28
        rob_uop_3_9_dst_rtype = _RANDOM[11'h585][27:26];	// rob.scala:310:28
        rob_uop_3_9_fp_val = _RANDOM[11'h586][1];	// rob.scala:310:28
        rob_uop_3_10_uopc = _RANDOM[11'h586][18:12];	// rob.scala:310:28
        rob_uop_3_10_is_rvc = _RANDOM[11'h588][19];	// rob.scala:310:28
        rob_uop_3_10_br_mask = _RANDOM[11'h58B][27:8];	// rob.scala:310:28
        rob_uop_3_10_ftq_idx = _RANDOM[11'h58C][6:1];	// rob.scala:310:28
        rob_uop_3_10_edge_inst = _RANDOM[11'h58C][7];	// rob.scala:310:28
        rob_uop_3_10_pc_lob = _RANDOM[11'h58C][13:8];	// rob.scala:310:28
        rob_uop_3_10_pdst = _RANDOM[11'h58E][8:2];	// rob.scala:310:28
        rob_uop_3_10_stale_pdst = _RANDOM[11'h58F][14:8];	// rob.scala:310:28
        rob_uop_3_10_is_fencei = _RANDOM[11'h591][26];	// rob.scala:310:28
        rob_uop_3_10_uses_ldq = _RANDOM[11'h591][28];	// rob.scala:310:28
        rob_uop_3_10_uses_stq = _RANDOM[11'h591][29];	// rob.scala:310:28
        rob_uop_3_10_is_sys_pc2epc = _RANDOM[11'h591][30];	// rob.scala:310:28
        rob_uop_3_10_flush_on_commit = _RANDOM[11'h592][0];	// rob.scala:310:28
        rob_uop_3_10_ldst = _RANDOM[11'h592][7:2];	// rob.scala:310:28
        rob_uop_3_10_ldst_val = _RANDOM[11'h592][26];	// rob.scala:310:28
        rob_uop_3_10_dst_rtype = _RANDOM[11'h592][28:27];	// rob.scala:310:28
        rob_uop_3_10_fp_val = _RANDOM[11'h593][2];	// rob.scala:310:28
        rob_uop_3_11_uopc = _RANDOM[11'h593][19:13];	// rob.scala:310:28
        rob_uop_3_11_is_rvc = _RANDOM[11'h595][20];	// rob.scala:310:28
        rob_uop_3_11_br_mask = _RANDOM[11'h598][28:9];	// rob.scala:310:28
        rob_uop_3_11_ftq_idx = _RANDOM[11'h599][7:2];	// rob.scala:310:28
        rob_uop_3_11_edge_inst = _RANDOM[11'h599][8];	// rob.scala:310:28
        rob_uop_3_11_pc_lob = _RANDOM[11'h599][14:9];	// rob.scala:310:28
        rob_uop_3_11_pdst = _RANDOM[11'h59B][9:3];	// rob.scala:310:28
        rob_uop_3_11_stale_pdst = _RANDOM[11'h59C][15:9];	// rob.scala:310:28
        rob_uop_3_11_is_fencei = _RANDOM[11'h59E][27];	// rob.scala:310:28
        rob_uop_3_11_uses_ldq = _RANDOM[11'h59E][29];	// rob.scala:310:28
        rob_uop_3_11_uses_stq = _RANDOM[11'h59E][30];	// rob.scala:310:28
        rob_uop_3_11_is_sys_pc2epc = _RANDOM[11'h59E][31];	// rob.scala:310:28
        rob_uop_3_11_flush_on_commit = _RANDOM[11'h59F][1];	// rob.scala:310:28
        rob_uop_3_11_ldst = _RANDOM[11'h59F][8:3];	// rob.scala:310:28
        rob_uop_3_11_ldst_val = _RANDOM[11'h59F][27];	// rob.scala:310:28
        rob_uop_3_11_dst_rtype = _RANDOM[11'h59F][29:28];	// rob.scala:310:28
        rob_uop_3_11_fp_val = _RANDOM[11'h5A0][3];	// rob.scala:310:28
        rob_uop_3_12_uopc = _RANDOM[11'h5A0][20:14];	// rob.scala:310:28
        rob_uop_3_12_is_rvc = _RANDOM[11'h5A2][21];	// rob.scala:310:28
        rob_uop_3_12_br_mask = _RANDOM[11'h5A5][29:10];	// rob.scala:310:28
        rob_uop_3_12_ftq_idx = _RANDOM[11'h5A6][8:3];	// rob.scala:310:28
        rob_uop_3_12_edge_inst = _RANDOM[11'h5A6][9];	// rob.scala:310:28
        rob_uop_3_12_pc_lob = _RANDOM[11'h5A6][15:10];	// rob.scala:310:28
        rob_uop_3_12_pdst = _RANDOM[11'h5A8][10:4];	// rob.scala:310:28
        rob_uop_3_12_stale_pdst = _RANDOM[11'h5A9][16:10];	// rob.scala:310:28
        rob_uop_3_12_is_fencei = _RANDOM[11'h5AB][28];	// rob.scala:310:28
        rob_uop_3_12_uses_ldq = _RANDOM[11'h5AB][30];	// rob.scala:310:28
        rob_uop_3_12_uses_stq = _RANDOM[11'h5AB][31];	// rob.scala:310:28
        rob_uop_3_12_is_sys_pc2epc = _RANDOM[11'h5AC][0];	// rob.scala:310:28
        rob_uop_3_12_flush_on_commit = _RANDOM[11'h5AC][2];	// rob.scala:310:28
        rob_uop_3_12_ldst = _RANDOM[11'h5AC][9:4];	// rob.scala:310:28
        rob_uop_3_12_ldst_val = _RANDOM[11'h5AC][28];	// rob.scala:310:28
        rob_uop_3_12_dst_rtype = _RANDOM[11'h5AC][30:29];	// rob.scala:310:28
        rob_uop_3_12_fp_val = _RANDOM[11'h5AD][4];	// rob.scala:310:28
        rob_uop_3_13_uopc = _RANDOM[11'h5AD][21:15];	// rob.scala:310:28
        rob_uop_3_13_is_rvc = _RANDOM[11'h5AF][22];	// rob.scala:310:28
        rob_uop_3_13_br_mask = _RANDOM[11'h5B2][30:11];	// rob.scala:310:28
        rob_uop_3_13_ftq_idx = _RANDOM[11'h5B3][9:4];	// rob.scala:310:28
        rob_uop_3_13_edge_inst = _RANDOM[11'h5B3][10];	// rob.scala:310:28
        rob_uop_3_13_pc_lob = _RANDOM[11'h5B3][16:11];	// rob.scala:310:28
        rob_uop_3_13_pdst = _RANDOM[11'h5B5][11:5];	// rob.scala:310:28
        rob_uop_3_13_stale_pdst = _RANDOM[11'h5B6][17:11];	// rob.scala:310:28
        rob_uop_3_13_is_fencei = _RANDOM[11'h5B8][29];	// rob.scala:310:28
        rob_uop_3_13_uses_ldq = _RANDOM[11'h5B8][31];	// rob.scala:310:28
        rob_uop_3_13_uses_stq = _RANDOM[11'h5B9][0];	// rob.scala:310:28
        rob_uop_3_13_is_sys_pc2epc = _RANDOM[11'h5B9][1];	// rob.scala:310:28
        rob_uop_3_13_flush_on_commit = _RANDOM[11'h5B9][3];	// rob.scala:310:28
        rob_uop_3_13_ldst = _RANDOM[11'h5B9][10:5];	// rob.scala:310:28
        rob_uop_3_13_ldst_val = _RANDOM[11'h5B9][29];	// rob.scala:310:28
        rob_uop_3_13_dst_rtype = _RANDOM[11'h5B9][31:30];	// rob.scala:310:28
        rob_uop_3_13_fp_val = _RANDOM[11'h5BA][5];	// rob.scala:310:28
        rob_uop_3_14_uopc = _RANDOM[11'h5BA][22:16];	// rob.scala:310:28
        rob_uop_3_14_is_rvc = _RANDOM[11'h5BC][23];	// rob.scala:310:28
        rob_uop_3_14_br_mask = _RANDOM[11'h5BF][31:12];	// rob.scala:310:28
        rob_uop_3_14_ftq_idx = _RANDOM[11'h5C0][10:5];	// rob.scala:310:28
        rob_uop_3_14_edge_inst = _RANDOM[11'h5C0][11];	// rob.scala:310:28
        rob_uop_3_14_pc_lob = _RANDOM[11'h5C0][17:12];	// rob.scala:310:28
        rob_uop_3_14_pdst = _RANDOM[11'h5C2][12:6];	// rob.scala:310:28
        rob_uop_3_14_stale_pdst = _RANDOM[11'h5C3][18:12];	// rob.scala:310:28
        rob_uop_3_14_is_fencei = _RANDOM[11'h5C5][30];	// rob.scala:310:28
        rob_uop_3_14_uses_ldq = _RANDOM[11'h5C6][0];	// rob.scala:310:28
        rob_uop_3_14_uses_stq = _RANDOM[11'h5C6][1];	// rob.scala:310:28
        rob_uop_3_14_is_sys_pc2epc = _RANDOM[11'h5C6][2];	// rob.scala:310:28
        rob_uop_3_14_flush_on_commit = _RANDOM[11'h5C6][4];	// rob.scala:310:28
        rob_uop_3_14_ldst = _RANDOM[11'h5C6][11:6];	// rob.scala:310:28
        rob_uop_3_14_ldst_val = _RANDOM[11'h5C6][30];	// rob.scala:310:28
        rob_uop_3_14_dst_rtype = {_RANDOM[11'h5C6][31], _RANDOM[11'h5C7][0]};	// rob.scala:310:28
        rob_uop_3_14_fp_val = _RANDOM[11'h5C7][6];	// rob.scala:310:28
        rob_uop_3_15_uopc = _RANDOM[11'h5C7][23:17];	// rob.scala:310:28
        rob_uop_3_15_is_rvc = _RANDOM[11'h5C9][24];	// rob.scala:310:28
        rob_uop_3_15_br_mask = {_RANDOM[11'h5CC][31:13], _RANDOM[11'h5CD][0]};	// rob.scala:310:28
        rob_uop_3_15_ftq_idx = _RANDOM[11'h5CD][11:6];	// rob.scala:310:28
        rob_uop_3_15_edge_inst = _RANDOM[11'h5CD][12];	// rob.scala:310:28
        rob_uop_3_15_pc_lob = _RANDOM[11'h5CD][18:13];	// rob.scala:310:28
        rob_uop_3_15_pdst = _RANDOM[11'h5CF][13:7];	// rob.scala:310:28
        rob_uop_3_15_stale_pdst = _RANDOM[11'h5D0][19:13];	// rob.scala:310:28
        rob_uop_3_15_is_fencei = _RANDOM[11'h5D2][31];	// rob.scala:310:28
        rob_uop_3_15_uses_ldq = _RANDOM[11'h5D3][1];	// rob.scala:310:28
        rob_uop_3_15_uses_stq = _RANDOM[11'h5D3][2];	// rob.scala:310:28
        rob_uop_3_15_is_sys_pc2epc = _RANDOM[11'h5D3][3];	// rob.scala:310:28
        rob_uop_3_15_flush_on_commit = _RANDOM[11'h5D3][5];	// rob.scala:310:28
        rob_uop_3_15_ldst = _RANDOM[11'h5D3][12:7];	// rob.scala:310:28
        rob_uop_3_15_ldst_val = _RANDOM[11'h5D3][31];	// rob.scala:310:28
        rob_uop_3_15_dst_rtype = _RANDOM[11'h5D4][1:0];	// rob.scala:310:28
        rob_uop_3_15_fp_val = _RANDOM[11'h5D4][7];	// rob.scala:310:28
        rob_uop_3_16_uopc = _RANDOM[11'h5D4][24:18];	// rob.scala:310:28
        rob_uop_3_16_is_rvc = _RANDOM[11'h5D6][25];	// rob.scala:310:28
        rob_uop_3_16_br_mask = {_RANDOM[11'h5D9][31:14], _RANDOM[11'h5DA][1:0]};	// rob.scala:310:28
        rob_uop_3_16_ftq_idx = _RANDOM[11'h5DA][12:7];	// rob.scala:310:28
        rob_uop_3_16_edge_inst = _RANDOM[11'h5DA][13];	// rob.scala:310:28
        rob_uop_3_16_pc_lob = _RANDOM[11'h5DA][19:14];	// rob.scala:310:28
        rob_uop_3_16_pdst = _RANDOM[11'h5DC][14:8];	// rob.scala:310:28
        rob_uop_3_16_stale_pdst = _RANDOM[11'h5DD][20:14];	// rob.scala:310:28
        rob_uop_3_16_is_fencei = _RANDOM[11'h5E0][0];	// rob.scala:310:28
        rob_uop_3_16_uses_ldq = _RANDOM[11'h5E0][2];	// rob.scala:310:28
        rob_uop_3_16_uses_stq = _RANDOM[11'h5E0][3];	// rob.scala:310:28
        rob_uop_3_16_is_sys_pc2epc = _RANDOM[11'h5E0][4];	// rob.scala:310:28
        rob_uop_3_16_flush_on_commit = _RANDOM[11'h5E0][6];	// rob.scala:310:28
        rob_uop_3_16_ldst = _RANDOM[11'h5E0][13:8];	// rob.scala:310:28
        rob_uop_3_16_ldst_val = _RANDOM[11'h5E1][0];	// rob.scala:310:28
        rob_uop_3_16_dst_rtype = _RANDOM[11'h5E1][2:1];	// rob.scala:310:28
        rob_uop_3_16_fp_val = _RANDOM[11'h5E1][8];	// rob.scala:310:28
        rob_uop_3_17_uopc = _RANDOM[11'h5E1][25:19];	// rob.scala:310:28
        rob_uop_3_17_is_rvc = _RANDOM[11'h5E3][26];	// rob.scala:310:28
        rob_uop_3_17_br_mask = {_RANDOM[11'h5E6][31:15], _RANDOM[11'h5E7][2:0]};	// rob.scala:310:28
        rob_uop_3_17_ftq_idx = _RANDOM[11'h5E7][13:8];	// rob.scala:310:28
        rob_uop_3_17_edge_inst = _RANDOM[11'h5E7][14];	// rob.scala:310:28
        rob_uop_3_17_pc_lob = _RANDOM[11'h5E7][20:15];	// rob.scala:310:28
        rob_uop_3_17_pdst = _RANDOM[11'h5E9][15:9];	// rob.scala:310:28
        rob_uop_3_17_stale_pdst = _RANDOM[11'h5EA][21:15];	// rob.scala:310:28
        rob_uop_3_17_is_fencei = _RANDOM[11'h5ED][1];	// rob.scala:310:28
        rob_uop_3_17_uses_ldq = _RANDOM[11'h5ED][3];	// rob.scala:310:28
        rob_uop_3_17_uses_stq = _RANDOM[11'h5ED][4];	// rob.scala:310:28
        rob_uop_3_17_is_sys_pc2epc = _RANDOM[11'h5ED][5];	// rob.scala:310:28
        rob_uop_3_17_flush_on_commit = _RANDOM[11'h5ED][7];	// rob.scala:310:28
        rob_uop_3_17_ldst = _RANDOM[11'h5ED][14:9];	// rob.scala:310:28
        rob_uop_3_17_ldst_val = _RANDOM[11'h5EE][1];	// rob.scala:310:28
        rob_uop_3_17_dst_rtype = _RANDOM[11'h5EE][3:2];	// rob.scala:310:28
        rob_uop_3_17_fp_val = _RANDOM[11'h5EE][9];	// rob.scala:310:28
        rob_uop_3_18_uopc = _RANDOM[11'h5EE][26:20];	// rob.scala:310:28
        rob_uop_3_18_is_rvc = _RANDOM[11'h5F0][27];	// rob.scala:310:28
        rob_uop_3_18_br_mask = {_RANDOM[11'h5F3][31:16], _RANDOM[11'h5F4][3:0]};	// rob.scala:310:28
        rob_uop_3_18_ftq_idx = _RANDOM[11'h5F4][14:9];	// rob.scala:310:28
        rob_uop_3_18_edge_inst = _RANDOM[11'h5F4][15];	// rob.scala:310:28
        rob_uop_3_18_pc_lob = _RANDOM[11'h5F4][21:16];	// rob.scala:310:28
        rob_uop_3_18_pdst = _RANDOM[11'h5F6][16:10];	// rob.scala:310:28
        rob_uop_3_18_stale_pdst = _RANDOM[11'h5F7][22:16];	// rob.scala:310:28
        rob_uop_3_18_is_fencei = _RANDOM[11'h5FA][2];	// rob.scala:310:28
        rob_uop_3_18_uses_ldq = _RANDOM[11'h5FA][4];	// rob.scala:310:28
        rob_uop_3_18_uses_stq = _RANDOM[11'h5FA][5];	// rob.scala:310:28
        rob_uop_3_18_is_sys_pc2epc = _RANDOM[11'h5FA][6];	// rob.scala:310:28
        rob_uop_3_18_flush_on_commit = _RANDOM[11'h5FA][8];	// rob.scala:310:28
        rob_uop_3_18_ldst = _RANDOM[11'h5FA][15:10];	// rob.scala:310:28
        rob_uop_3_18_ldst_val = _RANDOM[11'h5FB][2];	// rob.scala:310:28
        rob_uop_3_18_dst_rtype = _RANDOM[11'h5FB][4:3];	// rob.scala:310:28
        rob_uop_3_18_fp_val = _RANDOM[11'h5FB][10];	// rob.scala:310:28
        rob_uop_3_19_uopc = _RANDOM[11'h5FB][27:21];	// rob.scala:310:28
        rob_uop_3_19_is_rvc = _RANDOM[11'h5FD][28];	// rob.scala:310:28
        rob_uop_3_19_br_mask = {_RANDOM[11'h600][31:17], _RANDOM[11'h601][4:0]};	// rob.scala:310:28
        rob_uop_3_19_ftq_idx = _RANDOM[11'h601][15:10];	// rob.scala:310:28
        rob_uop_3_19_edge_inst = _RANDOM[11'h601][16];	// rob.scala:310:28
        rob_uop_3_19_pc_lob = _RANDOM[11'h601][22:17];	// rob.scala:310:28
        rob_uop_3_19_pdst = _RANDOM[11'h603][17:11];	// rob.scala:310:28
        rob_uop_3_19_stale_pdst = _RANDOM[11'h604][23:17];	// rob.scala:310:28
        rob_uop_3_19_is_fencei = _RANDOM[11'h607][3];	// rob.scala:310:28
        rob_uop_3_19_uses_ldq = _RANDOM[11'h607][5];	// rob.scala:310:28
        rob_uop_3_19_uses_stq = _RANDOM[11'h607][6];	// rob.scala:310:28
        rob_uop_3_19_is_sys_pc2epc = _RANDOM[11'h607][7];	// rob.scala:310:28
        rob_uop_3_19_flush_on_commit = _RANDOM[11'h607][9];	// rob.scala:310:28
        rob_uop_3_19_ldst = _RANDOM[11'h607][16:11];	// rob.scala:310:28
        rob_uop_3_19_ldst_val = _RANDOM[11'h608][3];	// rob.scala:310:28
        rob_uop_3_19_dst_rtype = _RANDOM[11'h608][5:4];	// rob.scala:310:28
        rob_uop_3_19_fp_val = _RANDOM[11'h608][11];	// rob.scala:310:28
        rob_uop_3_20_uopc = _RANDOM[11'h608][28:22];	// rob.scala:310:28
        rob_uop_3_20_is_rvc = _RANDOM[11'h60A][29];	// rob.scala:310:28
        rob_uop_3_20_br_mask = {_RANDOM[11'h60D][31:18], _RANDOM[11'h60E][5:0]};	// rob.scala:310:28
        rob_uop_3_20_ftq_idx = _RANDOM[11'h60E][16:11];	// rob.scala:310:28
        rob_uop_3_20_edge_inst = _RANDOM[11'h60E][17];	// rob.scala:310:28
        rob_uop_3_20_pc_lob = _RANDOM[11'h60E][23:18];	// rob.scala:310:28
        rob_uop_3_20_pdst = _RANDOM[11'h610][18:12];	// rob.scala:310:28
        rob_uop_3_20_stale_pdst = _RANDOM[11'h611][24:18];	// rob.scala:310:28
        rob_uop_3_20_is_fencei = _RANDOM[11'h614][4];	// rob.scala:310:28
        rob_uop_3_20_uses_ldq = _RANDOM[11'h614][6];	// rob.scala:310:28
        rob_uop_3_20_uses_stq = _RANDOM[11'h614][7];	// rob.scala:310:28
        rob_uop_3_20_is_sys_pc2epc = _RANDOM[11'h614][8];	// rob.scala:310:28
        rob_uop_3_20_flush_on_commit = _RANDOM[11'h614][10];	// rob.scala:310:28
        rob_uop_3_20_ldst = _RANDOM[11'h614][17:12];	// rob.scala:310:28
        rob_uop_3_20_ldst_val = _RANDOM[11'h615][4];	// rob.scala:310:28
        rob_uop_3_20_dst_rtype = _RANDOM[11'h615][6:5];	// rob.scala:310:28
        rob_uop_3_20_fp_val = _RANDOM[11'h615][12];	// rob.scala:310:28
        rob_uop_3_21_uopc = _RANDOM[11'h615][29:23];	// rob.scala:310:28
        rob_uop_3_21_is_rvc = _RANDOM[11'h617][30];	// rob.scala:310:28
        rob_uop_3_21_br_mask = {_RANDOM[11'h61A][31:19], _RANDOM[11'h61B][6:0]};	// rob.scala:310:28
        rob_uop_3_21_ftq_idx = _RANDOM[11'h61B][17:12];	// rob.scala:310:28
        rob_uop_3_21_edge_inst = _RANDOM[11'h61B][18];	// rob.scala:310:28
        rob_uop_3_21_pc_lob = _RANDOM[11'h61B][24:19];	// rob.scala:310:28
        rob_uop_3_21_pdst = _RANDOM[11'h61D][19:13];	// rob.scala:310:28
        rob_uop_3_21_stale_pdst = _RANDOM[11'h61E][25:19];	// rob.scala:310:28
        rob_uop_3_21_is_fencei = _RANDOM[11'h621][5];	// rob.scala:310:28
        rob_uop_3_21_uses_ldq = _RANDOM[11'h621][7];	// rob.scala:310:28
        rob_uop_3_21_uses_stq = _RANDOM[11'h621][8];	// rob.scala:310:28
        rob_uop_3_21_is_sys_pc2epc = _RANDOM[11'h621][9];	// rob.scala:310:28
        rob_uop_3_21_flush_on_commit = _RANDOM[11'h621][11];	// rob.scala:310:28
        rob_uop_3_21_ldst = _RANDOM[11'h621][18:13];	// rob.scala:310:28
        rob_uop_3_21_ldst_val = _RANDOM[11'h622][5];	// rob.scala:310:28
        rob_uop_3_21_dst_rtype = _RANDOM[11'h622][7:6];	// rob.scala:310:28
        rob_uop_3_21_fp_val = _RANDOM[11'h622][13];	// rob.scala:310:28
        rob_uop_3_22_uopc = _RANDOM[11'h622][30:24];	// rob.scala:310:28
        rob_uop_3_22_is_rvc = _RANDOM[11'h624][31];	// rob.scala:310:28
        rob_uop_3_22_br_mask = {_RANDOM[11'h627][31:20], _RANDOM[11'h628][7:0]};	// rob.scala:310:28
        rob_uop_3_22_ftq_idx = _RANDOM[11'h628][18:13];	// rob.scala:310:28
        rob_uop_3_22_edge_inst = _RANDOM[11'h628][19];	// rob.scala:310:28
        rob_uop_3_22_pc_lob = _RANDOM[11'h628][25:20];	// rob.scala:310:28
        rob_uop_3_22_pdst = _RANDOM[11'h62A][20:14];	// rob.scala:310:28
        rob_uop_3_22_stale_pdst = _RANDOM[11'h62B][26:20];	// rob.scala:310:28
        rob_uop_3_22_is_fencei = _RANDOM[11'h62E][6];	// rob.scala:310:28
        rob_uop_3_22_uses_ldq = _RANDOM[11'h62E][8];	// rob.scala:310:28
        rob_uop_3_22_uses_stq = _RANDOM[11'h62E][9];	// rob.scala:310:28
        rob_uop_3_22_is_sys_pc2epc = _RANDOM[11'h62E][10];	// rob.scala:310:28
        rob_uop_3_22_flush_on_commit = _RANDOM[11'h62E][12];	// rob.scala:310:28
        rob_uop_3_22_ldst = _RANDOM[11'h62E][19:14];	// rob.scala:310:28
        rob_uop_3_22_ldst_val = _RANDOM[11'h62F][6];	// rob.scala:310:28
        rob_uop_3_22_dst_rtype = _RANDOM[11'h62F][8:7];	// rob.scala:310:28
        rob_uop_3_22_fp_val = _RANDOM[11'h62F][14];	// rob.scala:310:28
        rob_uop_3_23_uopc = _RANDOM[11'h62F][31:25];	// rob.scala:310:28
        rob_uop_3_23_is_rvc = _RANDOM[11'h632][0];	// rob.scala:310:28
        rob_uop_3_23_br_mask = {_RANDOM[11'h634][31:21], _RANDOM[11'h635][8:0]};	// rob.scala:310:28
        rob_uop_3_23_ftq_idx = _RANDOM[11'h635][19:14];	// rob.scala:310:28
        rob_uop_3_23_edge_inst = _RANDOM[11'h635][20];	// rob.scala:310:28
        rob_uop_3_23_pc_lob = _RANDOM[11'h635][26:21];	// rob.scala:310:28
        rob_uop_3_23_pdst = _RANDOM[11'h637][21:15];	// rob.scala:310:28
        rob_uop_3_23_stale_pdst = _RANDOM[11'h638][27:21];	// rob.scala:310:28
        rob_uop_3_23_is_fencei = _RANDOM[11'h63B][7];	// rob.scala:310:28
        rob_uop_3_23_uses_ldq = _RANDOM[11'h63B][9];	// rob.scala:310:28
        rob_uop_3_23_uses_stq = _RANDOM[11'h63B][10];	// rob.scala:310:28
        rob_uop_3_23_is_sys_pc2epc = _RANDOM[11'h63B][11];	// rob.scala:310:28
        rob_uop_3_23_flush_on_commit = _RANDOM[11'h63B][13];	// rob.scala:310:28
        rob_uop_3_23_ldst = _RANDOM[11'h63B][20:15];	// rob.scala:310:28
        rob_uop_3_23_ldst_val = _RANDOM[11'h63C][7];	// rob.scala:310:28
        rob_uop_3_23_dst_rtype = _RANDOM[11'h63C][9:8];	// rob.scala:310:28
        rob_uop_3_23_fp_val = _RANDOM[11'h63C][15];	// rob.scala:310:28
        rob_uop_3_24_uopc = {_RANDOM[11'h63C][31:26], _RANDOM[11'h63D][0]};	// rob.scala:310:28
        rob_uop_3_24_is_rvc = _RANDOM[11'h63F][1];	// rob.scala:310:28
        rob_uop_3_24_br_mask = {_RANDOM[11'h641][31:22], _RANDOM[11'h642][9:0]};	// rob.scala:310:28
        rob_uop_3_24_ftq_idx = _RANDOM[11'h642][20:15];	// rob.scala:310:28
        rob_uop_3_24_edge_inst = _RANDOM[11'h642][21];	// rob.scala:310:28
        rob_uop_3_24_pc_lob = _RANDOM[11'h642][27:22];	// rob.scala:310:28
        rob_uop_3_24_pdst = _RANDOM[11'h644][22:16];	// rob.scala:310:28
        rob_uop_3_24_stale_pdst = _RANDOM[11'h645][28:22];	// rob.scala:310:28
        rob_uop_3_24_is_fencei = _RANDOM[11'h648][8];	// rob.scala:310:28
        rob_uop_3_24_uses_ldq = _RANDOM[11'h648][10];	// rob.scala:310:28
        rob_uop_3_24_uses_stq = _RANDOM[11'h648][11];	// rob.scala:310:28
        rob_uop_3_24_is_sys_pc2epc = _RANDOM[11'h648][12];	// rob.scala:310:28
        rob_uop_3_24_flush_on_commit = _RANDOM[11'h648][14];	// rob.scala:310:28
        rob_uop_3_24_ldst = _RANDOM[11'h648][21:16];	// rob.scala:310:28
        rob_uop_3_24_ldst_val = _RANDOM[11'h649][8];	// rob.scala:310:28
        rob_uop_3_24_dst_rtype = _RANDOM[11'h649][10:9];	// rob.scala:310:28
        rob_uop_3_24_fp_val = _RANDOM[11'h649][16];	// rob.scala:310:28
        rob_uop_3_25_uopc = {_RANDOM[11'h649][31:27], _RANDOM[11'h64A][1:0]};	// rob.scala:310:28
        rob_uop_3_25_is_rvc = _RANDOM[11'h64C][2];	// rob.scala:310:28
        rob_uop_3_25_br_mask = {_RANDOM[11'h64E][31:23], _RANDOM[11'h64F][10:0]};	// rob.scala:310:28
        rob_uop_3_25_ftq_idx = _RANDOM[11'h64F][21:16];	// rob.scala:310:28
        rob_uop_3_25_edge_inst = _RANDOM[11'h64F][22];	// rob.scala:310:28
        rob_uop_3_25_pc_lob = _RANDOM[11'h64F][28:23];	// rob.scala:310:28
        rob_uop_3_25_pdst = _RANDOM[11'h651][23:17];	// rob.scala:310:28
        rob_uop_3_25_stale_pdst = _RANDOM[11'h652][29:23];	// rob.scala:310:28
        rob_uop_3_25_is_fencei = _RANDOM[11'h655][9];	// rob.scala:310:28
        rob_uop_3_25_uses_ldq = _RANDOM[11'h655][11];	// rob.scala:310:28
        rob_uop_3_25_uses_stq = _RANDOM[11'h655][12];	// rob.scala:310:28
        rob_uop_3_25_is_sys_pc2epc = _RANDOM[11'h655][13];	// rob.scala:310:28
        rob_uop_3_25_flush_on_commit = _RANDOM[11'h655][15];	// rob.scala:310:28
        rob_uop_3_25_ldst = _RANDOM[11'h655][22:17];	// rob.scala:310:28
        rob_uop_3_25_ldst_val = _RANDOM[11'h656][9];	// rob.scala:310:28
        rob_uop_3_25_dst_rtype = _RANDOM[11'h656][11:10];	// rob.scala:310:28
        rob_uop_3_25_fp_val = _RANDOM[11'h656][17];	// rob.scala:310:28
        rob_uop_3_26_uopc = {_RANDOM[11'h656][31:28], _RANDOM[11'h657][2:0]};	// rob.scala:310:28
        rob_uop_3_26_is_rvc = _RANDOM[11'h659][3];	// rob.scala:310:28
        rob_uop_3_26_br_mask = {_RANDOM[11'h65B][31:24], _RANDOM[11'h65C][11:0]};	// rob.scala:310:28
        rob_uop_3_26_ftq_idx = _RANDOM[11'h65C][22:17];	// rob.scala:310:28
        rob_uop_3_26_edge_inst = _RANDOM[11'h65C][23];	// rob.scala:310:28
        rob_uop_3_26_pc_lob = _RANDOM[11'h65C][29:24];	// rob.scala:310:28
        rob_uop_3_26_pdst = _RANDOM[11'h65E][24:18];	// rob.scala:310:28
        rob_uop_3_26_stale_pdst = _RANDOM[11'h65F][30:24];	// rob.scala:310:28
        rob_uop_3_26_is_fencei = _RANDOM[11'h662][10];	// rob.scala:310:28
        rob_uop_3_26_uses_ldq = _RANDOM[11'h662][12];	// rob.scala:310:28
        rob_uop_3_26_uses_stq = _RANDOM[11'h662][13];	// rob.scala:310:28
        rob_uop_3_26_is_sys_pc2epc = _RANDOM[11'h662][14];	// rob.scala:310:28
        rob_uop_3_26_flush_on_commit = _RANDOM[11'h662][16];	// rob.scala:310:28
        rob_uop_3_26_ldst = _RANDOM[11'h662][23:18];	// rob.scala:310:28
        rob_uop_3_26_ldst_val = _RANDOM[11'h663][10];	// rob.scala:310:28
        rob_uop_3_26_dst_rtype = _RANDOM[11'h663][12:11];	// rob.scala:310:28
        rob_uop_3_26_fp_val = _RANDOM[11'h663][18];	// rob.scala:310:28
        rob_uop_3_27_uopc = {_RANDOM[11'h663][31:29], _RANDOM[11'h664][3:0]};	// rob.scala:310:28
        rob_uop_3_27_is_rvc = _RANDOM[11'h666][4];	// rob.scala:310:28
        rob_uop_3_27_br_mask = {_RANDOM[11'h668][31:25], _RANDOM[11'h669][12:0]};	// rob.scala:310:28
        rob_uop_3_27_ftq_idx = _RANDOM[11'h669][23:18];	// rob.scala:310:28
        rob_uop_3_27_edge_inst = _RANDOM[11'h669][24];	// rob.scala:310:28
        rob_uop_3_27_pc_lob = _RANDOM[11'h669][30:25];	// rob.scala:310:28
        rob_uop_3_27_pdst = _RANDOM[11'h66B][25:19];	// rob.scala:310:28
        rob_uop_3_27_stale_pdst = _RANDOM[11'h66C][31:25];	// rob.scala:310:28
        rob_uop_3_27_is_fencei = _RANDOM[11'h66F][11];	// rob.scala:310:28
        rob_uop_3_27_uses_ldq = _RANDOM[11'h66F][13];	// rob.scala:310:28
        rob_uop_3_27_uses_stq = _RANDOM[11'h66F][14];	// rob.scala:310:28
        rob_uop_3_27_is_sys_pc2epc = _RANDOM[11'h66F][15];	// rob.scala:310:28
        rob_uop_3_27_flush_on_commit = _RANDOM[11'h66F][17];	// rob.scala:310:28
        rob_uop_3_27_ldst = _RANDOM[11'h66F][24:19];	// rob.scala:310:28
        rob_uop_3_27_ldst_val = _RANDOM[11'h670][11];	// rob.scala:310:28
        rob_uop_3_27_dst_rtype = _RANDOM[11'h670][13:12];	// rob.scala:310:28
        rob_uop_3_27_fp_val = _RANDOM[11'h670][19];	// rob.scala:310:28
        rob_uop_3_28_uopc = {_RANDOM[11'h670][31:30], _RANDOM[11'h671][4:0]};	// rob.scala:310:28
        rob_uop_3_28_is_rvc = _RANDOM[11'h673][5];	// rob.scala:310:28
        rob_uop_3_28_br_mask = {_RANDOM[11'h675][31:26], _RANDOM[11'h676][13:0]};	// rob.scala:310:28
        rob_uop_3_28_ftq_idx = _RANDOM[11'h676][24:19];	// rob.scala:310:28
        rob_uop_3_28_edge_inst = _RANDOM[11'h676][25];	// rob.scala:310:28
        rob_uop_3_28_pc_lob = _RANDOM[11'h676][31:26];	// rob.scala:310:28
        rob_uop_3_28_pdst = _RANDOM[11'h678][26:20];	// rob.scala:310:28
        rob_uop_3_28_stale_pdst = {_RANDOM[11'h679][31:26], _RANDOM[11'h67A][0]};	// rob.scala:310:28
        rob_uop_3_28_is_fencei = _RANDOM[11'h67C][12];	// rob.scala:310:28
        rob_uop_3_28_uses_ldq = _RANDOM[11'h67C][14];	// rob.scala:310:28
        rob_uop_3_28_uses_stq = _RANDOM[11'h67C][15];	// rob.scala:310:28
        rob_uop_3_28_is_sys_pc2epc = _RANDOM[11'h67C][16];	// rob.scala:310:28
        rob_uop_3_28_flush_on_commit = _RANDOM[11'h67C][18];	// rob.scala:310:28
        rob_uop_3_28_ldst = _RANDOM[11'h67C][25:20];	// rob.scala:310:28
        rob_uop_3_28_ldst_val = _RANDOM[11'h67D][12];	// rob.scala:310:28
        rob_uop_3_28_dst_rtype = _RANDOM[11'h67D][14:13];	// rob.scala:310:28
        rob_uop_3_28_fp_val = _RANDOM[11'h67D][20];	// rob.scala:310:28
        rob_uop_3_29_uopc = {_RANDOM[11'h67D][31], _RANDOM[11'h67E][5:0]};	// rob.scala:310:28
        rob_uop_3_29_is_rvc = _RANDOM[11'h680][6];	// rob.scala:310:28
        rob_uop_3_29_br_mask = {_RANDOM[11'h682][31:27], _RANDOM[11'h683][14:0]};	// rob.scala:310:28
        rob_uop_3_29_ftq_idx = _RANDOM[11'h683][25:20];	// rob.scala:310:28
        rob_uop_3_29_edge_inst = _RANDOM[11'h683][26];	// rob.scala:310:28
        rob_uop_3_29_pc_lob = {_RANDOM[11'h683][31:27], _RANDOM[11'h684][0]};	// rob.scala:310:28
        rob_uop_3_29_pdst = _RANDOM[11'h685][27:21];	// rob.scala:310:28
        rob_uop_3_29_stale_pdst = {_RANDOM[11'h686][31:27], _RANDOM[11'h687][1:0]};	// rob.scala:310:28
        rob_uop_3_29_is_fencei = _RANDOM[11'h689][13];	// rob.scala:310:28
        rob_uop_3_29_uses_ldq = _RANDOM[11'h689][15];	// rob.scala:310:28
        rob_uop_3_29_uses_stq = _RANDOM[11'h689][16];	// rob.scala:310:28
        rob_uop_3_29_is_sys_pc2epc = _RANDOM[11'h689][17];	// rob.scala:310:28
        rob_uop_3_29_flush_on_commit = _RANDOM[11'h689][19];	// rob.scala:310:28
        rob_uop_3_29_ldst = _RANDOM[11'h689][26:21];	// rob.scala:310:28
        rob_uop_3_29_ldst_val = _RANDOM[11'h68A][13];	// rob.scala:310:28
        rob_uop_3_29_dst_rtype = _RANDOM[11'h68A][15:14];	// rob.scala:310:28
        rob_uop_3_29_fp_val = _RANDOM[11'h68A][21];	// rob.scala:310:28
        rob_uop_3_30_uopc = _RANDOM[11'h68B][6:0];	// rob.scala:310:28
        rob_uop_3_30_is_rvc = _RANDOM[11'h68D][7];	// rob.scala:310:28
        rob_uop_3_30_br_mask = {_RANDOM[11'h68F][31:28], _RANDOM[11'h690][15:0]};	// rob.scala:310:28
        rob_uop_3_30_ftq_idx = _RANDOM[11'h690][26:21];	// rob.scala:310:28
        rob_uop_3_30_edge_inst = _RANDOM[11'h690][27];	// rob.scala:310:28
        rob_uop_3_30_pc_lob = {_RANDOM[11'h690][31:28], _RANDOM[11'h691][1:0]};	// rob.scala:310:28
        rob_uop_3_30_pdst = _RANDOM[11'h692][28:22];	// rob.scala:310:28
        rob_uop_3_30_stale_pdst = {_RANDOM[11'h693][31:28], _RANDOM[11'h694][2:0]};	// rob.scala:310:28
        rob_uop_3_30_is_fencei = _RANDOM[11'h696][14];	// rob.scala:310:28
        rob_uop_3_30_uses_ldq = _RANDOM[11'h696][16];	// rob.scala:310:28
        rob_uop_3_30_uses_stq = _RANDOM[11'h696][17];	// rob.scala:310:28
        rob_uop_3_30_is_sys_pc2epc = _RANDOM[11'h696][18];	// rob.scala:310:28
        rob_uop_3_30_flush_on_commit = _RANDOM[11'h696][20];	// rob.scala:310:28
        rob_uop_3_30_ldst = _RANDOM[11'h696][27:22];	// rob.scala:310:28
        rob_uop_3_30_ldst_val = _RANDOM[11'h697][14];	// rob.scala:310:28
        rob_uop_3_30_dst_rtype = _RANDOM[11'h697][16:15];	// rob.scala:310:28
        rob_uop_3_30_fp_val = _RANDOM[11'h697][22];	// rob.scala:310:28
        rob_uop_3_31_uopc = _RANDOM[11'h698][7:1];	// rob.scala:310:28
        rob_uop_3_31_is_rvc = _RANDOM[11'h69A][8];	// rob.scala:310:28
        rob_uop_3_31_br_mask = {_RANDOM[11'h69C][31:29], _RANDOM[11'h69D][16:0]};	// rob.scala:310:28
        rob_uop_3_31_ftq_idx = _RANDOM[11'h69D][27:22];	// rob.scala:310:28
        rob_uop_3_31_edge_inst = _RANDOM[11'h69D][28];	// rob.scala:310:28
        rob_uop_3_31_pc_lob = {_RANDOM[11'h69D][31:29], _RANDOM[11'h69E][2:0]};	// rob.scala:310:28
        rob_uop_3_31_pdst = _RANDOM[11'h69F][29:23];	// rob.scala:310:28
        rob_uop_3_31_stale_pdst = {_RANDOM[11'h6A0][31:29], _RANDOM[11'h6A1][3:0]};	// rob.scala:310:28
        rob_uop_3_31_is_fencei = _RANDOM[11'h6A3][15];	// rob.scala:310:28
        rob_uop_3_31_uses_ldq = _RANDOM[11'h6A3][17];	// rob.scala:310:28
        rob_uop_3_31_uses_stq = _RANDOM[11'h6A3][18];	// rob.scala:310:28
        rob_uop_3_31_is_sys_pc2epc = _RANDOM[11'h6A3][19];	// rob.scala:310:28
        rob_uop_3_31_flush_on_commit = _RANDOM[11'h6A3][21];	// rob.scala:310:28
        rob_uop_3_31_ldst = _RANDOM[11'h6A3][28:23];	// rob.scala:310:28
        rob_uop_3_31_ldst_val = _RANDOM[11'h6A4][15];	// rob.scala:310:28
        rob_uop_3_31_dst_rtype = _RANDOM[11'h6A4][17:16];	// rob.scala:310:28
        rob_uop_3_31_fp_val = _RANDOM[11'h6A4][23];	// rob.scala:310:28
        rob_exception_3_0 = _RANDOM[11'h6A5][2];	// rob.scala:311:28
        rob_exception_3_1 = _RANDOM[11'h6A5][3];	// rob.scala:311:28
        rob_exception_3_2 = _RANDOM[11'h6A5][4];	// rob.scala:311:28
        rob_exception_3_3 = _RANDOM[11'h6A5][5];	// rob.scala:311:28
        rob_exception_3_4 = _RANDOM[11'h6A5][6];	// rob.scala:311:28
        rob_exception_3_5 = _RANDOM[11'h6A5][7];	// rob.scala:311:28
        rob_exception_3_6 = _RANDOM[11'h6A5][8];	// rob.scala:311:28
        rob_exception_3_7 = _RANDOM[11'h6A5][9];	// rob.scala:311:28
        rob_exception_3_8 = _RANDOM[11'h6A5][10];	// rob.scala:311:28
        rob_exception_3_9 = _RANDOM[11'h6A5][11];	// rob.scala:311:28
        rob_exception_3_10 = _RANDOM[11'h6A5][12];	// rob.scala:311:28
        rob_exception_3_11 = _RANDOM[11'h6A5][13];	// rob.scala:311:28
        rob_exception_3_12 = _RANDOM[11'h6A5][14];	// rob.scala:311:28
        rob_exception_3_13 = _RANDOM[11'h6A5][15];	// rob.scala:311:28
        rob_exception_3_14 = _RANDOM[11'h6A5][16];	// rob.scala:311:28
        rob_exception_3_15 = _RANDOM[11'h6A5][17];	// rob.scala:311:28
        rob_exception_3_16 = _RANDOM[11'h6A5][18];	// rob.scala:311:28
        rob_exception_3_17 = _RANDOM[11'h6A5][19];	// rob.scala:311:28
        rob_exception_3_18 = _RANDOM[11'h6A5][20];	// rob.scala:311:28
        rob_exception_3_19 = _RANDOM[11'h6A5][21];	// rob.scala:311:28
        rob_exception_3_20 = _RANDOM[11'h6A5][22];	// rob.scala:311:28
        rob_exception_3_21 = _RANDOM[11'h6A5][23];	// rob.scala:311:28
        rob_exception_3_22 = _RANDOM[11'h6A5][24];	// rob.scala:311:28
        rob_exception_3_23 = _RANDOM[11'h6A5][25];	// rob.scala:311:28
        rob_exception_3_24 = _RANDOM[11'h6A5][26];	// rob.scala:311:28
        rob_exception_3_25 = _RANDOM[11'h6A5][27];	// rob.scala:311:28
        rob_exception_3_26 = _RANDOM[11'h6A5][28];	// rob.scala:311:28
        rob_exception_3_27 = _RANDOM[11'h6A5][29];	// rob.scala:311:28
        rob_exception_3_28 = _RANDOM[11'h6A5][30];	// rob.scala:311:28
        rob_exception_3_29 = _RANDOM[11'h6A5][31];	// rob.scala:311:28
        rob_exception_3_30 = _RANDOM[11'h6A6][0];	// rob.scala:311:28
        rob_exception_3_31 = _RANDOM[11'h6A6][1];	// rob.scala:311:28
        rob_predicated_3_0 = _RANDOM[11'h6A6][2];	// rob.scala:311:28, :312:29
        rob_predicated_3_1 = _RANDOM[11'h6A6][3];	// rob.scala:311:28, :312:29
        rob_predicated_3_2 = _RANDOM[11'h6A6][4];	// rob.scala:311:28, :312:29
        rob_predicated_3_3 = _RANDOM[11'h6A6][5];	// rob.scala:311:28, :312:29
        rob_predicated_3_4 = _RANDOM[11'h6A6][6];	// rob.scala:311:28, :312:29
        rob_predicated_3_5 = _RANDOM[11'h6A6][7];	// rob.scala:311:28, :312:29
        rob_predicated_3_6 = _RANDOM[11'h6A6][8];	// rob.scala:311:28, :312:29
        rob_predicated_3_7 = _RANDOM[11'h6A6][9];	// rob.scala:311:28, :312:29
        rob_predicated_3_8 = _RANDOM[11'h6A6][10];	// rob.scala:311:28, :312:29
        rob_predicated_3_9 = _RANDOM[11'h6A6][11];	// rob.scala:311:28, :312:29
        rob_predicated_3_10 = _RANDOM[11'h6A6][12];	// rob.scala:311:28, :312:29
        rob_predicated_3_11 = _RANDOM[11'h6A6][13];	// rob.scala:311:28, :312:29
        rob_predicated_3_12 = _RANDOM[11'h6A6][14];	// rob.scala:311:28, :312:29
        rob_predicated_3_13 = _RANDOM[11'h6A6][15];	// rob.scala:311:28, :312:29
        rob_predicated_3_14 = _RANDOM[11'h6A6][16];	// rob.scala:311:28, :312:29
        rob_predicated_3_15 = _RANDOM[11'h6A6][17];	// rob.scala:311:28, :312:29
        rob_predicated_3_16 = _RANDOM[11'h6A6][18];	// rob.scala:311:28, :312:29
        rob_predicated_3_17 = _RANDOM[11'h6A6][19];	// rob.scala:311:28, :312:29
        rob_predicated_3_18 = _RANDOM[11'h6A6][20];	// rob.scala:311:28, :312:29
        rob_predicated_3_19 = _RANDOM[11'h6A6][21];	// rob.scala:311:28, :312:29
        rob_predicated_3_20 = _RANDOM[11'h6A6][22];	// rob.scala:311:28, :312:29
        rob_predicated_3_21 = _RANDOM[11'h6A6][23];	// rob.scala:311:28, :312:29
        rob_predicated_3_22 = _RANDOM[11'h6A6][24];	// rob.scala:311:28, :312:29
        rob_predicated_3_23 = _RANDOM[11'h6A6][25];	// rob.scala:311:28, :312:29
        rob_predicated_3_24 = _RANDOM[11'h6A6][26];	// rob.scala:311:28, :312:29
        rob_predicated_3_25 = _RANDOM[11'h6A6][27];	// rob.scala:311:28, :312:29
        rob_predicated_3_26 = _RANDOM[11'h6A6][28];	// rob.scala:311:28, :312:29
        rob_predicated_3_27 = _RANDOM[11'h6A6][29];	// rob.scala:311:28, :312:29
        rob_predicated_3_28 = _RANDOM[11'h6A6][30];	// rob.scala:311:28, :312:29
        rob_predicated_3_29 = _RANDOM[11'h6A6][31];	// rob.scala:311:28, :312:29
        rob_predicated_3_30 = _RANDOM[11'h6A7][0];	// rob.scala:312:29
        rob_predicated_3_31 = _RANDOM[11'h6A7][1];	// rob.scala:312:29
        block_commit_REG = _RANDOM[11'h6A7][2];	// rob.scala:312:29, :540:94
        block_commit_REG_1 = _RANDOM[11'h6A7][3];	// rob.scala:312:29, :540:131
        block_commit_REG_2 = _RANDOM[11'h6A7][4];	// rob.scala:312:29, :540:123
        r_partial_row = _RANDOM[11'h6A7][5];	// rob.scala:312:29, :677:30
        pnr_maybe_at_tail = _RANDOM[11'h6A7][6];	// rob.scala:312:29, :714:36
        REG = _RANDOM[11'h6A7][7];	// rob.scala:312:29, :808:30
        REG_1 = _RANDOM[11'h6A7][8];	// rob.scala:312:29, :808:22
        REG_2 = _RANDOM[11'h6A7][9];	// rob.scala:312:29, :824:22
        io_com_load_is_at_rob_head_REG = _RANDOM[11'h6A7][10];	// rob.scala:312:29, :865:40
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  rob_fflags_32x5 rob_fflags_ext (	// rob.scala:313:28
    .R0_addr (rob_head),	// rob.scala:224:29
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .W0_addr (io_fflags_3_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W0_en   (io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h0),	// rob.scala:221:26, :272:36, :304:53, :381:32
    .W0_clk  (clock),
    .W0_data (io_fflags_3_bits_flags),
    .W1_addr (io_fflags_2_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W1_en   (io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h0),	// rob.scala:221:26, :272:36, :304:53, :381:32
    .W1_clk  (clock),
    .W1_data (io_fflags_2_bits_flags),
    .W2_addr (io_fflags_0_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W2_en   (io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h0),	// rob.scala:221:26, :272:36, :304:53, :381:32
    .W2_clk  (clock),
    .W2_data (io_fflags_0_bits_flags),
    .W3_addr (rob_tail),	// rob.scala:228:29
    .W3_en   (io_enq_valids_0),
    .W3_clk  (clock),
    .W3_data (5'h0),	// rob.scala:236:31, :268:25
    .R0_data (_rob_fflags_ext_R0_data)
  );
  rob_fflags_32x5 rob_fflags_1_ext (	// rob.scala:313:28
    .R0_addr (rob_head),	// rob.scala:224:29
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .W0_addr (io_fflags_3_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W0_en   (io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h1),	// rob.scala:272:36, :304:53, :381:32, :540:33
    .W0_clk  (clock),
    .W0_data (io_fflags_3_bits_flags),
    .W1_addr (io_fflags_2_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W1_en   (io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h1),	// rob.scala:272:36, :304:53, :381:32, :540:33
    .W1_clk  (clock),
    .W1_data (io_fflags_2_bits_flags),
    .W2_addr (io_fflags_0_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W2_en   (io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h1),	// rob.scala:272:36, :304:53, :381:32, :540:33
    .W2_clk  (clock),
    .W2_data (io_fflags_0_bits_flags),
    .W3_addr (rob_tail),	// rob.scala:228:29
    .W3_en   (io_enq_valids_1),
    .W3_clk  (clock),
    .W3_data (5'h0),	// rob.scala:236:31, :268:25
    .R0_data (_rob_fflags_1_ext_R0_data)
  );
  rob_fflags_32x5 rob_fflags_2_ext (	// rob.scala:313:28
    .R0_addr (rob_head),	// rob.scala:224:29
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .W0_addr (io_fflags_3_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W0_en   (io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h2),	// rob.scala:236:31, :272:36, :304:53, :381:32
    .W0_clk  (clock),
    .W0_data (io_fflags_3_bits_flags),
    .W1_addr (io_fflags_2_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W1_en   (io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h2),	// rob.scala:236:31, :272:36, :304:53, :381:32
    .W1_clk  (clock),
    .W1_data (io_fflags_2_bits_flags),
    .W2_addr (io_fflags_0_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W2_en   (io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h2),	// rob.scala:236:31, :272:36, :304:53, :381:32
    .W2_clk  (clock),
    .W2_data (io_fflags_0_bits_flags),
    .W3_addr (rob_tail),	// rob.scala:228:29
    .W3_en   (io_enq_valids_2),
    .W3_clk  (clock),
    .W3_data (5'h0),	// rob.scala:236:31, :268:25
    .R0_data (_rob_fflags_2_ext_R0_data)
  );
  rob_fflags_32x5 rob_fflags_3_ext (	// rob.scala:313:28
    .R0_addr (rob_head),	// rob.scala:224:29
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .W0_addr (io_fflags_3_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W0_en   (io_fflags_3_valid & (&(io_fflags_3_bits_uop_rob_idx[1:0]))),	// rob.scala:272:36, :304:53, :381:32
    .W0_clk  (clock),
    .W0_data (io_fflags_3_bits_flags),
    .W1_addr (io_fflags_2_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W1_en   (io_fflags_2_valid & (&(io_fflags_2_bits_uop_rob_idx[1:0]))),	// rob.scala:272:36, :304:53, :381:32
    .W1_clk  (clock),
    .W1_data (io_fflags_2_bits_flags),
    .W2_addr (io_fflags_0_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W2_en   (io_fflags_0_valid & (&(io_fflags_0_bits_uop_rob_idx[1:0]))),	// rob.scala:272:36, :304:53, :381:32
    .W2_clk  (clock),
    .W2_data (io_fflags_0_bits_flags),
    .W3_addr (rob_tail),	// rob.scala:228:29
    .W3_en   (io_enq_valids_3),
    .W3_clk  (clock),
    .W3_data (5'h0),	// rob.scala:236:31, :268:25
    .R0_data (_rob_fflags_3_ext_R0_data)
  );
  assign io_rob_tail_idx = rob_tail_idx;	// Cat.scala:30:58
  assign io_rob_head_idx = rob_head_idx;	// Cat.scala:30:58
  assign io_commit_valids_0 = will_commit_0;	// rob.scala:547:70
  assign io_commit_valids_1 = will_commit_1;	// rob.scala:547:70
  assign io_commit_valids_2 = will_commit_2;	// rob.scala:547:70
  assign io_commit_valids_3 = will_commit_3;	// rob.scala:547:70
  assign io_commit_arch_valids_0 = will_commit_0 & ~_GEN_17[com_idx];	// rob.scala:236:20, :410:{48,51}, :547:70
  assign io_commit_arch_valids_1 = will_commit_1 & ~_GEN_52[com_idx];	// rob.scala:236:20, :410:{48,51}, :547:70
  assign io_commit_arch_valids_2 = will_commit_2 & ~_GEN_87[com_idx];	// rob.scala:236:20, :410:{48,51}, :547:70
  assign io_commit_arch_valids_3 = will_commit_3 & ~_GEN_122[com_idx];	// rob.scala:236:20, :410:{48,51}, :547:70
  assign io_commit_uops_0_ftq_idx = _GEN_20[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_pdst = _GEN_23[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_stale_pdst = _GEN_24[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_is_fencei = _GEN_25[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_uses_ldq = _GEN_26[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_uses_stq = _GEN_27[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_ldst = _GEN_30[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_ldst_val = _GEN_31[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_dst_rtype = _GEN_32[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_ftq_idx = _GEN_55[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_pdst = _GEN_58[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_stale_pdst = _GEN_59[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_is_fencei = _GEN_60[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_uses_ldq = _GEN_61[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_uses_stq = _GEN_62[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_ldst = _GEN_65[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_ldst_val = _GEN_66[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_dst_rtype = _GEN_67[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_ftq_idx = _GEN_90[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_pdst = _GEN_93[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_stale_pdst = _GEN_94[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_is_fencei = _GEN_95[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_uses_ldq = _GEN_96[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_uses_stq = _GEN_97[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_ldst = _GEN_100[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_ldst_val = _GEN_101[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_dst_rtype = _GEN_102[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_ftq_idx = _GEN_125[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_pdst = _GEN_128[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_stale_pdst = _GEN_129[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_is_fencei = _GEN_130[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_uses_ldq = _GEN_131[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_uses_stq = _GEN_132[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_ldst = _GEN_135[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_ldst_val = _GEN_136[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_3_dst_rtype = _GEN_137[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_fflags_valid =
    fflags_val_0 | fflags_val_1 | fflags_val_2 | fflags_val_3;	// rob.scala:602:32, :617:48
  assign io_commit_fflags_bits =
    (fflags_val_0 ? _rob_fflags_ext_R0_data : 5'h0)
    | (fflags_val_1 ? _rob_fflags_1_ext_R0_data : 5'h0)
    | (fflags_val_2 ? _rob_fflags_2_ext_R0_data : 5'h0)
    | (fflags_val_3 ? _rob_fflags_3_ext_R0_data : 5'h0);	// rob.scala:236:31, :268:25, :313:28, :602:32, :605:21, :618:44
  assign io_commit_rbk_valids_0 = _io_commit_rbk_valids_0_output;	// rob.scala:427:40
  assign io_commit_rbk_valids_1 = _io_commit_rbk_valids_1_output;	// rob.scala:427:40
  assign io_commit_rbk_valids_2 = _io_commit_rbk_valids_2_output;	// rob.scala:427:40
  assign io_commit_rbk_valids_3 = _io_commit_rbk_valids_3_output;	// rob.scala:427:40
  assign io_commit_rollback = _io_commit_rollback_T_3;	// rob.scala:236:31
  assign io_com_load_is_at_rob_head = io_com_load_is_at_rob_head_REG;	// rob.scala:865:40
  assign io_com_xcpt_valid = exception_thrown & _io_flush_bits_flush_typ_T;	// rob.scala:545:85, :556:50, :557:41
  assign io_com_xcpt_bits_ftq_idx = com_xcpt_uop_ftq_idx;	// Mux.scala:47:69
  assign io_com_xcpt_bits_edge_inst = com_xcpt_uop_edge_inst;	// Mux.scala:47:69
  assign io_com_xcpt_bits_pc_lob = com_xcpt_uop_pc_lob;	// Mux.scala:47:69
  assign io_com_xcpt_bits_cause = r_xcpt_uop_exc_cause;	// rob.scala:259:29
  assign io_com_xcpt_bits_badvaddr = {{24{r_xcpt_badvaddr[39]}}, r_xcpt_badvaddr};	// Bitwise.scala:72:12, Cat.scala:30:58, rob.scala:260:29, util.scala:261:46
  assign io_flush_valid = _io_flush_valid_output;	// rob.scala:573:36
  assign io_flush_bits_ftq_idx =
    exception_thrown
      ? com_xcpt_uop_ftq_idx
      : (flush_commit_mask_0 ? _GEN_20[com_idx] : 6'h0)
        | (flush_commit_mask_1 ? _GEN_55[com_idx] : 6'h0)
        | (flush_commit_mask_2 ? _GEN_90[com_idx] : 6'h0)
        | (flush_commit_mask_3 ? _GEN_125[com_idx] : 6'h0);	// Mux.scala:27:72, :47:69, rob.scala:236:20, :287:15, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_edge_inst =
    exception_thrown
      ? com_xcpt_uop_edge_inst
      : flush_commit_mask_0 & _GEN_21[com_idx] | flush_commit_mask_1 & _GEN_56[com_idx]
        | flush_commit_mask_2 & _GEN_91[com_idx] | flush_commit_mask_3
        & _GEN_126[com_idx];	// Mux.scala:27:72, :47:69, rob.scala:236:20, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_is_rvc =
    exception_thrown
      ? (rob_head_vals_0
           ? _GEN_19[com_idx]
           : rob_head_vals_1
               ? _GEN_54[com_idx]
               : rob_head_vals_2 ? _GEN_89[com_idx] : _GEN_124[com_idx])
      : flush_commit_mask_0 & _GEN_19[com_idx] | flush_commit_mask_1 & _GEN_54[com_idx]
        | flush_commit_mask_2 & _GEN_89[com_idx] | flush_commit_mask_3
        & _GEN_124[com_idx];	// Mux.scala:27:72, :47:69, rob.scala:236:20, :398:49, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_pc_lob =
    exception_thrown
      ? com_xcpt_uop_pc_lob
      : (flush_commit_mask_0 ? _GEN_22[com_idx] : 6'h0)
        | (flush_commit_mask_1 ? _GEN_57[com_idx] : 6'h0)
        | (flush_commit_mask_2 ? _GEN_92[com_idx] : 6'h0)
        | (flush_commit_mask_3 ? _GEN_127[com_idx] : 6'h0);	// Mux.scala:27:72, :47:69, rob.scala:236:20, :287:15, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_flush_typ =
    _io_flush_valid_output
      ? (flush_commit
         & (exception_thrown
              ? (rob_head_vals_0
                   ? _GEN_18[com_idx]
                   : rob_head_vals_1
                       ? _GEN_53[com_idx]
                       : rob_head_vals_2 ? _GEN_88[com_idx] : _GEN_123[com_idx])
              : (flush_commit_mask_0 ? _GEN_18[com_idx] : 7'h0)
                | (flush_commit_mask_1 ? _GEN_53[com_idx] : 7'h0)
                | (flush_commit_mask_2 ? _GEN_88[com_idx] : 7'h0)
                | (flush_commit_mask_3 ? _GEN_123[com_idx] : 7'h0)) == 7'h6A
           ? 3'h3
           : exception_thrown & _io_flush_bits_flush_typ_T
               ? 3'h1
               : exception_thrown
                 | (rob_head_vals_0 | rob_head_vals_1 | rob_head_vals_2 | rob_head_vals_3)
                 & (rob_head_vals_0
                      ? _GEN_28[com_idx]
                      : rob_head_vals_1
                          ? _GEN_63[com_idx]
                          : rob_head_vals_2 ? _GEN_98[com_idx] : _GEN_133[com_idx])
                   ? 3'h2
                   : 3'h4)
      : 3'h0;	// Mux.scala:27:72, :47:69, rob.scala:172:10, :173:10, :174:10, :175:10, :236:20, :287:15, :398:49, :411:25, :457:33, :545:85, :556:50, :562:{27,31}, :564:39, :571:75, :572:48, :573:36, :578:22, :587:66, :588:{62,80}
  assign io_empty = empty;	// rob.scala:788:41
  assign io_ready = _io_ready_T & ~full & ~r_xcpt_val;	// rob.scala:258:33, :425:47, :658:33, :716:33, :787:39, :794:56
  assign io_flush_frontend = r_xcpt_val;	// rob.scala:258:33
endmodule

