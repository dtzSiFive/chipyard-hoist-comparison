// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module IssueUnitCollapsing_5(
  input         clock,
                reset,
                io_dis_uops_0_valid,
  input  [6:0]  io_dis_uops_0_bits_uopc,
  input  [31:0] io_dis_uops_0_bits_inst,
                io_dis_uops_0_bits_debug_inst,
  input         io_dis_uops_0_bits_is_rvc,
  input  [39:0] io_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_dis_uops_0_bits_iq_type,
  input  [9:0]  io_dis_uops_0_bits_fu_code,
  input         io_dis_uops_0_bits_is_br,
                io_dis_uops_0_bits_is_jalr,
                io_dis_uops_0_bits_is_jal,
                io_dis_uops_0_bits_is_sfb,
  input  [15:0] io_dis_uops_0_bits_br_mask,
  input  [3:0]  io_dis_uops_0_bits_br_tag,
  input  [4:0]  io_dis_uops_0_bits_ftq_idx,
  input         io_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_dis_uops_0_bits_pc_lob,
  input         io_dis_uops_0_bits_taken,
  input  [19:0] io_dis_uops_0_bits_imm_packed,
  input  [11:0] io_dis_uops_0_bits_csr_addr,
  input  [6:0]  io_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_dis_uops_0_bits_ldq_idx,
                io_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_dis_uops_0_bits_pdst,
                io_dis_uops_0_bits_prs1,
                io_dis_uops_0_bits_prs2,
                io_dis_uops_0_bits_prs3,
  input         io_dis_uops_0_bits_prs1_busy,
                io_dis_uops_0_bits_prs2_busy,
  input  [6:0]  io_dis_uops_0_bits_stale_pdst,
  input         io_dis_uops_0_bits_exception,
  input  [63:0] io_dis_uops_0_bits_exc_cause,
  input         io_dis_uops_0_bits_bypassable,
  input  [4:0]  io_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_dis_uops_0_bits_mem_size,
  input         io_dis_uops_0_bits_mem_signed,
                io_dis_uops_0_bits_is_fence,
                io_dis_uops_0_bits_is_fencei,
                io_dis_uops_0_bits_is_amo,
                io_dis_uops_0_bits_uses_ldq,
                io_dis_uops_0_bits_uses_stq,
                io_dis_uops_0_bits_is_sys_pc2epc,
                io_dis_uops_0_bits_is_unique,
                io_dis_uops_0_bits_flush_on_commit,
                io_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_0_bits_ldst,
                io_dis_uops_0_bits_lrs1,
                io_dis_uops_0_bits_lrs2,
                io_dis_uops_0_bits_lrs3,
  input         io_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_dis_uops_0_bits_dst_rtype,
                io_dis_uops_0_bits_lrs1_rtype,
                io_dis_uops_0_bits_lrs2_rtype,
  input         io_dis_uops_0_bits_frs3_en,
                io_dis_uops_0_bits_fp_val,
                io_dis_uops_0_bits_fp_single,
                io_dis_uops_0_bits_xcpt_pf_if,
                io_dis_uops_0_bits_xcpt_ae_if,
                io_dis_uops_0_bits_xcpt_ma_if,
                io_dis_uops_0_bits_bp_debug_if,
                io_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_0_bits_debug_fsrc,
                io_dis_uops_0_bits_debug_tsrc,
  input         io_dis_uops_1_valid,
  input  [6:0]  io_dis_uops_1_bits_uopc,
  input  [31:0] io_dis_uops_1_bits_inst,
                io_dis_uops_1_bits_debug_inst,
  input         io_dis_uops_1_bits_is_rvc,
  input  [39:0] io_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_dis_uops_1_bits_iq_type,
  input  [9:0]  io_dis_uops_1_bits_fu_code,
  input         io_dis_uops_1_bits_is_br,
                io_dis_uops_1_bits_is_jalr,
                io_dis_uops_1_bits_is_jal,
                io_dis_uops_1_bits_is_sfb,
  input  [15:0] io_dis_uops_1_bits_br_mask,
  input  [3:0]  io_dis_uops_1_bits_br_tag,
  input  [4:0]  io_dis_uops_1_bits_ftq_idx,
  input         io_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_dis_uops_1_bits_pc_lob,
  input         io_dis_uops_1_bits_taken,
  input  [19:0] io_dis_uops_1_bits_imm_packed,
  input  [11:0] io_dis_uops_1_bits_csr_addr,
  input  [6:0]  io_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_dis_uops_1_bits_ldq_idx,
                io_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_dis_uops_1_bits_pdst,
                io_dis_uops_1_bits_prs1,
                io_dis_uops_1_bits_prs2,
                io_dis_uops_1_bits_prs3,
  input         io_dis_uops_1_bits_prs1_busy,
                io_dis_uops_1_bits_prs2_busy,
  input  [6:0]  io_dis_uops_1_bits_stale_pdst,
  input         io_dis_uops_1_bits_exception,
  input  [63:0] io_dis_uops_1_bits_exc_cause,
  input         io_dis_uops_1_bits_bypassable,
  input  [4:0]  io_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_dis_uops_1_bits_mem_size,
  input         io_dis_uops_1_bits_mem_signed,
                io_dis_uops_1_bits_is_fence,
                io_dis_uops_1_bits_is_fencei,
                io_dis_uops_1_bits_is_amo,
                io_dis_uops_1_bits_uses_ldq,
                io_dis_uops_1_bits_uses_stq,
                io_dis_uops_1_bits_is_sys_pc2epc,
                io_dis_uops_1_bits_is_unique,
                io_dis_uops_1_bits_flush_on_commit,
                io_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_1_bits_ldst,
                io_dis_uops_1_bits_lrs1,
                io_dis_uops_1_bits_lrs2,
                io_dis_uops_1_bits_lrs3,
  input         io_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_dis_uops_1_bits_dst_rtype,
                io_dis_uops_1_bits_lrs1_rtype,
                io_dis_uops_1_bits_lrs2_rtype,
  input         io_dis_uops_1_bits_frs3_en,
                io_dis_uops_1_bits_fp_val,
                io_dis_uops_1_bits_fp_single,
                io_dis_uops_1_bits_xcpt_pf_if,
                io_dis_uops_1_bits_xcpt_ae_if,
                io_dis_uops_1_bits_xcpt_ma_if,
                io_dis_uops_1_bits_bp_debug_if,
                io_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_1_bits_debug_fsrc,
                io_dis_uops_1_bits_debug_tsrc,
  input         io_dis_uops_2_valid,
  input  [6:0]  io_dis_uops_2_bits_uopc,
  input  [31:0] io_dis_uops_2_bits_inst,
                io_dis_uops_2_bits_debug_inst,
  input         io_dis_uops_2_bits_is_rvc,
  input  [39:0] io_dis_uops_2_bits_debug_pc,
  input  [2:0]  io_dis_uops_2_bits_iq_type,
  input  [9:0]  io_dis_uops_2_bits_fu_code,
  input         io_dis_uops_2_bits_is_br,
                io_dis_uops_2_bits_is_jalr,
                io_dis_uops_2_bits_is_jal,
                io_dis_uops_2_bits_is_sfb,
  input  [15:0] io_dis_uops_2_bits_br_mask,
  input  [3:0]  io_dis_uops_2_bits_br_tag,
  input  [4:0]  io_dis_uops_2_bits_ftq_idx,
  input         io_dis_uops_2_bits_edge_inst,
  input  [5:0]  io_dis_uops_2_bits_pc_lob,
  input         io_dis_uops_2_bits_taken,
  input  [19:0] io_dis_uops_2_bits_imm_packed,
  input  [11:0] io_dis_uops_2_bits_csr_addr,
  input  [6:0]  io_dis_uops_2_bits_rob_idx,
  input  [4:0]  io_dis_uops_2_bits_ldq_idx,
                io_dis_uops_2_bits_stq_idx,
  input  [1:0]  io_dis_uops_2_bits_rxq_idx,
  input  [6:0]  io_dis_uops_2_bits_pdst,
                io_dis_uops_2_bits_prs1,
                io_dis_uops_2_bits_prs2,
                io_dis_uops_2_bits_prs3,
  input         io_dis_uops_2_bits_prs1_busy,
                io_dis_uops_2_bits_prs2_busy,
  input  [6:0]  io_dis_uops_2_bits_stale_pdst,
  input         io_dis_uops_2_bits_exception,
  input  [63:0] io_dis_uops_2_bits_exc_cause,
  input         io_dis_uops_2_bits_bypassable,
  input  [4:0]  io_dis_uops_2_bits_mem_cmd,
  input  [1:0]  io_dis_uops_2_bits_mem_size,
  input         io_dis_uops_2_bits_mem_signed,
                io_dis_uops_2_bits_is_fence,
                io_dis_uops_2_bits_is_fencei,
                io_dis_uops_2_bits_is_amo,
                io_dis_uops_2_bits_uses_ldq,
                io_dis_uops_2_bits_uses_stq,
                io_dis_uops_2_bits_is_sys_pc2epc,
                io_dis_uops_2_bits_is_unique,
                io_dis_uops_2_bits_flush_on_commit,
                io_dis_uops_2_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_2_bits_ldst,
                io_dis_uops_2_bits_lrs1,
                io_dis_uops_2_bits_lrs2,
                io_dis_uops_2_bits_lrs3,
  input         io_dis_uops_2_bits_ldst_val,
  input  [1:0]  io_dis_uops_2_bits_dst_rtype,
                io_dis_uops_2_bits_lrs1_rtype,
                io_dis_uops_2_bits_lrs2_rtype,
  input         io_dis_uops_2_bits_frs3_en,
                io_dis_uops_2_bits_fp_val,
                io_dis_uops_2_bits_fp_single,
                io_dis_uops_2_bits_xcpt_pf_if,
                io_dis_uops_2_bits_xcpt_ae_if,
                io_dis_uops_2_bits_xcpt_ma_if,
                io_dis_uops_2_bits_bp_debug_if,
                io_dis_uops_2_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_2_bits_debug_fsrc,
                io_dis_uops_2_bits_debug_tsrc,
  input         io_wakeup_ports_0_valid,
  input  [6:0]  io_wakeup_ports_0_bits_pdst,
  input         io_wakeup_ports_1_valid,
  input  [6:0]  io_wakeup_ports_1_bits_pdst,
  input         io_wakeup_ports_2_valid,
  input  [6:0]  io_wakeup_ports_2_bits_pdst,
  input         io_wakeup_ports_3_valid,
  input  [6:0]  io_wakeup_ports_3_bits_pdst,
  input         io_wakeup_ports_4_valid,
  input  [6:0]  io_wakeup_ports_4_bits_pdst,
  input         io_wakeup_ports_5_valid,
  input  [6:0]  io_wakeup_ports_5_bits_pdst,
  input         io_wakeup_ports_6_valid,
  input  [6:0]  io_wakeup_ports_6_bits_pdst,
  input         io_spec_ld_wakeup_0_valid,
  input  [6:0]  io_spec_ld_wakeup_0_bits,
  input  [9:0]  io_fu_types_0,
                io_fu_types_1,
                io_fu_types_2,
  input  [15:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input         io_flush_pipeline,
                io_ld_miss,
  output        io_dis_uops_0_ready,
                io_dis_uops_1_ready,
                io_dis_uops_2_ready,
                io_iss_valids_0,
                io_iss_valids_1,
                io_iss_valids_2,
  output [6:0]  io_iss_uops_0_uopc,
  output        io_iss_uops_0_is_rvc,
  output [9:0]  io_iss_uops_0_fu_code,
  output        io_iss_uops_0_iw_p1_poisoned,
                io_iss_uops_0_iw_p2_poisoned,
                io_iss_uops_0_is_br,
                io_iss_uops_0_is_jalr,
                io_iss_uops_0_is_jal,
                io_iss_uops_0_is_sfb,
  output [15:0] io_iss_uops_0_br_mask,
  output [3:0]  io_iss_uops_0_br_tag,
  output [4:0]  io_iss_uops_0_ftq_idx,
  output        io_iss_uops_0_edge_inst,
  output [5:0]  io_iss_uops_0_pc_lob,
  output        io_iss_uops_0_taken,
  output [19:0] io_iss_uops_0_imm_packed,
  output [6:0]  io_iss_uops_0_rob_idx,
  output [4:0]  io_iss_uops_0_ldq_idx,
                io_iss_uops_0_stq_idx,
  output [6:0]  io_iss_uops_0_pdst,
                io_iss_uops_0_prs1,
                io_iss_uops_0_prs2,
  output        io_iss_uops_0_bypassable,
  output [4:0]  io_iss_uops_0_mem_cmd,
  output        io_iss_uops_0_is_amo,
                io_iss_uops_0_uses_stq,
                io_iss_uops_0_ldst_val,
  output [1:0]  io_iss_uops_0_dst_rtype,
                io_iss_uops_0_lrs1_rtype,
                io_iss_uops_0_lrs2_rtype,
  output [6:0]  io_iss_uops_1_uopc,
  output [31:0] io_iss_uops_1_inst,
                io_iss_uops_1_debug_inst,
  output        io_iss_uops_1_is_rvc,
  output [39:0] io_iss_uops_1_debug_pc,
  output [2:0]  io_iss_uops_1_iq_type,
  output [9:0]  io_iss_uops_1_fu_code,
  output [1:0]  io_iss_uops_1_iw_state,
  output        io_iss_uops_1_iw_p1_poisoned,
                io_iss_uops_1_iw_p2_poisoned,
                io_iss_uops_1_is_br,
                io_iss_uops_1_is_jalr,
                io_iss_uops_1_is_jal,
                io_iss_uops_1_is_sfb,
  output [15:0] io_iss_uops_1_br_mask,
  output [3:0]  io_iss_uops_1_br_tag,
  output [4:0]  io_iss_uops_1_ftq_idx,
  output        io_iss_uops_1_edge_inst,
  output [5:0]  io_iss_uops_1_pc_lob,
  output        io_iss_uops_1_taken,
  output [19:0] io_iss_uops_1_imm_packed,
  output [11:0] io_iss_uops_1_csr_addr,
  output [6:0]  io_iss_uops_1_rob_idx,
  output [4:0]  io_iss_uops_1_ldq_idx,
                io_iss_uops_1_stq_idx,
  output [1:0]  io_iss_uops_1_rxq_idx,
  output [6:0]  io_iss_uops_1_pdst,
                io_iss_uops_1_prs1,
                io_iss_uops_1_prs2,
                io_iss_uops_1_prs3,
  output [4:0]  io_iss_uops_1_ppred,
  output        io_iss_uops_1_prs1_busy,
                io_iss_uops_1_prs2_busy,
                io_iss_uops_1_prs3_busy,
                io_iss_uops_1_ppred_busy,
  output [6:0]  io_iss_uops_1_stale_pdst,
  output        io_iss_uops_1_exception,
  output [63:0] io_iss_uops_1_exc_cause,
  output        io_iss_uops_1_bypassable,
  output [4:0]  io_iss_uops_1_mem_cmd,
  output [1:0]  io_iss_uops_1_mem_size,
  output        io_iss_uops_1_mem_signed,
                io_iss_uops_1_is_fence,
                io_iss_uops_1_is_fencei,
                io_iss_uops_1_is_amo,
                io_iss_uops_1_uses_ldq,
                io_iss_uops_1_uses_stq,
                io_iss_uops_1_is_sys_pc2epc,
                io_iss_uops_1_is_unique,
                io_iss_uops_1_flush_on_commit,
                io_iss_uops_1_ldst_is_rs1,
  output [5:0]  io_iss_uops_1_ldst,
                io_iss_uops_1_lrs1,
                io_iss_uops_1_lrs2,
                io_iss_uops_1_lrs3,
  output        io_iss_uops_1_ldst_val,
  output [1:0]  io_iss_uops_1_dst_rtype,
                io_iss_uops_1_lrs1_rtype,
                io_iss_uops_1_lrs2_rtype,
  output        io_iss_uops_1_frs3_en,
                io_iss_uops_1_fp_val,
                io_iss_uops_1_fp_single,
                io_iss_uops_1_xcpt_pf_if,
                io_iss_uops_1_xcpt_ae_if,
                io_iss_uops_1_xcpt_ma_if,
                io_iss_uops_1_bp_debug_if,
                io_iss_uops_1_bp_xcpt_if,
  output [1:0]  io_iss_uops_1_debug_fsrc,
                io_iss_uops_1_debug_tsrc,
  output [6:0]  io_iss_uops_2_uopc,
  output        io_iss_uops_2_is_rvc,
  output [9:0]  io_iss_uops_2_fu_code,
  output        io_iss_uops_2_iw_p1_poisoned,
                io_iss_uops_2_iw_p2_poisoned,
                io_iss_uops_2_is_br,
                io_iss_uops_2_is_jalr,
                io_iss_uops_2_is_jal,
                io_iss_uops_2_is_sfb,
  output [15:0] io_iss_uops_2_br_mask,
  output [3:0]  io_iss_uops_2_br_tag,
  output [4:0]  io_iss_uops_2_ftq_idx,
  output        io_iss_uops_2_edge_inst,
  output [5:0]  io_iss_uops_2_pc_lob,
  output        io_iss_uops_2_taken,
  output [19:0] io_iss_uops_2_imm_packed,
  output [6:0]  io_iss_uops_2_rob_idx,
  output [4:0]  io_iss_uops_2_ldq_idx,
                io_iss_uops_2_stq_idx,
  output [6:0]  io_iss_uops_2_pdst,
                io_iss_uops_2_prs1,
                io_iss_uops_2_prs2,
  output        io_iss_uops_2_bypassable,
  output [4:0]  io_iss_uops_2_mem_cmd,
  output        io_iss_uops_2_is_amo,
                io_iss_uops_2_uses_stq,
                io_iss_uops_2_ldst_val,
  output [1:0]  io_iss_uops_2_dst_rtype,
                io_iss_uops_2_lrs1_rtype,
                io_iss_uops_2_lrs2_rtype
);

  wire        issue_slots_31_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_30_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_29_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_28_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_27_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_26_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_25_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_24_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_23_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_22_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_21_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_20_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_19_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_18_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_17_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_16_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_15_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_14_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_13_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_12_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_11_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_10_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_9_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_8_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_7_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_6_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_5_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_4_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_3_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_2_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_1_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire        issue_slots_0_grant;	// issue-unit-age-ordered.scala:118:76, :119:30
  wire [2:0]  next_30;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_29;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_28;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_27;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_26;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_25;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_24;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_23;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_22;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_21;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_20;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_19;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_18;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_17;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_16;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_15;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_14;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_13;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_12;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_11;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_10;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_9;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_8;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_7;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_6;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_5;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_3;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [2:0]  next_2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire [1:0]  _next_1_1to0;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  wire        _slots_31_io_valid;	// issue-unit.scala:153:73
  wire        _slots_31_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_31_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_31_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_31_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_31_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_31_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_31_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_31_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_31_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_31_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_31_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_31_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_31_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_31_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_31_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_31_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_31_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_31_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_31_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_31_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_31_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_31_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_31_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_31_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_31_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_31_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_31_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_30_io_valid;	// issue-unit.scala:153:73
  wire        _slots_30_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_30_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_30_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_30_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_30_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_30_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_30_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_30_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_30_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_30_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_30_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_30_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_30_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_30_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_30_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_30_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_30_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_30_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_30_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_30_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_30_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_30_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_30_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_30_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_30_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_30_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_30_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_29_io_valid;	// issue-unit.scala:153:73
  wire        _slots_29_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_29_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_29_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_29_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_29_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_29_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_29_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_29_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_29_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_29_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_29_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_29_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_29_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_29_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_29_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_29_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_29_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_29_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_29_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_29_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_29_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_29_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_29_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_29_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_29_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_29_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_29_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_28_io_valid;	// issue-unit.scala:153:73
  wire        _slots_28_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_28_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_28_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_28_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_28_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_28_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_28_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_28_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_28_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_28_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_28_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_28_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_28_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_28_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_28_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_28_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_28_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_28_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_28_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_28_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_28_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_28_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_28_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_28_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_28_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_28_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_28_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_27_io_valid;	// issue-unit.scala:153:73
  wire        _slots_27_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_27_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_27_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_27_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_27_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_27_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_27_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_27_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_27_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_27_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_27_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_27_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_27_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_27_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_27_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_27_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_27_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_27_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_27_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_27_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_27_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_27_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_27_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_27_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_27_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_27_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_27_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_26_io_valid;	// issue-unit.scala:153:73
  wire        _slots_26_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_26_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_26_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_26_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_26_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_26_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_26_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_26_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_26_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_26_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_26_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_26_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_26_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_26_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_26_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_26_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_26_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_26_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_26_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_26_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_26_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_26_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_26_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_26_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_26_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_26_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_26_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_25_io_valid;	// issue-unit.scala:153:73
  wire        _slots_25_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_25_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_25_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_25_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_25_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_25_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_25_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_25_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_25_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_25_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_25_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_25_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_25_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_25_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_25_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_25_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_25_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_25_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_25_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_25_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_25_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_25_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_25_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_25_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_25_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_25_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_25_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_24_io_valid;	// issue-unit.scala:153:73
  wire        _slots_24_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_24_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_24_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_24_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_24_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_24_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_24_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_24_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_24_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_24_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_24_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_24_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_24_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_24_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_24_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_24_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_24_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_24_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_24_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_24_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_24_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_24_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_24_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_24_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_24_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_24_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_24_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_23_io_valid;	// issue-unit.scala:153:73
  wire        _slots_23_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_23_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_23_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_23_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_23_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_23_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_23_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_23_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_23_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_23_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_23_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_23_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_23_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_23_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_23_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_23_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_23_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_23_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_23_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_23_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_23_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_23_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_23_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_23_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_23_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_23_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_23_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_22_io_valid;	// issue-unit.scala:153:73
  wire        _slots_22_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_22_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_22_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_22_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_22_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_22_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_22_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_22_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_22_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_22_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_22_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_22_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_22_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_22_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_22_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_22_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_22_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_22_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_22_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_22_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_22_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_22_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_22_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_22_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_22_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_22_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_22_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_21_io_valid;	// issue-unit.scala:153:73
  wire        _slots_21_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_21_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_21_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_21_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_21_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_21_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_21_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_21_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_21_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_21_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_21_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_21_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_21_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_21_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_21_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_21_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_21_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_21_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_21_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_21_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_21_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_21_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_21_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_21_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_21_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_21_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_21_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_20_io_valid;	// issue-unit.scala:153:73
  wire        _slots_20_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_20_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_20_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_20_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_20_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_20_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_20_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_20_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_20_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_20_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_20_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_20_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_20_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_20_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_20_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_20_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_20_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_20_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_20_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_20_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_20_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_20_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_20_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_20_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_20_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_20_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_20_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_19_io_valid;	// issue-unit.scala:153:73
  wire        _slots_19_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_19_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_19_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_19_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_19_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_19_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_19_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_19_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_19_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_19_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_19_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_19_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_19_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_19_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_19_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_19_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_19_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_19_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_19_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_19_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_19_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_19_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_19_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_19_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_19_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_19_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_19_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_18_io_valid;	// issue-unit.scala:153:73
  wire        _slots_18_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_18_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_18_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_18_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_18_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_18_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_18_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_18_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_18_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_18_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_18_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_18_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_18_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_18_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_18_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_18_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_18_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_18_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_18_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_18_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_18_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_18_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_18_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_18_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_18_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_18_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_18_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_17_io_valid;	// issue-unit.scala:153:73
  wire        _slots_17_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_17_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_17_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_17_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_17_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_17_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_17_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_17_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_17_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_17_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_17_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_17_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_17_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_17_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_17_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_17_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_17_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_17_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_17_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_17_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_17_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_17_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_17_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_17_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_17_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_17_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_17_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_16_io_valid;	// issue-unit.scala:153:73
  wire        _slots_16_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_16_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_16_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_16_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_16_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_16_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_16_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_16_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_16_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_16_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_16_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_16_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_16_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_16_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_16_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_16_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_16_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_16_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_16_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_16_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_16_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_16_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_16_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_16_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_16_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_16_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_16_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_15_io_valid;	// issue-unit.scala:153:73
  wire        _slots_15_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_15_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_15_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_15_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_15_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_15_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_15_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_15_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_15_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_15_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_15_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_15_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_15_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_15_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_15_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_15_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_15_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_15_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_15_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_15_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_15_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_15_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_15_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_15_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_15_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_15_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_15_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_14_io_valid;	// issue-unit.scala:153:73
  wire        _slots_14_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_14_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_14_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_14_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_14_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_14_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_14_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_14_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_14_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_14_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_14_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_14_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_14_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_14_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_14_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_14_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_14_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_14_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_14_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_14_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_14_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_14_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_14_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_14_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_14_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_14_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_14_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_13_io_valid;	// issue-unit.scala:153:73
  wire        _slots_13_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_13_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_13_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_13_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_13_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_13_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_13_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_13_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_13_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_13_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_13_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_13_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_13_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_13_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_13_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_13_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_13_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_13_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_13_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_13_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_13_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_13_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_13_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_13_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_13_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_13_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_13_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_12_io_valid;	// issue-unit.scala:153:73
  wire        _slots_12_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_12_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_12_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_12_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_12_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_12_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_12_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_12_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_12_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_12_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_12_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_12_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_12_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_12_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_12_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_12_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_12_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_12_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_12_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_12_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_12_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_12_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_12_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_12_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_12_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_12_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_12_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_11_io_valid;	// issue-unit.scala:153:73
  wire        _slots_11_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_11_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_11_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_11_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_11_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_11_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_11_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_11_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_11_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_11_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_11_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_11_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_11_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_11_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_11_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_11_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_11_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_11_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_11_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_11_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_11_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_11_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_11_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_11_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_11_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_11_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_11_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_10_io_valid;	// issue-unit.scala:153:73
  wire        _slots_10_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_10_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_10_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_10_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_10_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_10_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_10_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_10_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_10_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_10_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_10_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_10_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_10_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_10_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_10_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_10_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_10_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_10_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_10_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_10_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_10_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_10_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_10_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_10_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_10_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_10_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_10_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_9_io_valid;	// issue-unit.scala:153:73
  wire        _slots_9_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_9_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_9_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_9_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_9_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_9_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_9_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_9_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_9_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_9_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_9_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_9_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_9_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_9_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_9_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_9_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_9_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_9_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_9_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_9_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_9_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_9_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_9_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_9_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_9_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_9_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_9_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_8_io_valid;	// issue-unit.scala:153:73
  wire        _slots_8_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_8_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_8_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_8_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_8_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_8_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_8_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_8_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_8_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_8_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_8_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_8_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_8_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_8_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_8_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_8_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_8_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_8_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_8_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_8_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_8_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_8_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_8_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_8_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_8_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_8_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_8_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_7_io_valid;	// issue-unit.scala:153:73
  wire        _slots_7_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_7_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_7_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_7_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_7_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_7_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_7_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_7_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_7_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_7_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_7_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_7_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_7_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_7_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_7_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_7_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_7_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_7_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_7_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_7_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_7_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_7_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_7_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_7_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_7_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_7_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_7_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_6_io_valid;	// issue-unit.scala:153:73
  wire        _slots_6_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_6_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_6_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_6_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_6_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_6_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_6_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_6_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_6_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_6_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_6_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_6_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_6_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_6_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_6_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_6_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_6_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_6_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_6_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_6_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_6_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_6_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_6_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_6_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_6_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_6_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_6_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_5_io_valid;	// issue-unit.scala:153:73
  wire        _slots_5_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_5_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_5_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_5_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_5_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_5_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_5_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_5_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_5_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_5_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_5_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_5_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_5_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_5_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_5_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_5_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_5_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_5_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_5_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_5_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_5_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_5_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_5_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_5_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_5_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_5_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_5_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_4_io_valid;	// issue-unit.scala:153:73
  wire        _slots_4_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_4_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_4_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_4_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_4_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_4_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_4_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_4_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_4_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_4_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_4_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_4_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_4_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_4_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_4_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_4_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_4_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_4_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_4_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_4_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_4_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_4_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_4_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_4_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_4_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_4_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_4_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_3_io_valid;	// issue-unit.scala:153:73
  wire        _slots_3_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_3_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_3_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_3_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_3_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_3_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_3_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_3_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_3_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_3_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_3_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_3_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_3_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_3_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_3_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_3_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_3_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_3_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_3_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_3_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_3_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_3_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_3_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_3_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_3_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_3_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_3_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_2_io_valid;	// issue-unit.scala:153:73
  wire        _slots_2_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_2_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_2_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_2_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_2_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_2_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_2_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_2_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_2_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_2_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_2_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_2_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_2_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_2_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_2_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_2_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_2_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_2_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_2_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_2_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_2_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_2_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_2_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_2_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_2_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_2_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_2_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_1_io_valid;	// issue-unit.scala:153:73
  wire        _slots_1_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_1_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_out_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_1_io_out_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_1_io_out_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_1_io_out_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_1_io_out_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_1_io_out_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_1_io_out_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_1_io_out_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_out_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_out_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_1_io_out_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_1_io_out_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_out_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_out_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_out_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_out_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_out_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_out_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_out_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_out_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_out_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_1_io_out_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_out_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_out_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_out_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_out_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_out_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_out_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_out_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_1_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_1_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_1_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_1_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_1_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_1_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_1_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_1_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_1_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_1_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_1_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_1_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_1_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_1_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_1_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _slots_0_io_valid;	// issue-unit.scala:153:73
  wire        _slots_0_io_will_be_valid;	// issue-unit.scala:153:73
  wire        _slots_0_io_request;	// issue-unit.scala:153:73
  wire [6:0]  _slots_0_io_uop_uopc;	// issue-unit.scala:153:73
  wire [31:0] _slots_0_io_uop_inst;	// issue-unit.scala:153:73
  wire [31:0] _slots_0_io_uop_debug_inst;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_rvc;	// issue-unit.scala:153:73
  wire [39:0] _slots_0_io_uop_debug_pc;	// issue-unit.scala:153:73
  wire [2:0]  _slots_0_io_uop_iq_type;	// issue-unit.scala:153:73
  wire [9:0]  _slots_0_io_uop_fu_code;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_iw_state;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_iw_p1_poisoned;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_iw_p2_poisoned;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_br;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_jalr;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_jal;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_sfb;	// issue-unit.scala:153:73
  wire [15:0] _slots_0_io_uop_br_mask;	// issue-unit.scala:153:73
  wire [3:0]  _slots_0_io_uop_br_tag;	// issue-unit.scala:153:73
  wire [4:0]  _slots_0_io_uop_ftq_idx;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_edge_inst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_0_io_uop_pc_lob;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_taken;	// issue-unit.scala:153:73
  wire [19:0] _slots_0_io_uop_imm_packed;	// issue-unit.scala:153:73
  wire [11:0] _slots_0_io_uop_csr_addr;	// issue-unit.scala:153:73
  wire [6:0]  _slots_0_io_uop_rob_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_0_io_uop_ldq_idx;	// issue-unit.scala:153:73
  wire [4:0]  _slots_0_io_uop_stq_idx;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_rxq_idx;	// issue-unit.scala:153:73
  wire [6:0]  _slots_0_io_uop_pdst;	// issue-unit.scala:153:73
  wire [6:0]  _slots_0_io_uop_prs1;	// issue-unit.scala:153:73
  wire [6:0]  _slots_0_io_uop_prs2;	// issue-unit.scala:153:73
  wire [6:0]  _slots_0_io_uop_prs3;	// issue-unit.scala:153:73
  wire [4:0]  _slots_0_io_uop_ppred;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_prs1_busy;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_prs2_busy;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_prs3_busy;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_ppred_busy;	// issue-unit.scala:153:73
  wire [6:0]  _slots_0_io_uop_stale_pdst;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_exception;	// issue-unit.scala:153:73
  wire [63:0] _slots_0_io_uop_exc_cause;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_bypassable;	// issue-unit.scala:153:73
  wire [4:0]  _slots_0_io_uop_mem_cmd;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_mem_size;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_mem_signed;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_fence;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_fencei;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_amo;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_uses_ldq;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_uses_stq;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_sys_pc2epc;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_is_unique;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_flush_on_commit;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_ldst_is_rs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_0_io_uop_ldst;	// issue-unit.scala:153:73
  wire [5:0]  _slots_0_io_uop_lrs1;	// issue-unit.scala:153:73
  wire [5:0]  _slots_0_io_uop_lrs2;	// issue-unit.scala:153:73
  wire [5:0]  _slots_0_io_uop_lrs3;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_ldst_val;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_dst_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_lrs1_rtype;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_lrs2_rtype;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_frs3_en;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_fp_val;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_fp_single;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_xcpt_pf_if;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_xcpt_ae_if;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_xcpt_ma_if;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_bp_debug_if;	// issue-unit.scala:153:73
  wire        _slots_0_io_uop_bp_xcpt_if;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_debug_fsrc;	// issue-unit.scala:153:73
  wire [1:0]  _slots_0_io_uop_debug_tsrc;	// issue-unit.scala:153:73
  wire        _GEN = io_dis_uops_0_bits_uopc == 7'h2;	// issue-unit.scala:127:39
  wire        _GEN_0 =
    _GEN & ~(|io_dis_uops_0_bits_lrs2_rtype) | io_dis_uops_0_bits_uopc == 7'h43;	// issue-unit.scala:127:{39,50,84,96}, :128:39
  wire [1:0]  uops_32_iw_state = _GEN_0 ? 2'h2 : 2'h1;	// issue-unit.scala:123:26, :127:96, :128:54, :129:30
  wire        _GEN_1 = _GEN_0 | ~(_GEN & (|io_dis_uops_0_bits_lrs2_rtype));	// issue-unit.scala:120:17, :127:{39,84,96}, :128:54, :131:{56,102}
  wire [1:0]  uops_32_lrs2_rtype = _GEN_1 ? io_dis_uops_0_bits_lrs2_rtype : 2'h2;	// issue-unit.scala:120:17, :128:54, :129:30, :131:102
  wire        uops_32_prs2_busy = _GEN_1 & io_dis_uops_0_bits_prs2_busy;	// issue-unit.scala:120:17, :128:54, :131:102
  wire        _GEN_2 = io_dis_uops_1_bits_uopc == 7'h2;	// issue-unit.scala:127:39
  wire        _GEN_3 =
    _GEN_2 & ~(|io_dis_uops_1_bits_lrs2_rtype) | io_dis_uops_1_bits_uopc == 7'h43;	// issue-unit.scala:127:{39,50,84,96}, :128:39
  wire        _GEN_4 = _GEN_3 | ~(_GEN_2 & (|io_dis_uops_1_bits_lrs2_rtype));	// issue-unit.scala:120:17, :127:{39,84,96}, :128:54, :131:{56,102}
  wire [1:0]  uops_33_lrs2_rtype = _GEN_4 ? io_dis_uops_1_bits_lrs2_rtype : 2'h2;	// issue-unit.scala:120:17, :128:54, :129:30, :131:102
  wire        uops_33_prs2_busy = _GEN_4 & io_dis_uops_1_bits_prs2_busy;	// issue-unit.scala:120:17, :128:54, :131:102
  wire        _GEN_5 = io_dis_uops_2_bits_uopc == 7'h2;	// issue-unit.scala:127:39
  wire        _GEN_6 =
    _GEN_5 & ~(|io_dis_uops_2_bits_lrs2_rtype) | io_dis_uops_2_bits_uopc == 7'h43;	// issue-unit.scala:127:{39,50,84,96}, :128:39
  wire        _GEN_7 = _GEN_6 | ~(_GEN_5 & (|io_dis_uops_2_bits_lrs2_rtype));	// issue-unit.scala:120:17, :127:{39,84,96}, :128:54, :131:{56,102}
  `ifndef SYNTHESIS	// issue-unit.scala:172:10
    always @(posedge clock) begin	// issue-unit.scala:172:10
      if (~({1'h0,
             {1'h0,
              {1'h0,
               {1'h0, {1'h0, issue_slots_0_grant} + {1'h0, issue_slots_1_grant}}
                 + {1'h0, {1'h0, issue_slots_2_grant} + {1'h0, issue_slots_3_grant}}}
                + {1'h0,
                   {1'h0, {1'h0, issue_slots_4_grant} + {1'h0, issue_slots_5_grant}}
                     + {1'h0, {1'h0, issue_slots_6_grant} + {1'h0, issue_slots_7_grant}}}}
               + {1'h0,
                  {1'h0,
                   {1'h0, {1'h0, issue_slots_8_grant} + {1'h0, issue_slots_9_grant}}
                     + {1'h0,
                        {1'h0, issue_slots_10_grant} + {1'h0, issue_slots_11_grant}}}
                    + {1'h0,
                       {1'h0, {1'h0, issue_slots_12_grant} + {1'h0, issue_slots_13_grant}}
                         + {1'h0,
                            {1'h0, issue_slots_14_grant}
                              + {1'h0, issue_slots_15_grant}}}}}
            + {1'h0,
               {1'h0,
                {1'h0,
                 {1'h0, {1'h0, issue_slots_16_grant} + {1'h0, issue_slots_17_grant}}
                   + {1'h0, {1'h0, issue_slots_18_grant} + {1'h0, issue_slots_19_grant}}}
                  + {1'h0,
                     {1'h0, {1'h0, issue_slots_20_grant} + {1'h0, issue_slots_21_grant}}
                       + {1'h0,
                          {1'h0, issue_slots_22_grant} + {1'h0, issue_slots_23_grant}}}}
                 + {1'h0,
                    {1'h0,
                     {1'h0, {1'h0, issue_slots_24_grant} + {1'h0, issue_slots_25_grant}}
                       + {1'h0,
                          {1'h0, issue_slots_26_grant} + {1'h0, issue_slots_27_grant}}}
                      + {1'h0,
                         {1'h0,
                          {1'h0, issue_slots_28_grant} + {1'h0, issue_slots_29_grant}}
                           + {1'h0,
                              {1'h0, issue_slots_30_grant}
                                + {1'h0, issue_slots_31_grant}}}}} < 6'h4 | reset)) begin	// Bitwise.scala:47:55, issue-unit-age-ordered.scala:118:76, :119:30, issue-unit.scala:172:{10,51}
        if (`ASSERT_VERBOSE_COND_)	// issue-unit.scala:172:10
          $error("Assertion failed: [issue] window giving out too many grants.\n    at issue-unit.scala:172 assert (PopCount(issue_slots.map(s => s.grant)) <= issueWidth.U, \"[issue] window giving out too many grants.\")\n");	// issue-unit.scala:172:10
        if (`STOP_COND_)	// issue-unit.scala:172:10
          $fatal;	// issue-unit.scala:172:10
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire [2:0]  next_1 =
    _slots_0_io_valid & ~_slots_1_io_valid
      ? 3'h1
      : _slots_1_io_valid ? {2'h0, ~_slots_0_io_valid} : {1'h0, ~_slots_0_io_valid, 1'h0};	// issue-unit-age-ordered.scala:39:38, :44:11, :45:{29,37}, :46:13, :47:44, :48:13, issue-unit.scala:127:84, :153:73
  assign _next_1_1to0 = next_1[1:0];	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44
  assign next_2 =
    _next_1_1to0 == 2'h0 & ~_slots_2_io_valid
      ? 3'h1
      : next_1[2] | _slots_2_io_valid ? next_1 : {_next_1_1to0, 1'h0};	// issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:127:84, :153:73
  assign next_3 =
    next_2 == 3'h0 & ~_slots_3_io_valid
      ? 3'h1
      : next_2[2] | _slots_3_io_valid ? next_2 : {next_2[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_4 =
    next_3 == 3'h0 & ~_slots_4_io_valid
      ? 3'h1
      : next_3[2] | _slots_4_io_valid ? next_3 : {next_3[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_5 =
    next_4 == 3'h0 & ~_slots_5_io_valid
      ? 3'h1
      : next_4[2] | _slots_5_io_valid ? next_4 : {next_4[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_6 =
    next_5 == 3'h0 & ~_slots_6_io_valid
      ? 3'h1
      : next_5[2] | _slots_6_io_valid ? next_5 : {next_5[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_7 =
    next_6 == 3'h0 & ~_slots_7_io_valid
      ? 3'h1
      : next_6[2] | _slots_7_io_valid ? next_6 : {next_6[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_8 =
    next_7 == 3'h0 & ~_slots_8_io_valid
      ? 3'h1
      : next_7[2] | _slots_8_io_valid ? next_7 : {next_7[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_9 =
    next_8 == 3'h0 & ~_slots_9_io_valid
      ? 3'h1
      : next_8[2] | _slots_9_io_valid ? next_8 : {next_8[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_10 =
    next_9 == 3'h0 & ~_slots_10_io_valid
      ? 3'h1
      : next_9[2] | _slots_10_io_valid ? next_9 : {next_9[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_11 =
    next_10 == 3'h0 & ~_slots_11_io_valid
      ? 3'h1
      : next_10[2] | _slots_11_io_valid ? next_10 : {next_10[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_12 =
    next_11 == 3'h0 & ~_slots_12_io_valid
      ? 3'h1
      : next_11[2] | _slots_12_io_valid ? next_11 : {next_11[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_13 =
    next_12 == 3'h0 & ~_slots_13_io_valid
      ? 3'h1
      : next_12[2] | _slots_13_io_valid ? next_12 : {next_12[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_14 =
    next_13 == 3'h0 & ~_slots_14_io_valid
      ? 3'h1
      : next_13[2] | _slots_14_io_valid ? next_13 : {next_13[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_15 =
    next_14 == 3'h0 & ~_slots_15_io_valid
      ? 3'h1
      : next_14[2] | _slots_15_io_valid ? next_14 : {next_14[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_16 =
    next_15 == 3'h0 & ~_slots_16_io_valid
      ? 3'h1
      : next_15[2] | _slots_16_io_valid ? next_15 : {next_15[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_17 =
    next_16 == 3'h0 & ~_slots_17_io_valid
      ? 3'h1
      : next_16[2] | _slots_17_io_valid ? next_16 : {next_16[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_18 =
    next_17 == 3'h0 & ~_slots_18_io_valid
      ? 3'h1
      : next_17[2] | _slots_18_io_valid ? next_17 : {next_17[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_19 =
    next_18 == 3'h0 & ~_slots_19_io_valid
      ? 3'h1
      : next_18[2] | _slots_19_io_valid ? next_18 : {next_18[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_20 =
    next_19 == 3'h0 & ~_slots_20_io_valid
      ? 3'h1
      : next_19[2] | _slots_20_io_valid ? next_19 : {next_19[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_21 =
    next_20 == 3'h0 & ~_slots_21_io_valid
      ? 3'h1
      : next_20[2] | _slots_21_io_valid ? next_20 : {next_20[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_22 =
    next_21 == 3'h0 & ~_slots_22_io_valid
      ? 3'h1
      : next_21[2] | _slots_22_io_valid ? next_21 : {next_21[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_23 =
    next_22 == 3'h0 & ~_slots_23_io_valid
      ? 3'h1
      : next_22[2] | _slots_23_io_valid ? next_22 : {next_22[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_24 =
    next_23 == 3'h0 & ~_slots_24_io_valid
      ? 3'h1
      : next_23[2] | _slots_24_io_valid ? next_23 : {next_23[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_25 =
    next_24 == 3'h0 & ~_slots_25_io_valid
      ? 3'h1
      : next_24[2] | _slots_25_io_valid ? next_24 : {next_24[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_26 =
    next_25 == 3'h0 & ~_slots_26_io_valid
      ? 3'h1
      : next_25[2] | _slots_26_io_valid ? next_25 : {next_25[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_27 =
    next_26 == 3'h0 & ~_slots_27_io_valid
      ? 3'h1
      : next_26[2] | _slots_27_io_valid ? next_26 : {next_26[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_28 =
    next_27 == 3'h0 & ~_slots_28_io_valid
      ? 3'h1
      : next_27[2] | _slots_28_io_valid ? next_27 : {next_27[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_29 =
    next_28 == 3'h0 & ~_slots_29_io_valid
      ? 3'h1
      : next_28[2] | _slots_29_io_valid ? next_28 : {next_28[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  assign next_30 =
    next_29 == 3'h0 & ~_slots_30_io_valid
      ? 3'h1
      : next_29[2] | _slots_30_io_valid ? next_29 : {next_29[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  wire [2:0]  next_31 =
    next_30 == 3'h0 & ~_slots_31_io_valid
      ? 3'h1
      : next_30[2] | _slots_31_io_valid ? next_30 : {next_30[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:38, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, issue-unit.scala:153:73
  wire [2:0]  next_32 =
    next_31 == 3'h0 & ~io_dis_uops_0_valid
      ? 3'h1
      : next_31[2] | io_dis_uops_0_valid ? next_31 : {next_31[1:0], 1'h0};	// consts.scala:270:20, issue-unit-age-ordered.scala:39:82, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13
  wire        will_be_valid_32 =
    io_dis_uops_0_valid & ~io_dis_uops_0_bits_exception & ~io_dis_uops_0_bits_is_fence
    & ~io_dis_uops_0_bits_is_fencei;	// issue-unit-age-ordered.scala:62:57, :63:{57,79}, :64:57
  wire        will_be_valid_33 =
    io_dis_uops_1_valid & ~io_dis_uops_1_bits_exception & ~io_dis_uops_1_bits_is_fence
    & ~io_dis_uops_1_bits_is_fencei;	// issue-unit-age-ordered.scala:62:57, :63:{57,79}, :64:57
  wire        _GEN_8 = _next_1_1to0 == 2'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28, issue-unit.scala:129:30
  wire        _GEN_9 = next_2 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_0_in_uop_valid =
    _GEN_9
      ? _slots_3_io_will_be_valid
      : _GEN_8
          ? _slots_2_io_will_be_valid
          : ~_slots_0_io_valid & _slots_1_io_will_be_valid;	// issue-unit-age-ordered.scala:39:38, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_10 = next_2 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_11 = next_3 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_1_in_uop_valid =
    _GEN_11
      ? _slots_4_io_will_be_valid
      : _GEN_10
          ? _slots_3_io_will_be_valid
          : _next_1_1to0 == 2'h1 & _slots_2_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:123:26, :153:73
  wire        _GEN_12 = next_3 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_13 = next_4 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_2_in_uop_valid =
    _GEN_13
      ? _slots_5_io_will_be_valid
      : _GEN_12 ? _slots_4_io_will_be_valid : next_2 == 3'h1 & _slots_3_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_14 = next_4 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_15 = next_5 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_3_in_uop_valid =
    _GEN_15
      ? _slots_6_io_will_be_valid
      : _GEN_14 ? _slots_5_io_will_be_valid : next_3 == 3'h1 & _slots_4_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_16 = next_5 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_17 = next_6 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_4_in_uop_valid =
    _GEN_17
      ? _slots_7_io_will_be_valid
      : _GEN_16 ? _slots_6_io_will_be_valid : next_4 == 3'h1 & _slots_5_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_18 = next_6 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_19 = next_7 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_5_in_uop_valid =
    _GEN_19
      ? _slots_8_io_will_be_valid
      : _GEN_18 ? _slots_7_io_will_be_valid : next_5 == 3'h1 & _slots_6_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_20 = next_7 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_21 = next_8 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_6_in_uop_valid =
    _GEN_21
      ? _slots_9_io_will_be_valid
      : _GEN_20 ? _slots_8_io_will_be_valid : next_6 == 3'h1 & _slots_7_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_22 = next_8 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_23 = next_9 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_7_in_uop_valid =
    _GEN_23
      ? _slots_10_io_will_be_valid
      : _GEN_22 ? _slots_9_io_will_be_valid : next_7 == 3'h1 & _slots_8_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_24 = next_9 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_25 = next_10 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_8_in_uop_valid =
    _GEN_25
      ? _slots_11_io_will_be_valid
      : _GEN_24 ? _slots_10_io_will_be_valid : next_8 == 3'h1 & _slots_9_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_26 = next_10 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_27 = next_11 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_9_in_uop_valid =
    _GEN_27
      ? _slots_12_io_will_be_valid
      : _GEN_26
          ? _slots_11_io_will_be_valid
          : next_9 == 3'h1 & _slots_10_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_28 = next_11 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_29 = next_12 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_10_in_uop_valid =
    _GEN_29
      ? _slots_13_io_will_be_valid
      : _GEN_28
          ? _slots_12_io_will_be_valid
          : next_10 == 3'h1 & _slots_11_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_30 = next_12 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_31 = next_13 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_11_in_uop_valid =
    _GEN_31
      ? _slots_14_io_will_be_valid
      : _GEN_30
          ? _slots_13_io_will_be_valid
          : next_11 == 3'h1 & _slots_12_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_32 = next_13 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_33 = next_14 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_12_in_uop_valid =
    _GEN_33
      ? _slots_15_io_will_be_valid
      : _GEN_32
          ? _slots_14_io_will_be_valid
          : next_12 == 3'h1 & _slots_13_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_34 = next_14 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_35 = next_15 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_13_in_uop_valid =
    _GEN_35
      ? _slots_16_io_will_be_valid
      : _GEN_34
          ? _slots_15_io_will_be_valid
          : next_13 == 3'h1 & _slots_14_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_36 = next_15 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_37 = next_16 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_14_in_uop_valid =
    _GEN_37
      ? _slots_17_io_will_be_valid
      : _GEN_36
          ? _slots_16_io_will_be_valid
          : next_14 == 3'h1 & _slots_15_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_38 = next_16 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_39 = next_17 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_15_in_uop_valid =
    _GEN_39
      ? _slots_18_io_will_be_valid
      : _GEN_38
          ? _slots_17_io_will_be_valid
          : next_15 == 3'h1 & _slots_16_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_40 = next_17 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_41 = next_18 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_16_in_uop_valid =
    _GEN_41
      ? _slots_19_io_will_be_valid
      : _GEN_40
          ? _slots_18_io_will_be_valid
          : next_16 == 3'h1 & _slots_17_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_42 = next_18 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_43 = next_19 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_17_in_uop_valid =
    _GEN_43
      ? _slots_20_io_will_be_valid
      : _GEN_42
          ? _slots_19_io_will_be_valid
          : next_17 == 3'h1 & _slots_18_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_44 = next_19 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_45 = next_20 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_18_in_uop_valid =
    _GEN_45
      ? _slots_21_io_will_be_valid
      : _GEN_44
          ? _slots_20_io_will_be_valid
          : next_18 == 3'h1 & _slots_19_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_46 = next_20 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_47 = next_21 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_19_in_uop_valid =
    _GEN_47
      ? _slots_22_io_will_be_valid
      : _GEN_46
          ? _slots_21_io_will_be_valid
          : next_19 == 3'h1 & _slots_20_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_48 = next_21 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_49 = next_22 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_20_in_uop_valid =
    _GEN_49
      ? _slots_23_io_will_be_valid
      : _GEN_48
          ? _slots_22_io_will_be_valid
          : next_20 == 3'h1 & _slots_21_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_50 = next_22 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_51 = next_23 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_21_in_uop_valid =
    _GEN_51
      ? _slots_24_io_will_be_valid
      : _GEN_50
          ? _slots_23_io_will_be_valid
          : next_21 == 3'h1 & _slots_22_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_52 = next_23 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_53 = next_24 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_22_in_uop_valid =
    _GEN_53
      ? _slots_25_io_will_be_valid
      : _GEN_52
          ? _slots_24_io_will_be_valid
          : next_22 == 3'h1 & _slots_23_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_54 = next_24 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_55 = next_25 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_23_in_uop_valid =
    _GEN_55
      ? _slots_26_io_will_be_valid
      : _GEN_54
          ? _slots_25_io_will_be_valid
          : next_23 == 3'h1 & _slots_24_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_56 = next_25 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_57 = next_26 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_24_in_uop_valid =
    _GEN_57
      ? _slots_27_io_will_be_valid
      : _GEN_56
          ? _slots_26_io_will_be_valid
          : next_24 == 3'h1 & _slots_25_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_58 = next_26 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_59 = next_27 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_25_in_uop_valid =
    _GEN_59
      ? _slots_28_io_will_be_valid
      : _GEN_58
          ? _slots_27_io_will_be_valid
          : next_25 == 3'h1 & _slots_26_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_60 = next_27 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_61 = next_28 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_26_in_uop_valid =
    _GEN_61
      ? _slots_29_io_will_be_valid
      : _GEN_60
          ? _slots_28_io_will_be_valid
          : next_26 == 3'h1 & _slots_27_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_62 = next_28 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_63 = next_29 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_27_in_uop_valid =
    _GEN_63
      ? _slots_30_io_will_be_valid
      : _GEN_62
          ? _slots_29_io_will_be_valid
          : next_27 == 3'h1 & _slots_28_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_64 = next_29 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_65 = next_30 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_28_in_uop_valid =
    _GEN_65
      ? _slots_31_io_will_be_valid
      : _GEN_64
          ? _slots_30_io_will_be_valid
          : next_28 == 3'h1 & _slots_29_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_66 = next_30 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_67 = next_31 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_29_in_uop_valid =
    _GEN_67
      ? will_be_valid_32
      : _GEN_66
          ? _slots_31_io_will_be_valid
          : next_29 == 3'h1 & _slots_30_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :63:79, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_68 = next_31 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_69 = next_32 == 3'h4;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        issue_slots_30_in_uop_valid =
    _GEN_69
      ? will_be_valid_33
      : _GEN_68 ? will_be_valid_32 : next_30 == 3'h1 & _slots_31_io_will_be_valid;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :63:79, :68:33, :71:{28,48}, :72:37, issue-unit.scala:153:73
  wire        _GEN_70 = _GEN_69 | _GEN_68;	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
  wire        _GEN_71 = next_32 == 3'h2;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :71:28
  wire        _GEN_72 =
    (next_32 == 3'h0 & ~io_dis_uops_1_valid
       ? 3'h1
       : next_32[2] | io_dis_uops_1_valid ? next_32 : {next_32[1:0], 1'h0}) == 3'h4;	// consts.scala:270:20, issue-unit-age-ordered.scala:39:82, :44:11, :45:{21,29,37}, :46:13, :47:{28,44}, :48:13, :71:28
  wire        issue_slots_31_in_uop_valid =
    _GEN_72
      ? io_dis_uops_2_valid & ~io_dis_uops_2_bits_exception & ~io_dis_uops_2_bits_is_fence
        & ~io_dis_uops_2_bits_is_fencei
      : _GEN_71 ? will_be_valid_33 : next_31 == 3'h1 & will_be_valid_32;	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :62:57, :63:{57,79}, :64:57, :68:33, :71:{28,48}, :72:37
  reg         io_dis_uops_0_ready_REG;	// issue-unit-age-ordered.scala:87:36
  reg         io_dis_uops_1_ready_REG;	// issue-unit-age-ordered.scala:87:36
  reg         io_dis_uops_2_ready_REG;	// issue-unit-age-ordered.scala:87:36
  wire        _GEN_73 =
    _slots_0_io_request & (|(_slots_0_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire [9:0]  _can_allocate_T_1 = _slots_0_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_74 = _slots_0_io_request & ~_GEN_73 & (|_can_allocate_T_1);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40}, issue-unit.scala:153:73
  wire        _GEN_75 =
    _slots_0_io_request & ~(_slots_0_io_request & (|_can_allocate_T_1) | _GEN_73)
    & (|(_slots_0_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40}, :125:{33,74}, issue-unit.scala:153:73
  assign issue_slots_0_grant = _GEN_75 | _GEN_74 | _GEN_73;	// issue-unit-age-ordered.scala:118:{40,76}, :119:30
  wire        _GEN_76 =
    _slots_1_io_request & (|(_slots_1_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_77 = _GEN_76 & ~_GEN_73;	// issue-unit-age-ordered.scala:118:{28,40,56}
  wire        _GEN_78 = _GEN_76 | _GEN_73;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_4 = _slots_1_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_79 = _slots_1_io_request & ~_GEN_77 & (|_can_allocate_T_4);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_80 = _GEN_79 & ~_GEN_74;	// issue-unit-age-ordered.scala:118:{40,56,59}
  wire        _GEN_81 = _GEN_79 | _GEN_74;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_82 =
    _slots_1_io_request
    & ~(_slots_1_io_request & (|_can_allocate_T_4) & ~_GEN_74 | _GEN_77)
    & (|(_slots_1_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_83 = _GEN_82 & ~_GEN_75;	// issue-unit-age-ordered.scala:118:{40,56,59}
  assign issue_slots_1_grant = _GEN_83 | _GEN_80 | _GEN_77;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_84 = _GEN_82 | _GEN_75;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_85 =
    _slots_2_io_request & (|(_slots_2_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_86 = _GEN_85 & ~_GEN_78;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_87 = _GEN_85 | _GEN_78;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_7 = _slots_2_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_88 = _slots_2_io_request & ~_GEN_86 & (|_can_allocate_T_7);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_89 = _GEN_88 & ~_GEN_81;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_90 = _GEN_88 | _GEN_81;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_91 =
    _slots_2_io_request
    & ~(_slots_2_io_request & (|_can_allocate_T_7) & ~_GEN_81 | _GEN_86)
    & (|(_slots_2_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_92 = _GEN_91 & ~_GEN_84;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_2_grant = _GEN_92 | _GEN_89 | _GEN_86;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_93 = _GEN_91 | _GEN_84;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_94 =
    _slots_3_io_request & (|(_slots_3_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_95 = _GEN_94 & ~_GEN_87;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_96 = _GEN_94 | _GEN_87;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_10 = _slots_3_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_97 = _slots_3_io_request & ~_GEN_95 & (|_can_allocate_T_10);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_98 = _GEN_97 & ~_GEN_90;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_99 = _GEN_97 | _GEN_90;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_100 =
    _slots_3_io_request
    & ~(_slots_3_io_request & (|_can_allocate_T_10) & ~_GEN_90 | _GEN_95)
    & (|(_slots_3_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_101 = _GEN_100 & ~_GEN_93;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_3_grant = _GEN_101 | _GEN_98 | _GEN_95;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_102 = _GEN_100 | _GEN_93;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_103 =
    _slots_4_io_request & (|(_slots_4_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_104 = _GEN_103 & ~_GEN_96;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_105 = _GEN_103 | _GEN_96;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_13 = _slots_4_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_106 = _slots_4_io_request & ~_GEN_104 & (|_can_allocate_T_13);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_107 = _GEN_106 & ~_GEN_99;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_108 = _GEN_106 | _GEN_99;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_109 =
    _slots_4_io_request
    & ~(_slots_4_io_request & (|_can_allocate_T_13) & ~_GEN_99 | _GEN_104)
    & (|(_slots_4_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_110 = _GEN_109 & ~_GEN_102;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_4_grant = _GEN_110 | _GEN_107 | _GEN_104;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_111 = _GEN_109 | _GEN_102;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_112 =
    _slots_5_io_request & (|(_slots_5_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_113 = _GEN_112 & ~_GEN_105;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_114 = _GEN_112 | _GEN_105;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_16 = _slots_5_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_115 = _slots_5_io_request & ~_GEN_113 & (|_can_allocate_T_16);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_116 = _GEN_115 & ~_GEN_108;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_117 = _GEN_115 | _GEN_108;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_118 =
    _slots_5_io_request
    & ~(_slots_5_io_request & (|_can_allocate_T_16) & ~_GEN_108 | _GEN_113)
    & (|(_slots_5_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_119 = _GEN_118 & ~_GEN_111;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_5_grant = _GEN_119 | _GEN_116 | _GEN_113;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_120 = _GEN_118 | _GEN_111;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_121 =
    _slots_6_io_request & (|(_slots_6_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_122 = _GEN_121 & ~_GEN_114;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_123 = _GEN_121 | _GEN_114;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_19 = _slots_6_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_124 = _slots_6_io_request & ~_GEN_122 & (|_can_allocate_T_19);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_125 = _GEN_124 & ~_GEN_117;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_126 = _GEN_124 | _GEN_117;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_127 =
    _slots_6_io_request
    & ~(_slots_6_io_request & (|_can_allocate_T_19) & ~_GEN_117 | _GEN_122)
    & (|(_slots_6_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_128 = _GEN_127 & ~_GEN_120;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_6_grant = _GEN_128 | _GEN_125 | _GEN_122;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_129 = _GEN_127 | _GEN_120;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_130 =
    _slots_7_io_request & (|(_slots_7_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_131 = _GEN_130 & ~_GEN_123;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_132 = _GEN_130 | _GEN_123;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_22 = _slots_7_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_133 = _slots_7_io_request & ~_GEN_131 & (|_can_allocate_T_22);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_134 = _GEN_133 & ~_GEN_126;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_135 = _GEN_133 | _GEN_126;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_136 =
    _slots_7_io_request
    & ~(_slots_7_io_request & (|_can_allocate_T_22) & ~_GEN_126 | _GEN_131)
    & (|(_slots_7_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_137 = _GEN_136 & ~_GEN_129;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_7_grant = _GEN_137 | _GEN_134 | _GEN_131;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_138 = _GEN_136 | _GEN_129;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_139 =
    _slots_8_io_request & (|(_slots_8_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_140 = _GEN_139 & ~_GEN_132;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_141 = _GEN_139 | _GEN_132;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_25 = _slots_8_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_142 = _slots_8_io_request & ~_GEN_140 & (|_can_allocate_T_25);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_143 = _GEN_142 & ~_GEN_135;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_144 = _GEN_142 | _GEN_135;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_145 =
    _slots_8_io_request
    & ~(_slots_8_io_request & (|_can_allocate_T_25) & ~_GEN_135 | _GEN_140)
    & (|(_slots_8_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_146 = _GEN_145 & ~_GEN_138;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_8_grant = _GEN_146 | _GEN_143 | _GEN_140;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_147 = _GEN_145 | _GEN_138;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_148 =
    _slots_9_io_request & (|(_slots_9_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_149 = _GEN_148 & ~_GEN_141;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_150 = _GEN_148 | _GEN_141;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_28 = _slots_9_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_151 = _slots_9_io_request & ~_GEN_149 & (|_can_allocate_T_28);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_152 = _GEN_151 & ~_GEN_144;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_153 = _GEN_151 | _GEN_144;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_154 =
    _slots_9_io_request
    & ~(_slots_9_io_request & (|_can_allocate_T_28) & ~_GEN_144 | _GEN_149)
    & (|(_slots_9_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_155 = _GEN_154 & ~_GEN_147;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_9_grant = _GEN_155 | _GEN_152 | _GEN_149;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_156 = _GEN_154 | _GEN_147;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_157 =
    _slots_10_io_request & (|(_slots_10_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_158 = _GEN_157 & ~_GEN_150;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_159 = _GEN_157 | _GEN_150;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_31 = _slots_10_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_160 = _slots_10_io_request & ~_GEN_158 & (|_can_allocate_T_31);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_161 = _GEN_160 & ~_GEN_153;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_162 = _GEN_160 | _GEN_153;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_163 =
    _slots_10_io_request
    & ~(_slots_10_io_request & (|_can_allocate_T_31) & ~_GEN_153 | _GEN_158)
    & (|(_slots_10_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_164 = _GEN_163 & ~_GEN_156;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_10_grant = _GEN_164 | _GEN_161 | _GEN_158;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_165 = _GEN_163 | _GEN_156;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_166 =
    _slots_11_io_request & (|(_slots_11_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_167 = _GEN_166 & ~_GEN_159;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_168 = _GEN_166 | _GEN_159;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_34 = _slots_11_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_169 = _slots_11_io_request & ~_GEN_167 & (|_can_allocate_T_34);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_170 = _GEN_169 & ~_GEN_162;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_171 = _GEN_169 | _GEN_162;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_172 =
    _slots_11_io_request
    & ~(_slots_11_io_request & (|_can_allocate_T_34) & ~_GEN_162 | _GEN_167)
    & (|(_slots_11_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_173 = _GEN_172 & ~_GEN_165;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_11_grant = _GEN_173 | _GEN_170 | _GEN_167;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_174 = _GEN_172 | _GEN_165;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_175 =
    _slots_12_io_request & (|(_slots_12_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_176 = _GEN_175 & ~_GEN_168;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_177 = _GEN_175 | _GEN_168;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_37 = _slots_12_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_178 = _slots_12_io_request & ~_GEN_176 & (|_can_allocate_T_37);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_179 = _GEN_178 & ~_GEN_171;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_180 = _GEN_178 | _GEN_171;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_181 =
    _slots_12_io_request
    & ~(_slots_12_io_request & (|_can_allocate_T_37) & ~_GEN_171 | _GEN_176)
    & (|(_slots_12_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_182 = _GEN_181 & ~_GEN_174;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_12_grant = _GEN_182 | _GEN_179 | _GEN_176;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_183 = _GEN_181 | _GEN_174;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_184 =
    _slots_13_io_request & (|(_slots_13_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_185 = _GEN_184 & ~_GEN_177;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_186 = _GEN_184 | _GEN_177;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_40 = _slots_13_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_187 = _slots_13_io_request & ~_GEN_185 & (|_can_allocate_T_40);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_188 = _GEN_187 & ~_GEN_180;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_189 = _GEN_187 | _GEN_180;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_190 =
    _slots_13_io_request
    & ~(_slots_13_io_request & (|_can_allocate_T_40) & ~_GEN_180 | _GEN_185)
    & (|(_slots_13_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_191 = _GEN_190 & ~_GEN_183;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_13_grant = _GEN_191 | _GEN_188 | _GEN_185;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_192 = _GEN_190 | _GEN_183;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_193 =
    _slots_14_io_request & (|(_slots_14_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_194 = _GEN_193 & ~_GEN_186;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_195 = _GEN_193 | _GEN_186;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_43 = _slots_14_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_196 = _slots_14_io_request & ~_GEN_194 & (|_can_allocate_T_43);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_197 = _GEN_196 & ~_GEN_189;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_198 = _GEN_196 | _GEN_189;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_199 =
    _slots_14_io_request
    & ~(_slots_14_io_request & (|_can_allocate_T_43) & ~_GEN_189 | _GEN_194)
    & (|(_slots_14_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_200 = _GEN_199 & ~_GEN_192;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_14_grant = _GEN_200 | _GEN_197 | _GEN_194;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_201 = _GEN_199 | _GEN_192;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_202 =
    _slots_15_io_request & (|(_slots_15_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_203 = _GEN_202 & ~_GEN_195;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_204 = _GEN_202 | _GEN_195;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_46 = _slots_15_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_205 = _slots_15_io_request & ~_GEN_203 & (|_can_allocate_T_46);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_206 = _GEN_205 & ~_GEN_198;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_207 = _GEN_205 | _GEN_198;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_208 =
    _slots_15_io_request
    & ~(_slots_15_io_request & (|_can_allocate_T_46) & ~_GEN_198 | _GEN_203)
    & (|(_slots_15_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_209 = _GEN_208 & ~_GEN_201;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_15_grant = _GEN_209 | _GEN_206 | _GEN_203;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_210 = _GEN_208 | _GEN_201;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_211 =
    _slots_16_io_request & (|(_slots_16_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_212 = _GEN_211 & ~_GEN_204;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_213 = _GEN_211 | _GEN_204;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_49 = _slots_16_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_214 = _slots_16_io_request & ~_GEN_212 & (|_can_allocate_T_49);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_215 = _GEN_214 & ~_GEN_207;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_216 = _GEN_214 | _GEN_207;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_217 =
    _slots_16_io_request
    & ~(_slots_16_io_request & (|_can_allocate_T_49) & ~_GEN_207 | _GEN_212)
    & (|(_slots_16_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_218 = _GEN_217 & ~_GEN_210;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_16_grant = _GEN_218 | _GEN_215 | _GEN_212;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_219 = _GEN_217 | _GEN_210;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_220 =
    _slots_17_io_request & (|(_slots_17_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_221 = _GEN_220 & ~_GEN_213;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_222 = _GEN_220 | _GEN_213;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_52 = _slots_17_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_223 = _slots_17_io_request & ~_GEN_221 & (|_can_allocate_T_52);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_224 = _GEN_223 & ~_GEN_216;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_225 = _GEN_223 | _GEN_216;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_226 =
    _slots_17_io_request
    & ~(_slots_17_io_request & (|_can_allocate_T_52) & ~_GEN_216 | _GEN_221)
    & (|(_slots_17_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_227 = _GEN_226 & ~_GEN_219;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_17_grant = _GEN_227 | _GEN_224 | _GEN_221;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_228 = _GEN_226 | _GEN_219;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_229 =
    _slots_18_io_request & (|(_slots_18_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_230 = _GEN_229 & ~_GEN_222;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_231 = _GEN_229 | _GEN_222;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_55 = _slots_18_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_232 = _slots_18_io_request & ~_GEN_230 & (|_can_allocate_T_55);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_233 = _GEN_232 & ~_GEN_225;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_234 = _GEN_232 | _GEN_225;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_235 =
    _slots_18_io_request
    & ~(_slots_18_io_request & (|_can_allocate_T_55) & ~_GEN_225 | _GEN_230)
    & (|(_slots_18_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_236 = _GEN_235 & ~_GEN_228;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_18_grant = _GEN_236 | _GEN_233 | _GEN_230;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_237 = _GEN_235 | _GEN_228;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_238 =
    _slots_19_io_request & (|(_slots_19_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_239 = _GEN_238 & ~_GEN_231;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_240 = _GEN_238 | _GEN_231;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_58 = _slots_19_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_241 = _slots_19_io_request & ~_GEN_239 & (|_can_allocate_T_58);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_242 = _GEN_241 & ~_GEN_234;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_243 = _GEN_241 | _GEN_234;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_244 =
    _slots_19_io_request
    & ~(_slots_19_io_request & (|_can_allocate_T_58) & ~_GEN_234 | _GEN_239)
    & (|(_slots_19_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_245 = _GEN_244 & ~_GEN_237;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_19_grant = _GEN_245 | _GEN_242 | _GEN_239;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_246 = _GEN_244 | _GEN_237;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_247 =
    _slots_20_io_request & (|(_slots_20_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_248 = _GEN_247 & ~_GEN_240;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_249 = _GEN_247 | _GEN_240;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_61 = _slots_20_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_250 = _slots_20_io_request & ~_GEN_248 & (|_can_allocate_T_61);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_251 = _GEN_250 & ~_GEN_243;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_252 = _GEN_250 | _GEN_243;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_253 =
    _slots_20_io_request
    & ~(_slots_20_io_request & (|_can_allocate_T_61) & ~_GEN_243 | _GEN_248)
    & (|(_slots_20_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_254 = _GEN_253 & ~_GEN_246;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_20_grant = _GEN_254 | _GEN_251 | _GEN_248;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_255 = _GEN_253 | _GEN_246;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_256 =
    _slots_21_io_request & (|(_slots_21_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_257 = _GEN_256 & ~_GEN_249;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_258 = _GEN_256 | _GEN_249;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_64 = _slots_21_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_259 = _slots_21_io_request & ~_GEN_257 & (|_can_allocate_T_64);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_260 = _GEN_259 & ~_GEN_252;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_261 = _GEN_259 | _GEN_252;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_262 =
    _slots_21_io_request
    & ~(_slots_21_io_request & (|_can_allocate_T_64) & ~_GEN_252 | _GEN_257)
    & (|(_slots_21_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_263 = _GEN_262 & ~_GEN_255;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_21_grant = _GEN_263 | _GEN_260 | _GEN_257;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_264 = _GEN_262 | _GEN_255;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_265 =
    _slots_22_io_request & (|(_slots_22_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_266 = _GEN_265 & ~_GEN_258;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_267 = _GEN_265 | _GEN_258;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_67 = _slots_22_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_268 = _slots_22_io_request & ~_GEN_266 & (|_can_allocate_T_67);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_269 = _GEN_268 & ~_GEN_261;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_270 = _GEN_268 | _GEN_261;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_271 =
    _slots_22_io_request
    & ~(_slots_22_io_request & (|_can_allocate_T_67) & ~_GEN_261 | _GEN_266)
    & (|(_slots_22_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_272 = _GEN_271 & ~_GEN_264;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_22_grant = _GEN_272 | _GEN_269 | _GEN_266;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_273 = _GEN_271 | _GEN_264;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_274 =
    _slots_23_io_request & (|(_slots_23_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_275 = _GEN_274 & ~_GEN_267;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_276 = _GEN_274 | _GEN_267;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_70 = _slots_23_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_277 = _slots_23_io_request & ~_GEN_275 & (|_can_allocate_T_70);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_278 = _GEN_277 & ~_GEN_270;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_279 = _GEN_277 | _GEN_270;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_280 =
    _slots_23_io_request
    & ~(_slots_23_io_request & (|_can_allocate_T_70) & ~_GEN_270 | _GEN_275)
    & (|(_slots_23_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_281 = _GEN_280 & ~_GEN_273;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_23_grant = _GEN_281 | _GEN_278 | _GEN_275;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_282 = _GEN_280 | _GEN_273;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_283 =
    _slots_24_io_request & (|(_slots_24_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_284 = _GEN_283 & ~_GEN_276;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_285 = _GEN_283 | _GEN_276;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_73 = _slots_24_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_286 = _slots_24_io_request & ~_GEN_284 & (|_can_allocate_T_73);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_287 = _GEN_286 & ~_GEN_279;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_288 = _GEN_286 | _GEN_279;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_289 =
    _slots_24_io_request
    & ~(_slots_24_io_request & (|_can_allocate_T_73) & ~_GEN_279 | _GEN_284)
    & (|(_slots_24_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_290 = _GEN_289 & ~_GEN_282;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_24_grant = _GEN_290 | _GEN_287 | _GEN_284;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_291 = _GEN_289 | _GEN_282;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_292 =
    _slots_25_io_request & (|(_slots_25_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_293 = _GEN_292 & ~_GEN_285;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_294 = _GEN_292 | _GEN_285;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_76 = _slots_25_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_295 = _slots_25_io_request & ~_GEN_293 & (|_can_allocate_T_76);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_296 = _GEN_295 & ~_GEN_288;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_297 = _GEN_295 | _GEN_288;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_298 =
    _slots_25_io_request
    & ~(_slots_25_io_request & (|_can_allocate_T_76) & ~_GEN_288 | _GEN_293)
    & (|(_slots_25_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_299 = _GEN_298 & ~_GEN_291;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_25_grant = _GEN_299 | _GEN_296 | _GEN_293;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_300 = _GEN_298 | _GEN_291;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_301 =
    _slots_26_io_request & (|(_slots_26_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_302 = _GEN_301 & ~_GEN_294;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_303 = _GEN_301 | _GEN_294;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_79 = _slots_26_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_304 = _slots_26_io_request & ~_GEN_302 & (|_can_allocate_T_79);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_305 = _GEN_304 & ~_GEN_297;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_306 = _GEN_304 | _GEN_297;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_307 =
    _slots_26_io_request
    & ~(_slots_26_io_request & (|_can_allocate_T_79) & ~_GEN_297 | _GEN_302)
    & (|(_slots_26_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_308 = _GEN_307 & ~_GEN_300;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_26_grant = _GEN_308 | _GEN_305 | _GEN_302;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_309 = _GEN_307 | _GEN_300;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_310 =
    _slots_27_io_request & (|(_slots_27_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_311 = _GEN_310 & ~_GEN_303;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_312 = _GEN_310 | _GEN_303;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_82 = _slots_27_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_313 = _slots_27_io_request & ~_GEN_311 & (|_can_allocate_T_82);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_314 = _GEN_313 & ~_GEN_306;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_315 = _GEN_313 | _GEN_306;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_316 =
    _slots_27_io_request
    & ~(_slots_27_io_request & (|_can_allocate_T_82) & ~_GEN_306 | _GEN_311)
    & (|(_slots_27_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_317 = _GEN_316 & ~_GEN_309;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_27_grant = _GEN_317 | _GEN_314 | _GEN_311;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_318 = _GEN_316 | _GEN_309;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_319 =
    _slots_28_io_request & (|(_slots_28_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_320 = _GEN_319 & ~_GEN_312;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_321 = _GEN_319 | _GEN_312;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_85 = _slots_28_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_322 = _slots_28_io_request & ~_GEN_320 & (|_can_allocate_T_85);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_323 = _GEN_322 & ~_GEN_315;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_324 = _GEN_322 | _GEN_315;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_325 =
    _slots_28_io_request
    & ~(_slots_28_io_request & (|_can_allocate_T_85) & ~_GEN_315 | _GEN_320)
    & (|(_slots_28_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_326 = _GEN_325 & ~_GEN_318;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_28_grant = _GEN_326 | _GEN_323 | _GEN_320;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_327 = _GEN_325 | _GEN_318;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_328 =
    _slots_29_io_request & (|(_slots_29_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_329 = _GEN_328 & ~_GEN_321;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_330 = _GEN_328 | _GEN_321;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire [9:0]  _can_allocate_T_88 = _slots_29_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_331 = _slots_29_io_request & ~_GEN_329 & (|_can_allocate_T_88);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_332 = _GEN_331 & ~_GEN_324;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_333 = _GEN_331 | _GEN_324;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_334 =
    _slots_29_io_request
    & ~(_slots_29_io_request & (|_can_allocate_T_88) & ~_GEN_324 | _GEN_329)
    & (|(_slots_29_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_335 = _GEN_334 & ~_GEN_327;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_29_grant = _GEN_335 | _GEN_332 | _GEN_329;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_336 = _GEN_334 | _GEN_327;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_337 =
    _slots_30_io_request & (|(_slots_30_io_uop_fu_code & io_fu_types_0));	// issue-unit-age-ordered.scala:116:{54,72}, :118:40, issue-unit.scala:153:73
  wire        _GEN_338 = _GEN_337 & ~_GEN_330;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire [9:0]  _can_allocate_T_91 = _slots_30_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_339 = _slots_30_io_request & ~_GEN_338 & (|_can_allocate_T_91);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56}, issue-unit.scala:153:73
  wire        _GEN_340 = _GEN_339 & ~_GEN_333;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  wire        _GEN_341 = _GEN_339 | _GEN_333;	// issue-unit-age-ordered.scala:118:40, :124:69
  wire        _GEN_342 =
    _slots_30_io_request
    & ~(_slots_30_io_request & (|_can_allocate_T_91) & ~_GEN_333 | _GEN_338)
    & (|(_slots_30_io_uop_fu_code & io_fu_types_2));	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  wire        _GEN_343 = _GEN_342 & ~_GEN_336;	// issue-unit-age-ordered.scala:118:{40,56,59}, :124:69
  assign issue_slots_30_grant = _GEN_343 | _GEN_340 | _GEN_338;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  wire        _GEN_344 =
    _slots_31_io_request & (|(_slots_31_io_uop_fu_code & io_fu_types_0))
    & ~(_GEN_337 | _GEN_330);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{40,56,59}, :124:69, issue-unit.scala:153:73
  wire [9:0]  _can_allocate_T_94 = _slots_31_io_uop_fu_code & io_fu_types_1;	// issue-unit-age-ordered.scala:116:54, issue-unit.scala:153:73
  wire        _GEN_345 =
    _slots_31_io_request & ~_GEN_344 & (|_can_allocate_T_94) & ~_GEN_341;	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,56,59}, :124:69, issue-unit.scala:153:73
  wire        _GEN_346 =
    _slots_31_io_request
    & ~(_slots_31_io_request & (|_can_allocate_T_94) & ~_GEN_341 | _GEN_344)
    & (|(_slots_31_io_uop_fu_code & io_fu_types_2)) & ~(_GEN_342 | _GEN_336);	// issue-unit-age-ordered.scala:116:{54,72}, :118:{28,40,56,59}, :124:69, :125:{49,74}, issue-unit.scala:153:73
  assign issue_slots_31_grant = _GEN_346 | _GEN_345 | _GEN_344;	// issue-unit-age-ordered.scala:118:{56,76}, :119:30
  always @(posedge clock) begin
    automatic logic [5:0] num_available =
      {1'h0,
       {1'h0,
        {1'h0,
         {1'h0,
          {1'h0, ~_slots_0_io_will_be_valid & ~issue_slots_0_in_uop_valid}
            + {1'h0,
               (~_slots_1_io_will_be_valid | ~_slots_0_io_valid)
                 & ~issue_slots_1_in_uop_valid}}
           + {1'h0,
              {1'h0,
               (~_slots_2_io_will_be_valid | (|_next_1_1to0))
                 & ~issue_slots_2_in_uop_valid}
                + {1'h0,
                   (~_slots_3_io_will_be_valid | (|next_2))
                     & ~issue_slots_3_in_uop_valid}}}
          + {1'h0,
             {1'h0,
              {1'h0,
               (~_slots_4_io_will_be_valid | (|next_3)) & ~issue_slots_4_in_uop_valid}
                + {1'h0,
                   (~_slots_5_io_will_be_valid | (|next_4))
                     & ~issue_slots_5_in_uop_valid}}
               + {1'h0,
                  {1'h0,
                   (~_slots_6_io_will_be_valid | (|next_5)) & ~issue_slots_6_in_uop_valid}
                    + {1'h0,
                       (~_slots_7_io_will_be_valid | (|next_6))
                         & ~issue_slots_7_in_uop_valid}}}}
         + {1'h0,
            {1'h0,
             {1'h0,
              {1'h0,
               (~_slots_8_io_will_be_valid | (|next_7)) & ~issue_slots_8_in_uop_valid}
                + {1'h0,
                   (~_slots_9_io_will_be_valid | (|next_8))
                     & ~issue_slots_9_in_uop_valid}}
               + {1'h0,
                  {1'h0,
                   (~_slots_10_io_will_be_valid | (|next_9))
                     & ~issue_slots_10_in_uop_valid}
                    + {1'h0,
                       (~_slots_11_io_will_be_valid | (|next_10))
                         & ~issue_slots_11_in_uop_valid}}}
              + {1'h0,
                 {1'h0,
                  {1'h0,
                   (~_slots_12_io_will_be_valid | (|next_11))
                     & ~issue_slots_12_in_uop_valid}
                    + {1'h0,
                       (~_slots_13_io_will_be_valid | (|next_12))
                         & ~issue_slots_13_in_uop_valid}}
                   + {1'h0,
                      {1'h0,
                       (~_slots_14_io_will_be_valid | (|next_13))
                         & ~issue_slots_14_in_uop_valid}
                        + {1'h0,
                           (~_slots_15_io_will_be_valid | (|next_14))
                             & ~issue_slots_15_in_uop_valid}}}}}
      + {1'h0,
         {1'h0,
          {1'h0,
           {1'h0,
            {1'h0,
             (~_slots_16_io_will_be_valid | (|next_15)) & ~issue_slots_16_in_uop_valid}
              + {1'h0,
                 (~_slots_17_io_will_be_valid | (|next_16))
                   & ~issue_slots_17_in_uop_valid}}
             + {1'h0,
                {1'h0,
                 (~_slots_18_io_will_be_valid | (|next_17))
                   & ~issue_slots_18_in_uop_valid}
                  + {1'h0,
                     (~_slots_19_io_will_be_valid | (|next_18))
                       & ~issue_slots_19_in_uop_valid}}}
            + {1'h0,
               {1'h0,
                {1'h0,
                 (~_slots_20_io_will_be_valid | (|next_19))
                   & ~issue_slots_20_in_uop_valid}
                  + {1'h0,
                     (~_slots_21_io_will_be_valid | (|next_20))
                       & ~issue_slots_21_in_uop_valid}}
                 + {1'h0,
                    {1'h0,
                     (~_slots_22_io_will_be_valid | (|next_21))
                       & ~issue_slots_22_in_uop_valid}
                      + {1'h0,
                         (~_slots_23_io_will_be_valid | (|next_22))
                           & ~issue_slots_23_in_uop_valid}}}}
           + {1'h0,
              {1'h0,
               {1'h0,
                {1'h0,
                 (~_slots_24_io_will_be_valid | (|next_23))
                   & ~issue_slots_24_in_uop_valid}
                  + {1'h0,
                     (~_slots_25_io_will_be_valid | (|next_24))
                       & ~issue_slots_25_in_uop_valid}}
                 + {1'h0,
                    {1'h0,
                     (~_slots_26_io_will_be_valid | (|next_25))
                       & ~issue_slots_26_in_uop_valid}
                      + {1'h0,
                         (~_slots_27_io_will_be_valid | (|next_26))
                           & ~issue_slots_27_in_uop_valid}}}
                + {1'h0,
                   {1'h0,
                    {1'h0,
                     (~_slots_28_io_will_be_valid | (|next_27))
                       & ~issue_slots_28_in_uop_valid}
                      + {1'h0,
                         (~_slots_29_io_will_be_valid | (|next_28))
                           & ~issue_slots_29_in_uop_valid}}
                     + {1'h0,
                        {1'h0,
                         (~_slots_30_io_will_be_valid | (|next_29))
                           & ~issue_slots_30_in_uop_valid}
                          + {1'h0,
                             (~_slots_31_io_will_be_valid | (|next_30))
                               & ~issue_slots_31_in_uop_valid}}}}};	// Bitwise.scala:47:55, issue-unit-age-ordered.scala:39:38, :45:37, :46:13, :47:44, :71:48, :72:37, :76:49, :84:{30,60,85,88}, issue-unit.scala:153:73
    io_dis_uops_0_ready_REG <= |num_available;	// Bitwise.scala:47:55, issue-unit-age-ordered.scala:87:{36,51}
    io_dis_uops_1_ready_REG <= |(num_available[5:1]);	// Bitwise.scala:47:55, issue-unit-age-ordered.scala:87:{36,51}
    io_dis_uops_2_ready_REG <= num_available > 6'h2;	// Bitwise.scala:47:55, issue-unit-age-ordered.scala:87:{36,51}
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:0];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        _RANDOM[/*Zero width*/ 1'b0] = `RANDOM;
        io_dis_uops_0_ready_REG = _RANDOM[/*Zero width*/ 1'b0][0];	// issue-unit-age-ordered.scala:87:36
        io_dis_uops_1_ready_REG = _RANDOM[/*Zero width*/ 1'b0][1];	// issue-unit-age-ordered.scala:87:36
        io_dis_uops_2_ready_REG = _RANDOM[/*Zero width*/ 1'b0][2];	// issue-unit-age-ordered.scala:87:36
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  IssueSlot_120 slots_0 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_0_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (1'h0),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_0_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_9
         ? _slots_3_io_out_uop_uopc
         : _GEN_8 ? _slots_2_io_out_uop_uopc : _slots_1_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_9
         ? _slots_3_io_out_uop_inst
         : _GEN_8 ? _slots_2_io_out_uop_inst : _slots_1_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_9
         ? _slots_3_io_out_uop_debug_inst
         : _GEN_8 ? _slots_2_io_out_uop_debug_inst : _slots_1_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_9
         ? _slots_3_io_out_uop_is_rvc
         : _GEN_8 ? _slots_2_io_out_uop_is_rvc : _slots_1_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_9
         ? _slots_3_io_out_uop_debug_pc
         : _GEN_8 ? _slots_2_io_out_uop_debug_pc : _slots_1_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_9
         ? _slots_3_io_out_uop_iq_type
         : _GEN_8 ? _slots_2_io_out_uop_iq_type : _slots_1_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_9
         ? _slots_3_io_out_uop_fu_code
         : _GEN_8 ? _slots_2_io_out_uop_fu_code : _slots_1_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_9
         ? _slots_3_io_out_uop_iw_state
         : _GEN_8 ? _slots_2_io_out_uop_iw_state : _slots_1_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_9
         ? _slots_3_io_out_uop_iw_p1_poisoned
         : _GEN_8
             ? _slots_2_io_out_uop_iw_p1_poisoned
             : _slots_1_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_9
         ? _slots_3_io_out_uop_iw_p2_poisoned
         : _GEN_8
             ? _slots_2_io_out_uop_iw_p2_poisoned
             : _slots_1_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_9
         ? _slots_3_io_out_uop_is_br
         : _GEN_8 ? _slots_2_io_out_uop_is_br : _slots_1_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_9
         ? _slots_3_io_out_uop_is_jalr
         : _GEN_8 ? _slots_2_io_out_uop_is_jalr : _slots_1_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_9
         ? _slots_3_io_out_uop_is_jal
         : _GEN_8 ? _slots_2_io_out_uop_is_jal : _slots_1_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_9
         ? _slots_3_io_out_uop_is_sfb
         : _GEN_8 ? _slots_2_io_out_uop_is_sfb : _slots_1_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_9
         ? _slots_3_io_out_uop_br_mask
         : _GEN_8 ? _slots_2_io_out_uop_br_mask : _slots_1_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_9
         ? _slots_3_io_out_uop_br_tag
         : _GEN_8 ? _slots_2_io_out_uop_br_tag : _slots_1_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_9
         ? _slots_3_io_out_uop_ftq_idx
         : _GEN_8 ? _slots_2_io_out_uop_ftq_idx : _slots_1_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_9
         ? _slots_3_io_out_uop_edge_inst
         : _GEN_8 ? _slots_2_io_out_uop_edge_inst : _slots_1_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_9
         ? _slots_3_io_out_uop_pc_lob
         : _GEN_8 ? _slots_2_io_out_uop_pc_lob : _slots_1_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_9
         ? _slots_3_io_out_uop_taken
         : _GEN_8 ? _slots_2_io_out_uop_taken : _slots_1_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_9
         ? _slots_3_io_out_uop_imm_packed
         : _GEN_8 ? _slots_2_io_out_uop_imm_packed : _slots_1_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_9
         ? _slots_3_io_out_uop_csr_addr
         : _GEN_8 ? _slots_2_io_out_uop_csr_addr : _slots_1_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_9
         ? _slots_3_io_out_uop_rob_idx
         : _GEN_8 ? _slots_2_io_out_uop_rob_idx : _slots_1_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_9
         ? _slots_3_io_out_uop_ldq_idx
         : _GEN_8 ? _slots_2_io_out_uop_ldq_idx : _slots_1_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_9
         ? _slots_3_io_out_uop_stq_idx
         : _GEN_8 ? _slots_2_io_out_uop_stq_idx : _slots_1_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_9
         ? _slots_3_io_out_uop_rxq_idx
         : _GEN_8 ? _slots_2_io_out_uop_rxq_idx : _slots_1_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_9
         ? _slots_3_io_out_uop_pdst
         : _GEN_8 ? _slots_2_io_out_uop_pdst : _slots_1_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_9
         ? _slots_3_io_out_uop_prs1
         : _GEN_8 ? _slots_2_io_out_uop_prs1 : _slots_1_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_9
         ? _slots_3_io_out_uop_prs2
         : _GEN_8 ? _slots_2_io_out_uop_prs2 : _slots_1_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_9
         ? _slots_3_io_out_uop_prs3
         : _GEN_8 ? _slots_2_io_out_uop_prs3 : _slots_1_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_9
         ? _slots_3_io_out_uop_ppred
         : _GEN_8 ? _slots_2_io_out_uop_ppred : _slots_1_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_9
         ? _slots_3_io_out_uop_prs1_busy
         : _GEN_8 ? _slots_2_io_out_uop_prs1_busy : _slots_1_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_9
         ? _slots_3_io_out_uop_prs2_busy
         : _GEN_8 ? _slots_2_io_out_uop_prs2_busy : _slots_1_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_9
         ? _slots_3_io_out_uop_prs3_busy
         : _GEN_8 ? _slots_2_io_out_uop_prs3_busy : _slots_1_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_9
         ? _slots_3_io_out_uop_ppred_busy
         : _GEN_8 ? _slots_2_io_out_uop_ppred_busy : _slots_1_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_9
         ? _slots_3_io_out_uop_stale_pdst
         : _GEN_8 ? _slots_2_io_out_uop_stale_pdst : _slots_1_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_9
         ? _slots_3_io_out_uop_exception
         : _GEN_8 ? _slots_2_io_out_uop_exception : _slots_1_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_9
         ? _slots_3_io_out_uop_exc_cause
         : _GEN_8 ? _slots_2_io_out_uop_exc_cause : _slots_1_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_9
         ? _slots_3_io_out_uop_bypassable
         : _GEN_8 ? _slots_2_io_out_uop_bypassable : _slots_1_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_9
         ? _slots_3_io_out_uop_mem_cmd
         : _GEN_8 ? _slots_2_io_out_uop_mem_cmd : _slots_1_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_9
         ? _slots_3_io_out_uop_mem_size
         : _GEN_8 ? _slots_2_io_out_uop_mem_size : _slots_1_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_9
         ? _slots_3_io_out_uop_mem_signed
         : _GEN_8 ? _slots_2_io_out_uop_mem_signed : _slots_1_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_9
         ? _slots_3_io_out_uop_is_fence
         : _GEN_8 ? _slots_2_io_out_uop_is_fence : _slots_1_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_9
         ? _slots_3_io_out_uop_is_fencei
         : _GEN_8 ? _slots_2_io_out_uop_is_fencei : _slots_1_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_9
         ? _slots_3_io_out_uop_is_amo
         : _GEN_8 ? _slots_2_io_out_uop_is_amo : _slots_1_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_9
         ? _slots_3_io_out_uop_uses_ldq
         : _GEN_8 ? _slots_2_io_out_uop_uses_ldq : _slots_1_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_9
         ? _slots_3_io_out_uop_uses_stq
         : _GEN_8 ? _slots_2_io_out_uop_uses_stq : _slots_1_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_9
         ? _slots_3_io_out_uop_is_sys_pc2epc
         : _GEN_8
             ? _slots_2_io_out_uop_is_sys_pc2epc
             : _slots_1_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_9
         ? _slots_3_io_out_uop_is_unique
         : _GEN_8 ? _slots_2_io_out_uop_is_unique : _slots_1_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_9
         ? _slots_3_io_out_uop_flush_on_commit
         : _GEN_8
             ? _slots_2_io_out_uop_flush_on_commit
             : _slots_1_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_9
         ? _slots_3_io_out_uop_ldst_is_rs1
         : _GEN_8 ? _slots_2_io_out_uop_ldst_is_rs1 : _slots_1_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_9
         ? _slots_3_io_out_uop_ldst
         : _GEN_8 ? _slots_2_io_out_uop_ldst : _slots_1_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_9
         ? _slots_3_io_out_uop_lrs1
         : _GEN_8 ? _slots_2_io_out_uop_lrs1 : _slots_1_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_9
         ? _slots_3_io_out_uop_lrs2
         : _GEN_8 ? _slots_2_io_out_uop_lrs2 : _slots_1_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_9
         ? _slots_3_io_out_uop_lrs3
         : _GEN_8 ? _slots_2_io_out_uop_lrs3 : _slots_1_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_9
         ? _slots_3_io_out_uop_ldst_val
         : _GEN_8 ? _slots_2_io_out_uop_ldst_val : _slots_1_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_9
         ? _slots_3_io_out_uop_dst_rtype
         : _GEN_8 ? _slots_2_io_out_uop_dst_rtype : _slots_1_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_9
         ? _slots_3_io_out_uop_lrs1_rtype
         : _GEN_8 ? _slots_2_io_out_uop_lrs1_rtype : _slots_1_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_9
         ? _slots_3_io_out_uop_lrs2_rtype
         : _GEN_8 ? _slots_2_io_out_uop_lrs2_rtype : _slots_1_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_9
         ? _slots_3_io_out_uop_frs3_en
         : _GEN_8 ? _slots_2_io_out_uop_frs3_en : _slots_1_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_9
         ? _slots_3_io_out_uop_fp_val
         : _GEN_8 ? _slots_2_io_out_uop_fp_val : _slots_1_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_9
         ? _slots_3_io_out_uop_fp_single
         : _GEN_8 ? _slots_2_io_out_uop_fp_single : _slots_1_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_9
         ? _slots_3_io_out_uop_xcpt_pf_if
         : _GEN_8 ? _slots_2_io_out_uop_xcpt_pf_if : _slots_1_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_9
         ? _slots_3_io_out_uop_xcpt_ae_if
         : _GEN_8 ? _slots_2_io_out_uop_xcpt_ae_if : _slots_1_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_9
         ? _slots_3_io_out_uop_xcpt_ma_if
         : _GEN_8 ? _slots_2_io_out_uop_xcpt_ma_if : _slots_1_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_9
         ? _slots_3_io_out_uop_bp_debug_if
         : _GEN_8 ? _slots_2_io_out_uop_bp_debug_if : _slots_1_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_9
         ? _slots_3_io_out_uop_bp_xcpt_if
         : _GEN_8 ? _slots_2_io_out_uop_bp_xcpt_if : _slots_1_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_9
         ? _slots_3_io_out_uop_debug_fsrc
         : _GEN_8 ? _slots_2_io_out_uop_debug_fsrc : _slots_1_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_9
         ? _slots_3_io_out_uop_debug_tsrc
         : _GEN_8 ? _slots_2_io_out_uop_debug_tsrc : _slots_1_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_0_io_valid),
    .io_will_be_valid               (_slots_0_io_will_be_valid),
    .io_request                     (_slots_0_io_request),
    .io_out_uop_uopc                (/* unused */),
    .io_out_uop_inst                (/* unused */),
    .io_out_uop_debug_inst          (/* unused */),
    .io_out_uop_is_rvc              (/* unused */),
    .io_out_uop_debug_pc            (/* unused */),
    .io_out_uop_iq_type             (/* unused */),
    .io_out_uop_fu_code             (/* unused */),
    .io_out_uop_iw_state            (/* unused */),
    .io_out_uop_iw_p1_poisoned      (/* unused */),
    .io_out_uop_iw_p2_poisoned      (/* unused */),
    .io_out_uop_is_br               (/* unused */),
    .io_out_uop_is_jalr             (/* unused */),
    .io_out_uop_is_jal              (/* unused */),
    .io_out_uop_is_sfb              (/* unused */),
    .io_out_uop_br_mask             (/* unused */),
    .io_out_uop_br_tag              (/* unused */),
    .io_out_uop_ftq_idx             (/* unused */),
    .io_out_uop_edge_inst           (/* unused */),
    .io_out_uop_pc_lob              (/* unused */),
    .io_out_uop_taken               (/* unused */),
    .io_out_uop_imm_packed          (/* unused */),
    .io_out_uop_csr_addr            (/* unused */),
    .io_out_uop_rob_idx             (/* unused */),
    .io_out_uop_ldq_idx             (/* unused */),
    .io_out_uop_stq_idx             (/* unused */),
    .io_out_uop_rxq_idx             (/* unused */),
    .io_out_uop_pdst                (/* unused */),
    .io_out_uop_prs1                (/* unused */),
    .io_out_uop_prs2                (/* unused */),
    .io_out_uop_prs3                (/* unused */),
    .io_out_uop_ppred               (/* unused */),
    .io_out_uop_prs1_busy           (/* unused */),
    .io_out_uop_prs2_busy           (/* unused */),
    .io_out_uop_prs3_busy           (/* unused */),
    .io_out_uop_ppred_busy          (/* unused */),
    .io_out_uop_stale_pdst          (/* unused */),
    .io_out_uop_exception           (/* unused */),
    .io_out_uop_exc_cause           (/* unused */),
    .io_out_uop_bypassable          (/* unused */),
    .io_out_uop_mem_cmd             (/* unused */),
    .io_out_uop_mem_size            (/* unused */),
    .io_out_uop_mem_signed          (/* unused */),
    .io_out_uop_is_fence            (/* unused */),
    .io_out_uop_is_fencei           (/* unused */),
    .io_out_uop_is_amo              (/* unused */),
    .io_out_uop_uses_ldq            (/* unused */),
    .io_out_uop_uses_stq            (/* unused */),
    .io_out_uop_is_sys_pc2epc       (/* unused */),
    .io_out_uop_is_unique           (/* unused */),
    .io_out_uop_flush_on_commit     (/* unused */),
    .io_out_uop_ldst_is_rs1         (/* unused */),
    .io_out_uop_ldst                (/* unused */),
    .io_out_uop_lrs1                (/* unused */),
    .io_out_uop_lrs2                (/* unused */),
    .io_out_uop_lrs3                (/* unused */),
    .io_out_uop_ldst_val            (/* unused */),
    .io_out_uop_dst_rtype           (/* unused */),
    .io_out_uop_lrs1_rtype          (/* unused */),
    .io_out_uop_lrs2_rtype          (/* unused */),
    .io_out_uop_frs3_en             (/* unused */),
    .io_out_uop_fp_val              (/* unused */),
    .io_out_uop_fp_single           (/* unused */),
    .io_out_uop_xcpt_pf_if          (/* unused */),
    .io_out_uop_xcpt_ae_if          (/* unused */),
    .io_out_uop_xcpt_ma_if          (/* unused */),
    .io_out_uop_bp_debug_if         (/* unused */),
    .io_out_uop_bp_xcpt_if          (/* unused */),
    .io_out_uop_debug_fsrc          (/* unused */),
    .io_out_uop_debug_tsrc          (/* unused */),
    .io_uop_uopc                    (_slots_0_io_uop_uopc),
    .io_uop_inst                    (_slots_0_io_uop_inst),
    .io_uop_debug_inst              (_slots_0_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_0_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_0_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_0_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_0_io_uop_fu_code),
    .io_uop_iw_state                (_slots_0_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_0_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_0_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_0_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_0_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_0_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_0_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_0_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_0_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_0_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_0_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_0_io_uop_pc_lob),
    .io_uop_taken                   (_slots_0_io_uop_taken),
    .io_uop_imm_packed              (_slots_0_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_0_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_0_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_0_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_0_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_0_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_0_io_uop_pdst),
    .io_uop_prs1                    (_slots_0_io_uop_prs1),
    .io_uop_prs2                    (_slots_0_io_uop_prs2),
    .io_uop_prs3                    (_slots_0_io_uop_prs3),
    .io_uop_ppred                   (_slots_0_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_0_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_0_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_0_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_0_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_0_io_uop_stale_pdst),
    .io_uop_exception               (_slots_0_io_uop_exception),
    .io_uop_exc_cause               (_slots_0_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_0_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_0_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_0_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_0_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_0_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_0_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_0_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_0_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_0_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_0_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_0_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_0_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_0_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_0_io_uop_ldst),
    .io_uop_lrs1                    (_slots_0_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_0_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_0_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_0_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_0_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_0_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_0_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_0_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_0_io_uop_fp_val),
    .io_uop_fp_single               (_slots_0_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_0_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_0_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_0_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_0_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_0_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_0_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_0_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_1 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_1_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (~_slots_0_io_valid),	// issue-unit-age-ordered.scala:39:38, issue-unit.scala:153:73
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_1_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_11
         ? _slots_4_io_out_uop_uopc
         : _GEN_10 ? _slots_3_io_out_uop_uopc : _slots_2_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_11
         ? _slots_4_io_out_uop_inst
         : _GEN_10 ? _slots_3_io_out_uop_inst : _slots_2_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_11
         ? _slots_4_io_out_uop_debug_inst
         : _GEN_10 ? _slots_3_io_out_uop_debug_inst : _slots_2_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_11
         ? _slots_4_io_out_uop_is_rvc
         : _GEN_10 ? _slots_3_io_out_uop_is_rvc : _slots_2_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_11
         ? _slots_4_io_out_uop_debug_pc
         : _GEN_10 ? _slots_3_io_out_uop_debug_pc : _slots_2_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_11
         ? _slots_4_io_out_uop_iq_type
         : _GEN_10 ? _slots_3_io_out_uop_iq_type : _slots_2_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_11
         ? _slots_4_io_out_uop_fu_code
         : _GEN_10 ? _slots_3_io_out_uop_fu_code : _slots_2_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_11
         ? _slots_4_io_out_uop_iw_state
         : _GEN_10 ? _slots_3_io_out_uop_iw_state : _slots_2_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_11
         ? _slots_4_io_out_uop_iw_p1_poisoned
         : _GEN_10
             ? _slots_3_io_out_uop_iw_p1_poisoned
             : _slots_2_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_11
         ? _slots_4_io_out_uop_iw_p2_poisoned
         : _GEN_10
             ? _slots_3_io_out_uop_iw_p2_poisoned
             : _slots_2_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_11
         ? _slots_4_io_out_uop_is_br
         : _GEN_10 ? _slots_3_io_out_uop_is_br : _slots_2_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_11
         ? _slots_4_io_out_uop_is_jalr
         : _GEN_10 ? _slots_3_io_out_uop_is_jalr : _slots_2_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_11
         ? _slots_4_io_out_uop_is_jal
         : _GEN_10 ? _slots_3_io_out_uop_is_jal : _slots_2_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_11
         ? _slots_4_io_out_uop_is_sfb
         : _GEN_10 ? _slots_3_io_out_uop_is_sfb : _slots_2_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_11
         ? _slots_4_io_out_uop_br_mask
         : _GEN_10 ? _slots_3_io_out_uop_br_mask : _slots_2_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_11
         ? _slots_4_io_out_uop_br_tag
         : _GEN_10 ? _slots_3_io_out_uop_br_tag : _slots_2_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_11
         ? _slots_4_io_out_uop_ftq_idx
         : _GEN_10 ? _slots_3_io_out_uop_ftq_idx : _slots_2_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_11
         ? _slots_4_io_out_uop_edge_inst
         : _GEN_10 ? _slots_3_io_out_uop_edge_inst : _slots_2_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_11
         ? _slots_4_io_out_uop_pc_lob
         : _GEN_10 ? _slots_3_io_out_uop_pc_lob : _slots_2_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_11
         ? _slots_4_io_out_uop_taken
         : _GEN_10 ? _slots_3_io_out_uop_taken : _slots_2_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_11
         ? _slots_4_io_out_uop_imm_packed
         : _GEN_10 ? _slots_3_io_out_uop_imm_packed : _slots_2_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_11
         ? _slots_4_io_out_uop_csr_addr
         : _GEN_10 ? _slots_3_io_out_uop_csr_addr : _slots_2_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_11
         ? _slots_4_io_out_uop_rob_idx
         : _GEN_10 ? _slots_3_io_out_uop_rob_idx : _slots_2_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_11
         ? _slots_4_io_out_uop_ldq_idx
         : _GEN_10 ? _slots_3_io_out_uop_ldq_idx : _slots_2_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_11
         ? _slots_4_io_out_uop_stq_idx
         : _GEN_10 ? _slots_3_io_out_uop_stq_idx : _slots_2_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_11
         ? _slots_4_io_out_uop_rxq_idx
         : _GEN_10 ? _slots_3_io_out_uop_rxq_idx : _slots_2_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_11
         ? _slots_4_io_out_uop_pdst
         : _GEN_10 ? _slots_3_io_out_uop_pdst : _slots_2_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_11
         ? _slots_4_io_out_uop_prs1
         : _GEN_10 ? _slots_3_io_out_uop_prs1 : _slots_2_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_11
         ? _slots_4_io_out_uop_prs2
         : _GEN_10 ? _slots_3_io_out_uop_prs2 : _slots_2_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_11
         ? _slots_4_io_out_uop_prs3
         : _GEN_10 ? _slots_3_io_out_uop_prs3 : _slots_2_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_11
         ? _slots_4_io_out_uop_ppred
         : _GEN_10 ? _slots_3_io_out_uop_ppred : _slots_2_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_11
         ? _slots_4_io_out_uop_prs1_busy
         : _GEN_10 ? _slots_3_io_out_uop_prs1_busy : _slots_2_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_11
         ? _slots_4_io_out_uop_prs2_busy
         : _GEN_10 ? _slots_3_io_out_uop_prs2_busy : _slots_2_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_11
         ? _slots_4_io_out_uop_prs3_busy
         : _GEN_10 ? _slots_3_io_out_uop_prs3_busy : _slots_2_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_11
         ? _slots_4_io_out_uop_ppred_busy
         : _GEN_10 ? _slots_3_io_out_uop_ppred_busy : _slots_2_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_11
         ? _slots_4_io_out_uop_stale_pdst
         : _GEN_10 ? _slots_3_io_out_uop_stale_pdst : _slots_2_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_11
         ? _slots_4_io_out_uop_exception
         : _GEN_10 ? _slots_3_io_out_uop_exception : _slots_2_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_11
         ? _slots_4_io_out_uop_exc_cause
         : _GEN_10 ? _slots_3_io_out_uop_exc_cause : _slots_2_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_11
         ? _slots_4_io_out_uop_bypassable
         : _GEN_10 ? _slots_3_io_out_uop_bypassable : _slots_2_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_11
         ? _slots_4_io_out_uop_mem_cmd
         : _GEN_10 ? _slots_3_io_out_uop_mem_cmd : _slots_2_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_11
         ? _slots_4_io_out_uop_mem_size
         : _GEN_10 ? _slots_3_io_out_uop_mem_size : _slots_2_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_11
         ? _slots_4_io_out_uop_mem_signed
         : _GEN_10 ? _slots_3_io_out_uop_mem_signed : _slots_2_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_11
         ? _slots_4_io_out_uop_is_fence
         : _GEN_10 ? _slots_3_io_out_uop_is_fence : _slots_2_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_11
         ? _slots_4_io_out_uop_is_fencei
         : _GEN_10 ? _slots_3_io_out_uop_is_fencei : _slots_2_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_11
         ? _slots_4_io_out_uop_is_amo
         : _GEN_10 ? _slots_3_io_out_uop_is_amo : _slots_2_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_11
         ? _slots_4_io_out_uop_uses_ldq
         : _GEN_10 ? _slots_3_io_out_uop_uses_ldq : _slots_2_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_11
         ? _slots_4_io_out_uop_uses_stq
         : _GEN_10 ? _slots_3_io_out_uop_uses_stq : _slots_2_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_11
         ? _slots_4_io_out_uop_is_sys_pc2epc
         : _GEN_10
             ? _slots_3_io_out_uop_is_sys_pc2epc
             : _slots_2_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_11
         ? _slots_4_io_out_uop_is_unique
         : _GEN_10 ? _slots_3_io_out_uop_is_unique : _slots_2_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_11
         ? _slots_4_io_out_uop_flush_on_commit
         : _GEN_10
             ? _slots_3_io_out_uop_flush_on_commit
             : _slots_2_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_11
         ? _slots_4_io_out_uop_ldst_is_rs1
         : _GEN_10 ? _slots_3_io_out_uop_ldst_is_rs1 : _slots_2_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_11
         ? _slots_4_io_out_uop_ldst
         : _GEN_10 ? _slots_3_io_out_uop_ldst : _slots_2_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_11
         ? _slots_4_io_out_uop_lrs1
         : _GEN_10 ? _slots_3_io_out_uop_lrs1 : _slots_2_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_11
         ? _slots_4_io_out_uop_lrs2
         : _GEN_10 ? _slots_3_io_out_uop_lrs2 : _slots_2_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_11
         ? _slots_4_io_out_uop_lrs3
         : _GEN_10 ? _slots_3_io_out_uop_lrs3 : _slots_2_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_11
         ? _slots_4_io_out_uop_ldst_val
         : _GEN_10 ? _slots_3_io_out_uop_ldst_val : _slots_2_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_11
         ? _slots_4_io_out_uop_dst_rtype
         : _GEN_10 ? _slots_3_io_out_uop_dst_rtype : _slots_2_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_11
         ? _slots_4_io_out_uop_lrs1_rtype
         : _GEN_10 ? _slots_3_io_out_uop_lrs1_rtype : _slots_2_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_11
         ? _slots_4_io_out_uop_lrs2_rtype
         : _GEN_10 ? _slots_3_io_out_uop_lrs2_rtype : _slots_2_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_11
         ? _slots_4_io_out_uop_frs3_en
         : _GEN_10 ? _slots_3_io_out_uop_frs3_en : _slots_2_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_11
         ? _slots_4_io_out_uop_fp_val
         : _GEN_10 ? _slots_3_io_out_uop_fp_val : _slots_2_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_11
         ? _slots_4_io_out_uop_fp_single
         : _GEN_10 ? _slots_3_io_out_uop_fp_single : _slots_2_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_11
         ? _slots_4_io_out_uop_xcpt_pf_if
         : _GEN_10 ? _slots_3_io_out_uop_xcpt_pf_if : _slots_2_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_11
         ? _slots_4_io_out_uop_xcpt_ae_if
         : _GEN_10 ? _slots_3_io_out_uop_xcpt_ae_if : _slots_2_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_11
         ? _slots_4_io_out_uop_xcpt_ma_if
         : _GEN_10 ? _slots_3_io_out_uop_xcpt_ma_if : _slots_2_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_11
         ? _slots_4_io_out_uop_bp_debug_if
         : _GEN_10 ? _slots_3_io_out_uop_bp_debug_if : _slots_2_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_11
         ? _slots_4_io_out_uop_bp_xcpt_if
         : _GEN_10 ? _slots_3_io_out_uop_bp_xcpt_if : _slots_2_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_11
         ? _slots_4_io_out_uop_debug_fsrc
         : _GEN_10 ? _slots_3_io_out_uop_debug_fsrc : _slots_2_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_11
         ? _slots_4_io_out_uop_debug_tsrc
         : _GEN_10 ? _slots_3_io_out_uop_debug_tsrc : _slots_2_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_1_io_valid),
    .io_will_be_valid               (_slots_1_io_will_be_valid),
    .io_request                     (_slots_1_io_request),
    .io_out_uop_uopc                (_slots_1_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_1_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_1_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_1_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_1_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_1_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_1_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_1_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_1_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_1_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_1_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_1_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_1_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_1_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_1_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_1_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_1_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_1_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_1_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_1_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_1_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_1_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_1_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_1_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_1_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_1_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_1_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_1_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_1_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_1_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_1_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_1_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_1_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_1_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_1_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_1_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_1_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_1_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_1_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_1_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_1_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_1_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_1_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_1_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_1_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_1_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_1_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_1_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_1_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_1_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_1_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_1_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_1_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_1_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_1_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_1_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_1_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_1_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_1_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_1_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_1_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_1_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_1_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_1_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_1_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_1_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_1_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_1_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_1_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_1_io_uop_uopc),
    .io_uop_inst                    (_slots_1_io_uop_inst),
    .io_uop_debug_inst              (_slots_1_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_1_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_1_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_1_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_1_io_uop_fu_code),
    .io_uop_iw_state                (_slots_1_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_1_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_1_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_1_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_1_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_1_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_1_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_1_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_1_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_1_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_1_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_1_io_uop_pc_lob),
    .io_uop_taken                   (_slots_1_io_uop_taken),
    .io_uop_imm_packed              (_slots_1_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_1_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_1_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_1_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_1_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_1_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_1_io_uop_pdst),
    .io_uop_prs1                    (_slots_1_io_uop_prs1),
    .io_uop_prs2                    (_slots_1_io_uop_prs2),
    .io_uop_prs3                    (_slots_1_io_uop_prs3),
    .io_uop_ppred                   (_slots_1_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_1_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_1_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_1_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_1_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_1_io_uop_stale_pdst),
    .io_uop_exception               (_slots_1_io_uop_exception),
    .io_uop_exc_cause               (_slots_1_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_1_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_1_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_1_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_1_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_1_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_1_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_1_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_1_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_1_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_1_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_1_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_1_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_1_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_1_io_uop_ldst),
    .io_uop_lrs1                    (_slots_1_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_1_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_1_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_1_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_1_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_1_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_1_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_1_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_1_io_uop_fp_val),
    .io_uop_fp_single               (_slots_1_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_1_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_1_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_1_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_1_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_1_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_1_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_1_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_2 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_2_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_next_1_1to0),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_2_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_13
         ? _slots_5_io_out_uop_uopc
         : _GEN_12 ? _slots_4_io_out_uop_uopc : _slots_3_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_13
         ? _slots_5_io_out_uop_inst
         : _GEN_12 ? _slots_4_io_out_uop_inst : _slots_3_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_13
         ? _slots_5_io_out_uop_debug_inst
         : _GEN_12 ? _slots_4_io_out_uop_debug_inst : _slots_3_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_13
         ? _slots_5_io_out_uop_is_rvc
         : _GEN_12 ? _slots_4_io_out_uop_is_rvc : _slots_3_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_13
         ? _slots_5_io_out_uop_debug_pc
         : _GEN_12 ? _slots_4_io_out_uop_debug_pc : _slots_3_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_13
         ? _slots_5_io_out_uop_iq_type
         : _GEN_12 ? _slots_4_io_out_uop_iq_type : _slots_3_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_13
         ? _slots_5_io_out_uop_fu_code
         : _GEN_12 ? _slots_4_io_out_uop_fu_code : _slots_3_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_13
         ? _slots_5_io_out_uop_iw_state
         : _GEN_12 ? _slots_4_io_out_uop_iw_state : _slots_3_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_13
         ? _slots_5_io_out_uop_iw_p1_poisoned
         : _GEN_12
             ? _slots_4_io_out_uop_iw_p1_poisoned
             : _slots_3_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_13
         ? _slots_5_io_out_uop_iw_p2_poisoned
         : _GEN_12
             ? _slots_4_io_out_uop_iw_p2_poisoned
             : _slots_3_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_13
         ? _slots_5_io_out_uop_is_br
         : _GEN_12 ? _slots_4_io_out_uop_is_br : _slots_3_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_13
         ? _slots_5_io_out_uop_is_jalr
         : _GEN_12 ? _slots_4_io_out_uop_is_jalr : _slots_3_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_13
         ? _slots_5_io_out_uop_is_jal
         : _GEN_12 ? _slots_4_io_out_uop_is_jal : _slots_3_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_13
         ? _slots_5_io_out_uop_is_sfb
         : _GEN_12 ? _slots_4_io_out_uop_is_sfb : _slots_3_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_13
         ? _slots_5_io_out_uop_br_mask
         : _GEN_12 ? _slots_4_io_out_uop_br_mask : _slots_3_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_13
         ? _slots_5_io_out_uop_br_tag
         : _GEN_12 ? _slots_4_io_out_uop_br_tag : _slots_3_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_13
         ? _slots_5_io_out_uop_ftq_idx
         : _GEN_12 ? _slots_4_io_out_uop_ftq_idx : _slots_3_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_13
         ? _slots_5_io_out_uop_edge_inst
         : _GEN_12 ? _slots_4_io_out_uop_edge_inst : _slots_3_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_13
         ? _slots_5_io_out_uop_pc_lob
         : _GEN_12 ? _slots_4_io_out_uop_pc_lob : _slots_3_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_13
         ? _slots_5_io_out_uop_taken
         : _GEN_12 ? _slots_4_io_out_uop_taken : _slots_3_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_13
         ? _slots_5_io_out_uop_imm_packed
         : _GEN_12 ? _slots_4_io_out_uop_imm_packed : _slots_3_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_13
         ? _slots_5_io_out_uop_csr_addr
         : _GEN_12 ? _slots_4_io_out_uop_csr_addr : _slots_3_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_13
         ? _slots_5_io_out_uop_rob_idx
         : _GEN_12 ? _slots_4_io_out_uop_rob_idx : _slots_3_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_13
         ? _slots_5_io_out_uop_ldq_idx
         : _GEN_12 ? _slots_4_io_out_uop_ldq_idx : _slots_3_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_13
         ? _slots_5_io_out_uop_stq_idx
         : _GEN_12 ? _slots_4_io_out_uop_stq_idx : _slots_3_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_13
         ? _slots_5_io_out_uop_rxq_idx
         : _GEN_12 ? _slots_4_io_out_uop_rxq_idx : _slots_3_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_13
         ? _slots_5_io_out_uop_pdst
         : _GEN_12 ? _slots_4_io_out_uop_pdst : _slots_3_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_13
         ? _slots_5_io_out_uop_prs1
         : _GEN_12 ? _slots_4_io_out_uop_prs1 : _slots_3_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_13
         ? _slots_5_io_out_uop_prs2
         : _GEN_12 ? _slots_4_io_out_uop_prs2 : _slots_3_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_13
         ? _slots_5_io_out_uop_prs3
         : _GEN_12 ? _slots_4_io_out_uop_prs3 : _slots_3_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_13
         ? _slots_5_io_out_uop_ppred
         : _GEN_12 ? _slots_4_io_out_uop_ppred : _slots_3_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_13
         ? _slots_5_io_out_uop_prs1_busy
         : _GEN_12 ? _slots_4_io_out_uop_prs1_busy : _slots_3_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_13
         ? _slots_5_io_out_uop_prs2_busy
         : _GEN_12 ? _slots_4_io_out_uop_prs2_busy : _slots_3_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_13
         ? _slots_5_io_out_uop_prs3_busy
         : _GEN_12 ? _slots_4_io_out_uop_prs3_busy : _slots_3_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_13
         ? _slots_5_io_out_uop_ppred_busy
         : _GEN_12 ? _slots_4_io_out_uop_ppred_busy : _slots_3_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_13
         ? _slots_5_io_out_uop_stale_pdst
         : _GEN_12 ? _slots_4_io_out_uop_stale_pdst : _slots_3_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_13
         ? _slots_5_io_out_uop_exception
         : _GEN_12 ? _slots_4_io_out_uop_exception : _slots_3_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_13
         ? _slots_5_io_out_uop_exc_cause
         : _GEN_12 ? _slots_4_io_out_uop_exc_cause : _slots_3_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_13
         ? _slots_5_io_out_uop_bypassable
         : _GEN_12 ? _slots_4_io_out_uop_bypassable : _slots_3_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_13
         ? _slots_5_io_out_uop_mem_cmd
         : _GEN_12 ? _slots_4_io_out_uop_mem_cmd : _slots_3_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_13
         ? _slots_5_io_out_uop_mem_size
         : _GEN_12 ? _slots_4_io_out_uop_mem_size : _slots_3_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_13
         ? _slots_5_io_out_uop_mem_signed
         : _GEN_12 ? _slots_4_io_out_uop_mem_signed : _slots_3_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_13
         ? _slots_5_io_out_uop_is_fence
         : _GEN_12 ? _slots_4_io_out_uop_is_fence : _slots_3_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_13
         ? _slots_5_io_out_uop_is_fencei
         : _GEN_12 ? _slots_4_io_out_uop_is_fencei : _slots_3_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_13
         ? _slots_5_io_out_uop_is_amo
         : _GEN_12 ? _slots_4_io_out_uop_is_amo : _slots_3_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_13
         ? _slots_5_io_out_uop_uses_ldq
         : _GEN_12 ? _slots_4_io_out_uop_uses_ldq : _slots_3_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_13
         ? _slots_5_io_out_uop_uses_stq
         : _GEN_12 ? _slots_4_io_out_uop_uses_stq : _slots_3_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_13
         ? _slots_5_io_out_uop_is_sys_pc2epc
         : _GEN_12
             ? _slots_4_io_out_uop_is_sys_pc2epc
             : _slots_3_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_13
         ? _slots_5_io_out_uop_is_unique
         : _GEN_12 ? _slots_4_io_out_uop_is_unique : _slots_3_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_13
         ? _slots_5_io_out_uop_flush_on_commit
         : _GEN_12
             ? _slots_4_io_out_uop_flush_on_commit
             : _slots_3_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_13
         ? _slots_5_io_out_uop_ldst_is_rs1
         : _GEN_12 ? _slots_4_io_out_uop_ldst_is_rs1 : _slots_3_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_13
         ? _slots_5_io_out_uop_ldst
         : _GEN_12 ? _slots_4_io_out_uop_ldst : _slots_3_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_13
         ? _slots_5_io_out_uop_lrs1
         : _GEN_12 ? _slots_4_io_out_uop_lrs1 : _slots_3_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_13
         ? _slots_5_io_out_uop_lrs2
         : _GEN_12 ? _slots_4_io_out_uop_lrs2 : _slots_3_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_13
         ? _slots_5_io_out_uop_lrs3
         : _GEN_12 ? _slots_4_io_out_uop_lrs3 : _slots_3_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_13
         ? _slots_5_io_out_uop_ldst_val
         : _GEN_12 ? _slots_4_io_out_uop_ldst_val : _slots_3_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_13
         ? _slots_5_io_out_uop_dst_rtype
         : _GEN_12 ? _slots_4_io_out_uop_dst_rtype : _slots_3_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_13
         ? _slots_5_io_out_uop_lrs1_rtype
         : _GEN_12 ? _slots_4_io_out_uop_lrs1_rtype : _slots_3_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_13
         ? _slots_5_io_out_uop_lrs2_rtype
         : _GEN_12 ? _slots_4_io_out_uop_lrs2_rtype : _slots_3_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_13
         ? _slots_5_io_out_uop_frs3_en
         : _GEN_12 ? _slots_4_io_out_uop_frs3_en : _slots_3_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_13
         ? _slots_5_io_out_uop_fp_val
         : _GEN_12 ? _slots_4_io_out_uop_fp_val : _slots_3_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_13
         ? _slots_5_io_out_uop_fp_single
         : _GEN_12 ? _slots_4_io_out_uop_fp_single : _slots_3_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_13
         ? _slots_5_io_out_uop_xcpt_pf_if
         : _GEN_12 ? _slots_4_io_out_uop_xcpt_pf_if : _slots_3_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_13
         ? _slots_5_io_out_uop_xcpt_ae_if
         : _GEN_12 ? _slots_4_io_out_uop_xcpt_ae_if : _slots_3_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_13
         ? _slots_5_io_out_uop_xcpt_ma_if
         : _GEN_12 ? _slots_4_io_out_uop_xcpt_ma_if : _slots_3_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_13
         ? _slots_5_io_out_uop_bp_debug_if
         : _GEN_12 ? _slots_4_io_out_uop_bp_debug_if : _slots_3_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_13
         ? _slots_5_io_out_uop_bp_xcpt_if
         : _GEN_12 ? _slots_4_io_out_uop_bp_xcpt_if : _slots_3_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_13
         ? _slots_5_io_out_uop_debug_fsrc
         : _GEN_12 ? _slots_4_io_out_uop_debug_fsrc : _slots_3_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_13
         ? _slots_5_io_out_uop_debug_tsrc
         : _GEN_12 ? _slots_4_io_out_uop_debug_tsrc : _slots_3_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_2_io_valid),
    .io_will_be_valid               (_slots_2_io_will_be_valid),
    .io_request                     (_slots_2_io_request),
    .io_out_uop_uopc                (_slots_2_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_2_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_2_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_2_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_2_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_2_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_2_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_2_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_2_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_2_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_2_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_2_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_2_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_2_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_2_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_2_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_2_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_2_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_2_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_2_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_2_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_2_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_2_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_2_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_2_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_2_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_2_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_2_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_2_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_2_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_2_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_2_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_2_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_2_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_2_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_2_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_2_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_2_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_2_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_2_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_2_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_2_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_2_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_2_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_2_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_2_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_2_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_2_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_2_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_2_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_2_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_2_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_2_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_2_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_2_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_2_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_2_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_2_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_2_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_2_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_2_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_2_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_2_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_2_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_2_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_2_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_2_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_2_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_2_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_2_io_uop_uopc),
    .io_uop_inst                    (_slots_2_io_uop_inst),
    .io_uop_debug_inst              (_slots_2_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_2_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_2_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_2_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_2_io_uop_fu_code),
    .io_uop_iw_state                (_slots_2_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_2_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_2_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_2_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_2_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_2_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_2_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_2_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_2_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_2_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_2_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_2_io_uop_pc_lob),
    .io_uop_taken                   (_slots_2_io_uop_taken),
    .io_uop_imm_packed              (_slots_2_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_2_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_2_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_2_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_2_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_2_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_2_io_uop_pdst),
    .io_uop_prs1                    (_slots_2_io_uop_prs1),
    .io_uop_prs2                    (_slots_2_io_uop_prs2),
    .io_uop_prs3                    (_slots_2_io_uop_prs3),
    .io_uop_ppred                   (_slots_2_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_2_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_2_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_2_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_2_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_2_io_uop_stale_pdst),
    .io_uop_exception               (_slots_2_io_uop_exception),
    .io_uop_exc_cause               (_slots_2_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_2_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_2_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_2_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_2_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_2_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_2_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_2_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_2_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_2_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_2_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_2_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_2_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_2_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_2_io_uop_ldst),
    .io_uop_lrs1                    (_slots_2_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_2_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_2_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_2_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_2_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_2_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_2_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_2_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_2_io_uop_fp_val),
    .io_uop_fp_single               (_slots_2_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_2_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_2_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_2_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_2_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_2_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_2_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_2_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_3 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_3_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_2),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_3_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_15
         ? _slots_6_io_out_uop_uopc
         : _GEN_14 ? _slots_5_io_out_uop_uopc : _slots_4_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_15
         ? _slots_6_io_out_uop_inst
         : _GEN_14 ? _slots_5_io_out_uop_inst : _slots_4_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_15
         ? _slots_6_io_out_uop_debug_inst
         : _GEN_14 ? _slots_5_io_out_uop_debug_inst : _slots_4_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_15
         ? _slots_6_io_out_uop_is_rvc
         : _GEN_14 ? _slots_5_io_out_uop_is_rvc : _slots_4_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_15
         ? _slots_6_io_out_uop_debug_pc
         : _GEN_14 ? _slots_5_io_out_uop_debug_pc : _slots_4_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_15
         ? _slots_6_io_out_uop_iq_type
         : _GEN_14 ? _slots_5_io_out_uop_iq_type : _slots_4_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_15
         ? _slots_6_io_out_uop_fu_code
         : _GEN_14 ? _slots_5_io_out_uop_fu_code : _slots_4_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_15
         ? _slots_6_io_out_uop_iw_state
         : _GEN_14 ? _slots_5_io_out_uop_iw_state : _slots_4_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_15
         ? _slots_6_io_out_uop_iw_p1_poisoned
         : _GEN_14
             ? _slots_5_io_out_uop_iw_p1_poisoned
             : _slots_4_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_15
         ? _slots_6_io_out_uop_iw_p2_poisoned
         : _GEN_14
             ? _slots_5_io_out_uop_iw_p2_poisoned
             : _slots_4_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_15
         ? _slots_6_io_out_uop_is_br
         : _GEN_14 ? _slots_5_io_out_uop_is_br : _slots_4_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_15
         ? _slots_6_io_out_uop_is_jalr
         : _GEN_14 ? _slots_5_io_out_uop_is_jalr : _slots_4_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_15
         ? _slots_6_io_out_uop_is_jal
         : _GEN_14 ? _slots_5_io_out_uop_is_jal : _slots_4_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_15
         ? _slots_6_io_out_uop_is_sfb
         : _GEN_14 ? _slots_5_io_out_uop_is_sfb : _slots_4_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_15
         ? _slots_6_io_out_uop_br_mask
         : _GEN_14 ? _slots_5_io_out_uop_br_mask : _slots_4_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_15
         ? _slots_6_io_out_uop_br_tag
         : _GEN_14 ? _slots_5_io_out_uop_br_tag : _slots_4_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_15
         ? _slots_6_io_out_uop_ftq_idx
         : _GEN_14 ? _slots_5_io_out_uop_ftq_idx : _slots_4_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_15
         ? _slots_6_io_out_uop_edge_inst
         : _GEN_14 ? _slots_5_io_out_uop_edge_inst : _slots_4_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_15
         ? _slots_6_io_out_uop_pc_lob
         : _GEN_14 ? _slots_5_io_out_uop_pc_lob : _slots_4_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_15
         ? _slots_6_io_out_uop_taken
         : _GEN_14 ? _slots_5_io_out_uop_taken : _slots_4_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_15
         ? _slots_6_io_out_uop_imm_packed
         : _GEN_14 ? _slots_5_io_out_uop_imm_packed : _slots_4_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_15
         ? _slots_6_io_out_uop_csr_addr
         : _GEN_14 ? _slots_5_io_out_uop_csr_addr : _slots_4_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_15
         ? _slots_6_io_out_uop_rob_idx
         : _GEN_14 ? _slots_5_io_out_uop_rob_idx : _slots_4_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_15
         ? _slots_6_io_out_uop_ldq_idx
         : _GEN_14 ? _slots_5_io_out_uop_ldq_idx : _slots_4_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_15
         ? _slots_6_io_out_uop_stq_idx
         : _GEN_14 ? _slots_5_io_out_uop_stq_idx : _slots_4_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_15
         ? _slots_6_io_out_uop_rxq_idx
         : _GEN_14 ? _slots_5_io_out_uop_rxq_idx : _slots_4_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_15
         ? _slots_6_io_out_uop_pdst
         : _GEN_14 ? _slots_5_io_out_uop_pdst : _slots_4_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_15
         ? _slots_6_io_out_uop_prs1
         : _GEN_14 ? _slots_5_io_out_uop_prs1 : _slots_4_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_15
         ? _slots_6_io_out_uop_prs2
         : _GEN_14 ? _slots_5_io_out_uop_prs2 : _slots_4_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_15
         ? _slots_6_io_out_uop_prs3
         : _GEN_14 ? _slots_5_io_out_uop_prs3 : _slots_4_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_15
         ? _slots_6_io_out_uop_ppred
         : _GEN_14 ? _slots_5_io_out_uop_ppred : _slots_4_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_15
         ? _slots_6_io_out_uop_prs1_busy
         : _GEN_14 ? _slots_5_io_out_uop_prs1_busy : _slots_4_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_15
         ? _slots_6_io_out_uop_prs2_busy
         : _GEN_14 ? _slots_5_io_out_uop_prs2_busy : _slots_4_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_15
         ? _slots_6_io_out_uop_prs3_busy
         : _GEN_14 ? _slots_5_io_out_uop_prs3_busy : _slots_4_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_15
         ? _slots_6_io_out_uop_ppred_busy
         : _GEN_14 ? _slots_5_io_out_uop_ppred_busy : _slots_4_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_15
         ? _slots_6_io_out_uop_stale_pdst
         : _GEN_14 ? _slots_5_io_out_uop_stale_pdst : _slots_4_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_15
         ? _slots_6_io_out_uop_exception
         : _GEN_14 ? _slots_5_io_out_uop_exception : _slots_4_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_15
         ? _slots_6_io_out_uop_exc_cause
         : _GEN_14 ? _slots_5_io_out_uop_exc_cause : _slots_4_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_15
         ? _slots_6_io_out_uop_bypassable
         : _GEN_14 ? _slots_5_io_out_uop_bypassable : _slots_4_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_15
         ? _slots_6_io_out_uop_mem_cmd
         : _GEN_14 ? _slots_5_io_out_uop_mem_cmd : _slots_4_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_15
         ? _slots_6_io_out_uop_mem_size
         : _GEN_14 ? _slots_5_io_out_uop_mem_size : _slots_4_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_15
         ? _slots_6_io_out_uop_mem_signed
         : _GEN_14 ? _slots_5_io_out_uop_mem_signed : _slots_4_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_15
         ? _slots_6_io_out_uop_is_fence
         : _GEN_14 ? _slots_5_io_out_uop_is_fence : _slots_4_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_15
         ? _slots_6_io_out_uop_is_fencei
         : _GEN_14 ? _slots_5_io_out_uop_is_fencei : _slots_4_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_15
         ? _slots_6_io_out_uop_is_amo
         : _GEN_14 ? _slots_5_io_out_uop_is_amo : _slots_4_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_15
         ? _slots_6_io_out_uop_uses_ldq
         : _GEN_14 ? _slots_5_io_out_uop_uses_ldq : _slots_4_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_15
         ? _slots_6_io_out_uop_uses_stq
         : _GEN_14 ? _slots_5_io_out_uop_uses_stq : _slots_4_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_15
         ? _slots_6_io_out_uop_is_sys_pc2epc
         : _GEN_14
             ? _slots_5_io_out_uop_is_sys_pc2epc
             : _slots_4_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_15
         ? _slots_6_io_out_uop_is_unique
         : _GEN_14 ? _slots_5_io_out_uop_is_unique : _slots_4_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_15
         ? _slots_6_io_out_uop_flush_on_commit
         : _GEN_14
             ? _slots_5_io_out_uop_flush_on_commit
             : _slots_4_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_15
         ? _slots_6_io_out_uop_ldst_is_rs1
         : _GEN_14 ? _slots_5_io_out_uop_ldst_is_rs1 : _slots_4_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_15
         ? _slots_6_io_out_uop_ldst
         : _GEN_14 ? _slots_5_io_out_uop_ldst : _slots_4_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_15
         ? _slots_6_io_out_uop_lrs1
         : _GEN_14 ? _slots_5_io_out_uop_lrs1 : _slots_4_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_15
         ? _slots_6_io_out_uop_lrs2
         : _GEN_14 ? _slots_5_io_out_uop_lrs2 : _slots_4_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_15
         ? _slots_6_io_out_uop_lrs3
         : _GEN_14 ? _slots_5_io_out_uop_lrs3 : _slots_4_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_15
         ? _slots_6_io_out_uop_ldst_val
         : _GEN_14 ? _slots_5_io_out_uop_ldst_val : _slots_4_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_15
         ? _slots_6_io_out_uop_dst_rtype
         : _GEN_14 ? _slots_5_io_out_uop_dst_rtype : _slots_4_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_15
         ? _slots_6_io_out_uop_lrs1_rtype
         : _GEN_14 ? _slots_5_io_out_uop_lrs1_rtype : _slots_4_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_15
         ? _slots_6_io_out_uop_lrs2_rtype
         : _GEN_14 ? _slots_5_io_out_uop_lrs2_rtype : _slots_4_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_15
         ? _slots_6_io_out_uop_frs3_en
         : _GEN_14 ? _slots_5_io_out_uop_frs3_en : _slots_4_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_15
         ? _slots_6_io_out_uop_fp_val
         : _GEN_14 ? _slots_5_io_out_uop_fp_val : _slots_4_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_15
         ? _slots_6_io_out_uop_fp_single
         : _GEN_14 ? _slots_5_io_out_uop_fp_single : _slots_4_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_15
         ? _slots_6_io_out_uop_xcpt_pf_if
         : _GEN_14 ? _slots_5_io_out_uop_xcpt_pf_if : _slots_4_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_15
         ? _slots_6_io_out_uop_xcpt_ae_if
         : _GEN_14 ? _slots_5_io_out_uop_xcpt_ae_if : _slots_4_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_15
         ? _slots_6_io_out_uop_xcpt_ma_if
         : _GEN_14 ? _slots_5_io_out_uop_xcpt_ma_if : _slots_4_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_15
         ? _slots_6_io_out_uop_bp_debug_if
         : _GEN_14 ? _slots_5_io_out_uop_bp_debug_if : _slots_4_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_15
         ? _slots_6_io_out_uop_bp_xcpt_if
         : _GEN_14 ? _slots_5_io_out_uop_bp_xcpt_if : _slots_4_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_15
         ? _slots_6_io_out_uop_debug_fsrc
         : _GEN_14 ? _slots_5_io_out_uop_debug_fsrc : _slots_4_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_15
         ? _slots_6_io_out_uop_debug_tsrc
         : _GEN_14 ? _slots_5_io_out_uop_debug_tsrc : _slots_4_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_3_io_valid),
    .io_will_be_valid               (_slots_3_io_will_be_valid),
    .io_request                     (_slots_3_io_request),
    .io_out_uop_uopc                (_slots_3_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_3_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_3_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_3_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_3_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_3_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_3_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_3_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_3_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_3_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_3_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_3_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_3_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_3_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_3_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_3_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_3_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_3_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_3_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_3_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_3_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_3_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_3_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_3_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_3_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_3_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_3_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_3_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_3_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_3_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_3_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_3_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_3_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_3_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_3_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_3_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_3_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_3_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_3_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_3_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_3_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_3_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_3_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_3_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_3_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_3_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_3_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_3_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_3_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_3_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_3_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_3_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_3_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_3_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_3_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_3_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_3_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_3_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_3_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_3_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_3_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_3_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_3_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_3_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_3_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_3_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_3_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_3_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_3_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_3_io_uop_uopc),
    .io_uop_inst                    (_slots_3_io_uop_inst),
    .io_uop_debug_inst              (_slots_3_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_3_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_3_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_3_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_3_io_uop_fu_code),
    .io_uop_iw_state                (_slots_3_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_3_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_3_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_3_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_3_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_3_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_3_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_3_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_3_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_3_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_3_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_3_io_uop_pc_lob),
    .io_uop_taken                   (_slots_3_io_uop_taken),
    .io_uop_imm_packed              (_slots_3_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_3_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_3_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_3_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_3_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_3_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_3_io_uop_pdst),
    .io_uop_prs1                    (_slots_3_io_uop_prs1),
    .io_uop_prs2                    (_slots_3_io_uop_prs2),
    .io_uop_prs3                    (_slots_3_io_uop_prs3),
    .io_uop_ppred                   (_slots_3_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_3_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_3_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_3_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_3_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_3_io_uop_stale_pdst),
    .io_uop_exception               (_slots_3_io_uop_exception),
    .io_uop_exc_cause               (_slots_3_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_3_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_3_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_3_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_3_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_3_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_3_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_3_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_3_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_3_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_3_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_3_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_3_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_3_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_3_io_uop_ldst),
    .io_uop_lrs1                    (_slots_3_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_3_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_3_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_3_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_3_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_3_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_3_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_3_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_3_io_uop_fp_val),
    .io_uop_fp_single               (_slots_3_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_3_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_3_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_3_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_3_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_3_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_3_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_3_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_4 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_4_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_3),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_4_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_17
         ? _slots_7_io_out_uop_uopc
         : _GEN_16 ? _slots_6_io_out_uop_uopc : _slots_5_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_17
         ? _slots_7_io_out_uop_inst
         : _GEN_16 ? _slots_6_io_out_uop_inst : _slots_5_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_17
         ? _slots_7_io_out_uop_debug_inst
         : _GEN_16 ? _slots_6_io_out_uop_debug_inst : _slots_5_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_17
         ? _slots_7_io_out_uop_is_rvc
         : _GEN_16 ? _slots_6_io_out_uop_is_rvc : _slots_5_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_17
         ? _slots_7_io_out_uop_debug_pc
         : _GEN_16 ? _slots_6_io_out_uop_debug_pc : _slots_5_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_17
         ? _slots_7_io_out_uop_iq_type
         : _GEN_16 ? _slots_6_io_out_uop_iq_type : _slots_5_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_17
         ? _slots_7_io_out_uop_fu_code
         : _GEN_16 ? _slots_6_io_out_uop_fu_code : _slots_5_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_17
         ? _slots_7_io_out_uop_iw_state
         : _GEN_16 ? _slots_6_io_out_uop_iw_state : _slots_5_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_17
         ? _slots_7_io_out_uop_iw_p1_poisoned
         : _GEN_16
             ? _slots_6_io_out_uop_iw_p1_poisoned
             : _slots_5_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_17
         ? _slots_7_io_out_uop_iw_p2_poisoned
         : _GEN_16
             ? _slots_6_io_out_uop_iw_p2_poisoned
             : _slots_5_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_17
         ? _slots_7_io_out_uop_is_br
         : _GEN_16 ? _slots_6_io_out_uop_is_br : _slots_5_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_17
         ? _slots_7_io_out_uop_is_jalr
         : _GEN_16 ? _slots_6_io_out_uop_is_jalr : _slots_5_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_17
         ? _slots_7_io_out_uop_is_jal
         : _GEN_16 ? _slots_6_io_out_uop_is_jal : _slots_5_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_17
         ? _slots_7_io_out_uop_is_sfb
         : _GEN_16 ? _slots_6_io_out_uop_is_sfb : _slots_5_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_17
         ? _slots_7_io_out_uop_br_mask
         : _GEN_16 ? _slots_6_io_out_uop_br_mask : _slots_5_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_17
         ? _slots_7_io_out_uop_br_tag
         : _GEN_16 ? _slots_6_io_out_uop_br_tag : _slots_5_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_17
         ? _slots_7_io_out_uop_ftq_idx
         : _GEN_16 ? _slots_6_io_out_uop_ftq_idx : _slots_5_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_17
         ? _slots_7_io_out_uop_edge_inst
         : _GEN_16 ? _slots_6_io_out_uop_edge_inst : _slots_5_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_17
         ? _slots_7_io_out_uop_pc_lob
         : _GEN_16 ? _slots_6_io_out_uop_pc_lob : _slots_5_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_17
         ? _slots_7_io_out_uop_taken
         : _GEN_16 ? _slots_6_io_out_uop_taken : _slots_5_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_17
         ? _slots_7_io_out_uop_imm_packed
         : _GEN_16 ? _slots_6_io_out_uop_imm_packed : _slots_5_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_17
         ? _slots_7_io_out_uop_csr_addr
         : _GEN_16 ? _slots_6_io_out_uop_csr_addr : _slots_5_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_17
         ? _slots_7_io_out_uop_rob_idx
         : _GEN_16 ? _slots_6_io_out_uop_rob_idx : _slots_5_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_17
         ? _slots_7_io_out_uop_ldq_idx
         : _GEN_16 ? _slots_6_io_out_uop_ldq_idx : _slots_5_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_17
         ? _slots_7_io_out_uop_stq_idx
         : _GEN_16 ? _slots_6_io_out_uop_stq_idx : _slots_5_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_17
         ? _slots_7_io_out_uop_rxq_idx
         : _GEN_16 ? _slots_6_io_out_uop_rxq_idx : _slots_5_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_17
         ? _slots_7_io_out_uop_pdst
         : _GEN_16 ? _slots_6_io_out_uop_pdst : _slots_5_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_17
         ? _slots_7_io_out_uop_prs1
         : _GEN_16 ? _slots_6_io_out_uop_prs1 : _slots_5_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_17
         ? _slots_7_io_out_uop_prs2
         : _GEN_16 ? _slots_6_io_out_uop_prs2 : _slots_5_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_17
         ? _slots_7_io_out_uop_prs3
         : _GEN_16 ? _slots_6_io_out_uop_prs3 : _slots_5_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_17
         ? _slots_7_io_out_uop_ppred
         : _GEN_16 ? _slots_6_io_out_uop_ppred : _slots_5_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_17
         ? _slots_7_io_out_uop_prs1_busy
         : _GEN_16 ? _slots_6_io_out_uop_prs1_busy : _slots_5_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_17
         ? _slots_7_io_out_uop_prs2_busy
         : _GEN_16 ? _slots_6_io_out_uop_prs2_busy : _slots_5_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_17
         ? _slots_7_io_out_uop_prs3_busy
         : _GEN_16 ? _slots_6_io_out_uop_prs3_busy : _slots_5_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_17
         ? _slots_7_io_out_uop_ppred_busy
         : _GEN_16 ? _slots_6_io_out_uop_ppred_busy : _slots_5_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_17
         ? _slots_7_io_out_uop_stale_pdst
         : _GEN_16 ? _slots_6_io_out_uop_stale_pdst : _slots_5_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_17
         ? _slots_7_io_out_uop_exception
         : _GEN_16 ? _slots_6_io_out_uop_exception : _slots_5_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_17
         ? _slots_7_io_out_uop_exc_cause
         : _GEN_16 ? _slots_6_io_out_uop_exc_cause : _slots_5_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_17
         ? _slots_7_io_out_uop_bypassable
         : _GEN_16 ? _slots_6_io_out_uop_bypassable : _slots_5_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_17
         ? _slots_7_io_out_uop_mem_cmd
         : _GEN_16 ? _slots_6_io_out_uop_mem_cmd : _slots_5_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_17
         ? _slots_7_io_out_uop_mem_size
         : _GEN_16 ? _slots_6_io_out_uop_mem_size : _slots_5_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_17
         ? _slots_7_io_out_uop_mem_signed
         : _GEN_16 ? _slots_6_io_out_uop_mem_signed : _slots_5_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_17
         ? _slots_7_io_out_uop_is_fence
         : _GEN_16 ? _slots_6_io_out_uop_is_fence : _slots_5_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_17
         ? _slots_7_io_out_uop_is_fencei
         : _GEN_16 ? _slots_6_io_out_uop_is_fencei : _slots_5_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_17
         ? _slots_7_io_out_uop_is_amo
         : _GEN_16 ? _slots_6_io_out_uop_is_amo : _slots_5_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_17
         ? _slots_7_io_out_uop_uses_ldq
         : _GEN_16 ? _slots_6_io_out_uop_uses_ldq : _slots_5_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_17
         ? _slots_7_io_out_uop_uses_stq
         : _GEN_16 ? _slots_6_io_out_uop_uses_stq : _slots_5_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_17
         ? _slots_7_io_out_uop_is_sys_pc2epc
         : _GEN_16
             ? _slots_6_io_out_uop_is_sys_pc2epc
             : _slots_5_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_17
         ? _slots_7_io_out_uop_is_unique
         : _GEN_16 ? _slots_6_io_out_uop_is_unique : _slots_5_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_17
         ? _slots_7_io_out_uop_flush_on_commit
         : _GEN_16
             ? _slots_6_io_out_uop_flush_on_commit
             : _slots_5_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_17
         ? _slots_7_io_out_uop_ldst_is_rs1
         : _GEN_16 ? _slots_6_io_out_uop_ldst_is_rs1 : _slots_5_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_17
         ? _slots_7_io_out_uop_ldst
         : _GEN_16 ? _slots_6_io_out_uop_ldst : _slots_5_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_17
         ? _slots_7_io_out_uop_lrs1
         : _GEN_16 ? _slots_6_io_out_uop_lrs1 : _slots_5_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_17
         ? _slots_7_io_out_uop_lrs2
         : _GEN_16 ? _slots_6_io_out_uop_lrs2 : _slots_5_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_17
         ? _slots_7_io_out_uop_lrs3
         : _GEN_16 ? _slots_6_io_out_uop_lrs3 : _slots_5_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_17
         ? _slots_7_io_out_uop_ldst_val
         : _GEN_16 ? _slots_6_io_out_uop_ldst_val : _slots_5_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_17
         ? _slots_7_io_out_uop_dst_rtype
         : _GEN_16 ? _slots_6_io_out_uop_dst_rtype : _slots_5_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_17
         ? _slots_7_io_out_uop_lrs1_rtype
         : _GEN_16 ? _slots_6_io_out_uop_lrs1_rtype : _slots_5_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_17
         ? _slots_7_io_out_uop_lrs2_rtype
         : _GEN_16 ? _slots_6_io_out_uop_lrs2_rtype : _slots_5_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_17
         ? _slots_7_io_out_uop_frs3_en
         : _GEN_16 ? _slots_6_io_out_uop_frs3_en : _slots_5_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_17
         ? _slots_7_io_out_uop_fp_val
         : _GEN_16 ? _slots_6_io_out_uop_fp_val : _slots_5_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_17
         ? _slots_7_io_out_uop_fp_single
         : _GEN_16 ? _slots_6_io_out_uop_fp_single : _slots_5_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_17
         ? _slots_7_io_out_uop_xcpt_pf_if
         : _GEN_16 ? _slots_6_io_out_uop_xcpt_pf_if : _slots_5_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_17
         ? _slots_7_io_out_uop_xcpt_ae_if
         : _GEN_16 ? _slots_6_io_out_uop_xcpt_ae_if : _slots_5_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_17
         ? _slots_7_io_out_uop_xcpt_ma_if
         : _GEN_16 ? _slots_6_io_out_uop_xcpt_ma_if : _slots_5_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_17
         ? _slots_7_io_out_uop_bp_debug_if
         : _GEN_16 ? _slots_6_io_out_uop_bp_debug_if : _slots_5_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_17
         ? _slots_7_io_out_uop_bp_xcpt_if
         : _GEN_16 ? _slots_6_io_out_uop_bp_xcpt_if : _slots_5_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_17
         ? _slots_7_io_out_uop_debug_fsrc
         : _GEN_16 ? _slots_6_io_out_uop_debug_fsrc : _slots_5_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_17
         ? _slots_7_io_out_uop_debug_tsrc
         : _GEN_16 ? _slots_6_io_out_uop_debug_tsrc : _slots_5_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_4_io_valid),
    .io_will_be_valid               (_slots_4_io_will_be_valid),
    .io_request                     (_slots_4_io_request),
    .io_out_uop_uopc                (_slots_4_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_4_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_4_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_4_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_4_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_4_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_4_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_4_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_4_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_4_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_4_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_4_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_4_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_4_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_4_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_4_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_4_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_4_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_4_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_4_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_4_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_4_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_4_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_4_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_4_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_4_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_4_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_4_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_4_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_4_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_4_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_4_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_4_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_4_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_4_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_4_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_4_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_4_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_4_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_4_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_4_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_4_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_4_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_4_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_4_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_4_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_4_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_4_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_4_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_4_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_4_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_4_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_4_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_4_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_4_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_4_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_4_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_4_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_4_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_4_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_4_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_4_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_4_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_4_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_4_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_4_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_4_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_4_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_4_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_4_io_uop_uopc),
    .io_uop_inst                    (_slots_4_io_uop_inst),
    .io_uop_debug_inst              (_slots_4_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_4_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_4_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_4_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_4_io_uop_fu_code),
    .io_uop_iw_state                (_slots_4_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_4_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_4_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_4_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_4_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_4_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_4_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_4_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_4_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_4_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_4_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_4_io_uop_pc_lob),
    .io_uop_taken                   (_slots_4_io_uop_taken),
    .io_uop_imm_packed              (_slots_4_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_4_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_4_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_4_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_4_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_4_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_4_io_uop_pdst),
    .io_uop_prs1                    (_slots_4_io_uop_prs1),
    .io_uop_prs2                    (_slots_4_io_uop_prs2),
    .io_uop_prs3                    (_slots_4_io_uop_prs3),
    .io_uop_ppred                   (_slots_4_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_4_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_4_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_4_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_4_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_4_io_uop_stale_pdst),
    .io_uop_exception               (_slots_4_io_uop_exception),
    .io_uop_exc_cause               (_slots_4_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_4_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_4_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_4_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_4_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_4_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_4_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_4_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_4_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_4_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_4_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_4_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_4_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_4_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_4_io_uop_ldst),
    .io_uop_lrs1                    (_slots_4_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_4_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_4_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_4_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_4_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_4_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_4_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_4_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_4_io_uop_fp_val),
    .io_uop_fp_single               (_slots_4_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_4_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_4_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_4_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_4_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_4_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_4_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_4_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_5 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_5_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_4),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_5_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_19
         ? _slots_8_io_out_uop_uopc
         : _GEN_18 ? _slots_7_io_out_uop_uopc : _slots_6_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_19
         ? _slots_8_io_out_uop_inst
         : _GEN_18 ? _slots_7_io_out_uop_inst : _slots_6_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_19
         ? _slots_8_io_out_uop_debug_inst
         : _GEN_18 ? _slots_7_io_out_uop_debug_inst : _slots_6_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_19
         ? _slots_8_io_out_uop_is_rvc
         : _GEN_18 ? _slots_7_io_out_uop_is_rvc : _slots_6_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_19
         ? _slots_8_io_out_uop_debug_pc
         : _GEN_18 ? _slots_7_io_out_uop_debug_pc : _slots_6_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_19
         ? _slots_8_io_out_uop_iq_type
         : _GEN_18 ? _slots_7_io_out_uop_iq_type : _slots_6_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_19
         ? _slots_8_io_out_uop_fu_code
         : _GEN_18 ? _slots_7_io_out_uop_fu_code : _slots_6_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_19
         ? _slots_8_io_out_uop_iw_state
         : _GEN_18 ? _slots_7_io_out_uop_iw_state : _slots_6_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_19
         ? _slots_8_io_out_uop_iw_p1_poisoned
         : _GEN_18
             ? _slots_7_io_out_uop_iw_p1_poisoned
             : _slots_6_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_19
         ? _slots_8_io_out_uop_iw_p2_poisoned
         : _GEN_18
             ? _slots_7_io_out_uop_iw_p2_poisoned
             : _slots_6_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_19
         ? _slots_8_io_out_uop_is_br
         : _GEN_18 ? _slots_7_io_out_uop_is_br : _slots_6_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_19
         ? _slots_8_io_out_uop_is_jalr
         : _GEN_18 ? _slots_7_io_out_uop_is_jalr : _slots_6_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_19
         ? _slots_8_io_out_uop_is_jal
         : _GEN_18 ? _slots_7_io_out_uop_is_jal : _slots_6_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_19
         ? _slots_8_io_out_uop_is_sfb
         : _GEN_18 ? _slots_7_io_out_uop_is_sfb : _slots_6_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_19
         ? _slots_8_io_out_uop_br_mask
         : _GEN_18 ? _slots_7_io_out_uop_br_mask : _slots_6_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_19
         ? _slots_8_io_out_uop_br_tag
         : _GEN_18 ? _slots_7_io_out_uop_br_tag : _slots_6_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_19
         ? _slots_8_io_out_uop_ftq_idx
         : _GEN_18 ? _slots_7_io_out_uop_ftq_idx : _slots_6_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_19
         ? _slots_8_io_out_uop_edge_inst
         : _GEN_18 ? _slots_7_io_out_uop_edge_inst : _slots_6_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_19
         ? _slots_8_io_out_uop_pc_lob
         : _GEN_18 ? _slots_7_io_out_uop_pc_lob : _slots_6_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_19
         ? _slots_8_io_out_uop_taken
         : _GEN_18 ? _slots_7_io_out_uop_taken : _slots_6_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_19
         ? _slots_8_io_out_uop_imm_packed
         : _GEN_18 ? _slots_7_io_out_uop_imm_packed : _slots_6_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_19
         ? _slots_8_io_out_uop_csr_addr
         : _GEN_18 ? _slots_7_io_out_uop_csr_addr : _slots_6_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_19
         ? _slots_8_io_out_uop_rob_idx
         : _GEN_18 ? _slots_7_io_out_uop_rob_idx : _slots_6_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_19
         ? _slots_8_io_out_uop_ldq_idx
         : _GEN_18 ? _slots_7_io_out_uop_ldq_idx : _slots_6_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_19
         ? _slots_8_io_out_uop_stq_idx
         : _GEN_18 ? _slots_7_io_out_uop_stq_idx : _slots_6_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_19
         ? _slots_8_io_out_uop_rxq_idx
         : _GEN_18 ? _slots_7_io_out_uop_rxq_idx : _slots_6_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_19
         ? _slots_8_io_out_uop_pdst
         : _GEN_18 ? _slots_7_io_out_uop_pdst : _slots_6_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_19
         ? _slots_8_io_out_uop_prs1
         : _GEN_18 ? _slots_7_io_out_uop_prs1 : _slots_6_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_19
         ? _slots_8_io_out_uop_prs2
         : _GEN_18 ? _slots_7_io_out_uop_prs2 : _slots_6_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_19
         ? _slots_8_io_out_uop_prs3
         : _GEN_18 ? _slots_7_io_out_uop_prs3 : _slots_6_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_19
         ? _slots_8_io_out_uop_ppred
         : _GEN_18 ? _slots_7_io_out_uop_ppred : _slots_6_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_19
         ? _slots_8_io_out_uop_prs1_busy
         : _GEN_18 ? _slots_7_io_out_uop_prs1_busy : _slots_6_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_19
         ? _slots_8_io_out_uop_prs2_busy
         : _GEN_18 ? _slots_7_io_out_uop_prs2_busy : _slots_6_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_19
         ? _slots_8_io_out_uop_prs3_busy
         : _GEN_18 ? _slots_7_io_out_uop_prs3_busy : _slots_6_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_19
         ? _slots_8_io_out_uop_ppred_busy
         : _GEN_18 ? _slots_7_io_out_uop_ppred_busy : _slots_6_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_19
         ? _slots_8_io_out_uop_stale_pdst
         : _GEN_18 ? _slots_7_io_out_uop_stale_pdst : _slots_6_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_19
         ? _slots_8_io_out_uop_exception
         : _GEN_18 ? _slots_7_io_out_uop_exception : _slots_6_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_19
         ? _slots_8_io_out_uop_exc_cause
         : _GEN_18 ? _slots_7_io_out_uop_exc_cause : _slots_6_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_19
         ? _slots_8_io_out_uop_bypassable
         : _GEN_18 ? _slots_7_io_out_uop_bypassable : _slots_6_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_19
         ? _slots_8_io_out_uop_mem_cmd
         : _GEN_18 ? _slots_7_io_out_uop_mem_cmd : _slots_6_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_19
         ? _slots_8_io_out_uop_mem_size
         : _GEN_18 ? _slots_7_io_out_uop_mem_size : _slots_6_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_19
         ? _slots_8_io_out_uop_mem_signed
         : _GEN_18 ? _slots_7_io_out_uop_mem_signed : _slots_6_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_19
         ? _slots_8_io_out_uop_is_fence
         : _GEN_18 ? _slots_7_io_out_uop_is_fence : _slots_6_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_19
         ? _slots_8_io_out_uop_is_fencei
         : _GEN_18 ? _slots_7_io_out_uop_is_fencei : _slots_6_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_19
         ? _slots_8_io_out_uop_is_amo
         : _GEN_18 ? _slots_7_io_out_uop_is_amo : _slots_6_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_19
         ? _slots_8_io_out_uop_uses_ldq
         : _GEN_18 ? _slots_7_io_out_uop_uses_ldq : _slots_6_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_19
         ? _slots_8_io_out_uop_uses_stq
         : _GEN_18 ? _slots_7_io_out_uop_uses_stq : _slots_6_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_19
         ? _slots_8_io_out_uop_is_sys_pc2epc
         : _GEN_18
             ? _slots_7_io_out_uop_is_sys_pc2epc
             : _slots_6_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_19
         ? _slots_8_io_out_uop_is_unique
         : _GEN_18 ? _slots_7_io_out_uop_is_unique : _slots_6_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_19
         ? _slots_8_io_out_uop_flush_on_commit
         : _GEN_18
             ? _slots_7_io_out_uop_flush_on_commit
             : _slots_6_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_19
         ? _slots_8_io_out_uop_ldst_is_rs1
         : _GEN_18 ? _slots_7_io_out_uop_ldst_is_rs1 : _slots_6_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_19
         ? _slots_8_io_out_uop_ldst
         : _GEN_18 ? _slots_7_io_out_uop_ldst : _slots_6_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_19
         ? _slots_8_io_out_uop_lrs1
         : _GEN_18 ? _slots_7_io_out_uop_lrs1 : _slots_6_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_19
         ? _slots_8_io_out_uop_lrs2
         : _GEN_18 ? _slots_7_io_out_uop_lrs2 : _slots_6_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_19
         ? _slots_8_io_out_uop_lrs3
         : _GEN_18 ? _slots_7_io_out_uop_lrs3 : _slots_6_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_19
         ? _slots_8_io_out_uop_ldst_val
         : _GEN_18 ? _slots_7_io_out_uop_ldst_val : _slots_6_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_19
         ? _slots_8_io_out_uop_dst_rtype
         : _GEN_18 ? _slots_7_io_out_uop_dst_rtype : _slots_6_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_19
         ? _slots_8_io_out_uop_lrs1_rtype
         : _GEN_18 ? _slots_7_io_out_uop_lrs1_rtype : _slots_6_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_19
         ? _slots_8_io_out_uop_lrs2_rtype
         : _GEN_18 ? _slots_7_io_out_uop_lrs2_rtype : _slots_6_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_19
         ? _slots_8_io_out_uop_frs3_en
         : _GEN_18 ? _slots_7_io_out_uop_frs3_en : _slots_6_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_19
         ? _slots_8_io_out_uop_fp_val
         : _GEN_18 ? _slots_7_io_out_uop_fp_val : _slots_6_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_19
         ? _slots_8_io_out_uop_fp_single
         : _GEN_18 ? _slots_7_io_out_uop_fp_single : _slots_6_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_19
         ? _slots_8_io_out_uop_xcpt_pf_if
         : _GEN_18 ? _slots_7_io_out_uop_xcpt_pf_if : _slots_6_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_19
         ? _slots_8_io_out_uop_xcpt_ae_if
         : _GEN_18 ? _slots_7_io_out_uop_xcpt_ae_if : _slots_6_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_19
         ? _slots_8_io_out_uop_xcpt_ma_if
         : _GEN_18 ? _slots_7_io_out_uop_xcpt_ma_if : _slots_6_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_19
         ? _slots_8_io_out_uop_bp_debug_if
         : _GEN_18 ? _slots_7_io_out_uop_bp_debug_if : _slots_6_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_19
         ? _slots_8_io_out_uop_bp_xcpt_if
         : _GEN_18 ? _slots_7_io_out_uop_bp_xcpt_if : _slots_6_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_19
         ? _slots_8_io_out_uop_debug_fsrc
         : _GEN_18 ? _slots_7_io_out_uop_debug_fsrc : _slots_6_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_19
         ? _slots_8_io_out_uop_debug_tsrc
         : _GEN_18 ? _slots_7_io_out_uop_debug_tsrc : _slots_6_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_5_io_valid),
    .io_will_be_valid               (_slots_5_io_will_be_valid),
    .io_request                     (_slots_5_io_request),
    .io_out_uop_uopc                (_slots_5_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_5_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_5_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_5_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_5_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_5_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_5_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_5_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_5_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_5_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_5_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_5_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_5_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_5_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_5_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_5_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_5_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_5_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_5_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_5_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_5_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_5_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_5_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_5_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_5_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_5_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_5_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_5_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_5_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_5_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_5_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_5_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_5_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_5_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_5_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_5_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_5_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_5_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_5_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_5_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_5_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_5_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_5_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_5_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_5_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_5_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_5_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_5_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_5_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_5_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_5_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_5_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_5_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_5_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_5_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_5_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_5_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_5_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_5_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_5_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_5_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_5_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_5_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_5_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_5_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_5_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_5_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_5_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_5_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_5_io_uop_uopc),
    .io_uop_inst                    (_slots_5_io_uop_inst),
    .io_uop_debug_inst              (_slots_5_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_5_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_5_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_5_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_5_io_uop_fu_code),
    .io_uop_iw_state                (_slots_5_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_5_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_5_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_5_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_5_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_5_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_5_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_5_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_5_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_5_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_5_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_5_io_uop_pc_lob),
    .io_uop_taken                   (_slots_5_io_uop_taken),
    .io_uop_imm_packed              (_slots_5_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_5_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_5_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_5_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_5_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_5_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_5_io_uop_pdst),
    .io_uop_prs1                    (_slots_5_io_uop_prs1),
    .io_uop_prs2                    (_slots_5_io_uop_prs2),
    .io_uop_prs3                    (_slots_5_io_uop_prs3),
    .io_uop_ppred                   (_slots_5_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_5_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_5_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_5_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_5_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_5_io_uop_stale_pdst),
    .io_uop_exception               (_slots_5_io_uop_exception),
    .io_uop_exc_cause               (_slots_5_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_5_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_5_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_5_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_5_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_5_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_5_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_5_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_5_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_5_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_5_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_5_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_5_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_5_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_5_io_uop_ldst),
    .io_uop_lrs1                    (_slots_5_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_5_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_5_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_5_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_5_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_5_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_5_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_5_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_5_io_uop_fp_val),
    .io_uop_fp_single               (_slots_5_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_5_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_5_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_5_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_5_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_5_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_5_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_5_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_6 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_6_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_5),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_6_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_21
         ? _slots_9_io_out_uop_uopc
         : _GEN_20 ? _slots_8_io_out_uop_uopc : _slots_7_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_21
         ? _slots_9_io_out_uop_inst
         : _GEN_20 ? _slots_8_io_out_uop_inst : _slots_7_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_21
         ? _slots_9_io_out_uop_debug_inst
         : _GEN_20 ? _slots_8_io_out_uop_debug_inst : _slots_7_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_21
         ? _slots_9_io_out_uop_is_rvc
         : _GEN_20 ? _slots_8_io_out_uop_is_rvc : _slots_7_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_21
         ? _slots_9_io_out_uop_debug_pc
         : _GEN_20 ? _slots_8_io_out_uop_debug_pc : _slots_7_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_21
         ? _slots_9_io_out_uop_iq_type
         : _GEN_20 ? _slots_8_io_out_uop_iq_type : _slots_7_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_21
         ? _slots_9_io_out_uop_fu_code
         : _GEN_20 ? _slots_8_io_out_uop_fu_code : _slots_7_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_21
         ? _slots_9_io_out_uop_iw_state
         : _GEN_20 ? _slots_8_io_out_uop_iw_state : _slots_7_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_21
         ? _slots_9_io_out_uop_iw_p1_poisoned
         : _GEN_20
             ? _slots_8_io_out_uop_iw_p1_poisoned
             : _slots_7_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_21
         ? _slots_9_io_out_uop_iw_p2_poisoned
         : _GEN_20
             ? _slots_8_io_out_uop_iw_p2_poisoned
             : _slots_7_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_21
         ? _slots_9_io_out_uop_is_br
         : _GEN_20 ? _slots_8_io_out_uop_is_br : _slots_7_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_21
         ? _slots_9_io_out_uop_is_jalr
         : _GEN_20 ? _slots_8_io_out_uop_is_jalr : _slots_7_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_21
         ? _slots_9_io_out_uop_is_jal
         : _GEN_20 ? _slots_8_io_out_uop_is_jal : _slots_7_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_21
         ? _slots_9_io_out_uop_is_sfb
         : _GEN_20 ? _slots_8_io_out_uop_is_sfb : _slots_7_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_21
         ? _slots_9_io_out_uop_br_mask
         : _GEN_20 ? _slots_8_io_out_uop_br_mask : _slots_7_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_21
         ? _slots_9_io_out_uop_br_tag
         : _GEN_20 ? _slots_8_io_out_uop_br_tag : _slots_7_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_21
         ? _slots_9_io_out_uop_ftq_idx
         : _GEN_20 ? _slots_8_io_out_uop_ftq_idx : _slots_7_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_21
         ? _slots_9_io_out_uop_edge_inst
         : _GEN_20 ? _slots_8_io_out_uop_edge_inst : _slots_7_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_21
         ? _slots_9_io_out_uop_pc_lob
         : _GEN_20 ? _slots_8_io_out_uop_pc_lob : _slots_7_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_21
         ? _slots_9_io_out_uop_taken
         : _GEN_20 ? _slots_8_io_out_uop_taken : _slots_7_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_21
         ? _slots_9_io_out_uop_imm_packed
         : _GEN_20 ? _slots_8_io_out_uop_imm_packed : _slots_7_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_21
         ? _slots_9_io_out_uop_csr_addr
         : _GEN_20 ? _slots_8_io_out_uop_csr_addr : _slots_7_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_21
         ? _slots_9_io_out_uop_rob_idx
         : _GEN_20 ? _slots_8_io_out_uop_rob_idx : _slots_7_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_21
         ? _slots_9_io_out_uop_ldq_idx
         : _GEN_20 ? _slots_8_io_out_uop_ldq_idx : _slots_7_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_21
         ? _slots_9_io_out_uop_stq_idx
         : _GEN_20 ? _slots_8_io_out_uop_stq_idx : _slots_7_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_21
         ? _slots_9_io_out_uop_rxq_idx
         : _GEN_20 ? _slots_8_io_out_uop_rxq_idx : _slots_7_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_21
         ? _slots_9_io_out_uop_pdst
         : _GEN_20 ? _slots_8_io_out_uop_pdst : _slots_7_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_21
         ? _slots_9_io_out_uop_prs1
         : _GEN_20 ? _slots_8_io_out_uop_prs1 : _slots_7_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_21
         ? _slots_9_io_out_uop_prs2
         : _GEN_20 ? _slots_8_io_out_uop_prs2 : _slots_7_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_21
         ? _slots_9_io_out_uop_prs3
         : _GEN_20 ? _slots_8_io_out_uop_prs3 : _slots_7_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_21
         ? _slots_9_io_out_uop_ppred
         : _GEN_20 ? _slots_8_io_out_uop_ppred : _slots_7_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_21
         ? _slots_9_io_out_uop_prs1_busy
         : _GEN_20 ? _slots_8_io_out_uop_prs1_busy : _slots_7_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_21
         ? _slots_9_io_out_uop_prs2_busy
         : _GEN_20 ? _slots_8_io_out_uop_prs2_busy : _slots_7_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_21
         ? _slots_9_io_out_uop_prs3_busy
         : _GEN_20 ? _slots_8_io_out_uop_prs3_busy : _slots_7_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_21
         ? _slots_9_io_out_uop_ppred_busy
         : _GEN_20 ? _slots_8_io_out_uop_ppred_busy : _slots_7_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_21
         ? _slots_9_io_out_uop_stale_pdst
         : _GEN_20 ? _slots_8_io_out_uop_stale_pdst : _slots_7_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_21
         ? _slots_9_io_out_uop_exception
         : _GEN_20 ? _slots_8_io_out_uop_exception : _slots_7_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_21
         ? _slots_9_io_out_uop_exc_cause
         : _GEN_20 ? _slots_8_io_out_uop_exc_cause : _slots_7_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_21
         ? _slots_9_io_out_uop_bypassable
         : _GEN_20 ? _slots_8_io_out_uop_bypassable : _slots_7_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_21
         ? _slots_9_io_out_uop_mem_cmd
         : _GEN_20 ? _slots_8_io_out_uop_mem_cmd : _slots_7_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_21
         ? _slots_9_io_out_uop_mem_size
         : _GEN_20 ? _slots_8_io_out_uop_mem_size : _slots_7_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_21
         ? _slots_9_io_out_uop_mem_signed
         : _GEN_20 ? _slots_8_io_out_uop_mem_signed : _slots_7_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_21
         ? _slots_9_io_out_uop_is_fence
         : _GEN_20 ? _slots_8_io_out_uop_is_fence : _slots_7_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_21
         ? _slots_9_io_out_uop_is_fencei
         : _GEN_20 ? _slots_8_io_out_uop_is_fencei : _slots_7_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_21
         ? _slots_9_io_out_uop_is_amo
         : _GEN_20 ? _slots_8_io_out_uop_is_amo : _slots_7_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_21
         ? _slots_9_io_out_uop_uses_ldq
         : _GEN_20 ? _slots_8_io_out_uop_uses_ldq : _slots_7_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_21
         ? _slots_9_io_out_uop_uses_stq
         : _GEN_20 ? _slots_8_io_out_uop_uses_stq : _slots_7_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_21
         ? _slots_9_io_out_uop_is_sys_pc2epc
         : _GEN_20
             ? _slots_8_io_out_uop_is_sys_pc2epc
             : _slots_7_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_21
         ? _slots_9_io_out_uop_is_unique
         : _GEN_20 ? _slots_8_io_out_uop_is_unique : _slots_7_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_21
         ? _slots_9_io_out_uop_flush_on_commit
         : _GEN_20
             ? _slots_8_io_out_uop_flush_on_commit
             : _slots_7_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_21
         ? _slots_9_io_out_uop_ldst_is_rs1
         : _GEN_20 ? _slots_8_io_out_uop_ldst_is_rs1 : _slots_7_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_21
         ? _slots_9_io_out_uop_ldst
         : _GEN_20 ? _slots_8_io_out_uop_ldst : _slots_7_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_21
         ? _slots_9_io_out_uop_lrs1
         : _GEN_20 ? _slots_8_io_out_uop_lrs1 : _slots_7_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_21
         ? _slots_9_io_out_uop_lrs2
         : _GEN_20 ? _slots_8_io_out_uop_lrs2 : _slots_7_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_21
         ? _slots_9_io_out_uop_lrs3
         : _GEN_20 ? _slots_8_io_out_uop_lrs3 : _slots_7_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_21
         ? _slots_9_io_out_uop_ldst_val
         : _GEN_20 ? _slots_8_io_out_uop_ldst_val : _slots_7_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_21
         ? _slots_9_io_out_uop_dst_rtype
         : _GEN_20 ? _slots_8_io_out_uop_dst_rtype : _slots_7_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_21
         ? _slots_9_io_out_uop_lrs1_rtype
         : _GEN_20 ? _slots_8_io_out_uop_lrs1_rtype : _slots_7_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_21
         ? _slots_9_io_out_uop_lrs2_rtype
         : _GEN_20 ? _slots_8_io_out_uop_lrs2_rtype : _slots_7_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_21
         ? _slots_9_io_out_uop_frs3_en
         : _GEN_20 ? _slots_8_io_out_uop_frs3_en : _slots_7_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_21
         ? _slots_9_io_out_uop_fp_val
         : _GEN_20 ? _slots_8_io_out_uop_fp_val : _slots_7_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_21
         ? _slots_9_io_out_uop_fp_single
         : _GEN_20 ? _slots_8_io_out_uop_fp_single : _slots_7_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_21
         ? _slots_9_io_out_uop_xcpt_pf_if
         : _GEN_20 ? _slots_8_io_out_uop_xcpt_pf_if : _slots_7_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_21
         ? _slots_9_io_out_uop_xcpt_ae_if
         : _GEN_20 ? _slots_8_io_out_uop_xcpt_ae_if : _slots_7_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_21
         ? _slots_9_io_out_uop_xcpt_ma_if
         : _GEN_20 ? _slots_8_io_out_uop_xcpt_ma_if : _slots_7_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_21
         ? _slots_9_io_out_uop_bp_debug_if
         : _GEN_20 ? _slots_8_io_out_uop_bp_debug_if : _slots_7_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_21
         ? _slots_9_io_out_uop_bp_xcpt_if
         : _GEN_20 ? _slots_8_io_out_uop_bp_xcpt_if : _slots_7_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_21
         ? _slots_9_io_out_uop_debug_fsrc
         : _GEN_20 ? _slots_8_io_out_uop_debug_fsrc : _slots_7_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_21
         ? _slots_9_io_out_uop_debug_tsrc
         : _GEN_20 ? _slots_8_io_out_uop_debug_tsrc : _slots_7_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_6_io_valid),
    .io_will_be_valid               (_slots_6_io_will_be_valid),
    .io_request                     (_slots_6_io_request),
    .io_out_uop_uopc                (_slots_6_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_6_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_6_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_6_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_6_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_6_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_6_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_6_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_6_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_6_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_6_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_6_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_6_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_6_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_6_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_6_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_6_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_6_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_6_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_6_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_6_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_6_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_6_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_6_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_6_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_6_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_6_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_6_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_6_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_6_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_6_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_6_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_6_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_6_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_6_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_6_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_6_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_6_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_6_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_6_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_6_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_6_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_6_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_6_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_6_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_6_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_6_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_6_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_6_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_6_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_6_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_6_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_6_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_6_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_6_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_6_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_6_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_6_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_6_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_6_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_6_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_6_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_6_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_6_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_6_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_6_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_6_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_6_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_6_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_6_io_uop_uopc),
    .io_uop_inst                    (_slots_6_io_uop_inst),
    .io_uop_debug_inst              (_slots_6_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_6_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_6_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_6_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_6_io_uop_fu_code),
    .io_uop_iw_state                (_slots_6_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_6_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_6_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_6_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_6_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_6_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_6_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_6_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_6_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_6_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_6_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_6_io_uop_pc_lob),
    .io_uop_taken                   (_slots_6_io_uop_taken),
    .io_uop_imm_packed              (_slots_6_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_6_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_6_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_6_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_6_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_6_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_6_io_uop_pdst),
    .io_uop_prs1                    (_slots_6_io_uop_prs1),
    .io_uop_prs2                    (_slots_6_io_uop_prs2),
    .io_uop_prs3                    (_slots_6_io_uop_prs3),
    .io_uop_ppred                   (_slots_6_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_6_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_6_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_6_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_6_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_6_io_uop_stale_pdst),
    .io_uop_exception               (_slots_6_io_uop_exception),
    .io_uop_exc_cause               (_slots_6_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_6_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_6_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_6_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_6_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_6_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_6_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_6_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_6_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_6_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_6_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_6_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_6_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_6_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_6_io_uop_ldst),
    .io_uop_lrs1                    (_slots_6_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_6_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_6_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_6_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_6_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_6_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_6_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_6_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_6_io_uop_fp_val),
    .io_uop_fp_single               (_slots_6_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_6_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_6_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_6_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_6_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_6_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_6_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_6_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_7 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_7_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_6),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_7_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_23
         ? _slots_10_io_out_uop_uopc
         : _GEN_22 ? _slots_9_io_out_uop_uopc : _slots_8_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_23
         ? _slots_10_io_out_uop_inst
         : _GEN_22 ? _slots_9_io_out_uop_inst : _slots_8_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_23
         ? _slots_10_io_out_uop_debug_inst
         : _GEN_22 ? _slots_9_io_out_uop_debug_inst : _slots_8_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_23
         ? _slots_10_io_out_uop_is_rvc
         : _GEN_22 ? _slots_9_io_out_uop_is_rvc : _slots_8_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_23
         ? _slots_10_io_out_uop_debug_pc
         : _GEN_22 ? _slots_9_io_out_uop_debug_pc : _slots_8_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_23
         ? _slots_10_io_out_uop_iq_type
         : _GEN_22 ? _slots_9_io_out_uop_iq_type : _slots_8_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_23
         ? _slots_10_io_out_uop_fu_code
         : _GEN_22 ? _slots_9_io_out_uop_fu_code : _slots_8_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_23
         ? _slots_10_io_out_uop_iw_state
         : _GEN_22 ? _slots_9_io_out_uop_iw_state : _slots_8_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_23
         ? _slots_10_io_out_uop_iw_p1_poisoned
         : _GEN_22
             ? _slots_9_io_out_uop_iw_p1_poisoned
             : _slots_8_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_23
         ? _slots_10_io_out_uop_iw_p2_poisoned
         : _GEN_22
             ? _slots_9_io_out_uop_iw_p2_poisoned
             : _slots_8_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_23
         ? _slots_10_io_out_uop_is_br
         : _GEN_22 ? _slots_9_io_out_uop_is_br : _slots_8_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_23
         ? _slots_10_io_out_uop_is_jalr
         : _GEN_22 ? _slots_9_io_out_uop_is_jalr : _slots_8_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_23
         ? _slots_10_io_out_uop_is_jal
         : _GEN_22 ? _slots_9_io_out_uop_is_jal : _slots_8_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_23
         ? _slots_10_io_out_uop_is_sfb
         : _GEN_22 ? _slots_9_io_out_uop_is_sfb : _slots_8_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_23
         ? _slots_10_io_out_uop_br_mask
         : _GEN_22 ? _slots_9_io_out_uop_br_mask : _slots_8_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_23
         ? _slots_10_io_out_uop_br_tag
         : _GEN_22 ? _slots_9_io_out_uop_br_tag : _slots_8_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_23
         ? _slots_10_io_out_uop_ftq_idx
         : _GEN_22 ? _slots_9_io_out_uop_ftq_idx : _slots_8_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_23
         ? _slots_10_io_out_uop_edge_inst
         : _GEN_22 ? _slots_9_io_out_uop_edge_inst : _slots_8_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_23
         ? _slots_10_io_out_uop_pc_lob
         : _GEN_22 ? _slots_9_io_out_uop_pc_lob : _slots_8_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_23
         ? _slots_10_io_out_uop_taken
         : _GEN_22 ? _slots_9_io_out_uop_taken : _slots_8_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_23
         ? _slots_10_io_out_uop_imm_packed
         : _GEN_22 ? _slots_9_io_out_uop_imm_packed : _slots_8_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_23
         ? _slots_10_io_out_uop_csr_addr
         : _GEN_22 ? _slots_9_io_out_uop_csr_addr : _slots_8_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_23
         ? _slots_10_io_out_uop_rob_idx
         : _GEN_22 ? _slots_9_io_out_uop_rob_idx : _slots_8_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_23
         ? _slots_10_io_out_uop_ldq_idx
         : _GEN_22 ? _slots_9_io_out_uop_ldq_idx : _slots_8_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_23
         ? _slots_10_io_out_uop_stq_idx
         : _GEN_22 ? _slots_9_io_out_uop_stq_idx : _slots_8_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_23
         ? _slots_10_io_out_uop_rxq_idx
         : _GEN_22 ? _slots_9_io_out_uop_rxq_idx : _slots_8_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_23
         ? _slots_10_io_out_uop_pdst
         : _GEN_22 ? _slots_9_io_out_uop_pdst : _slots_8_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_23
         ? _slots_10_io_out_uop_prs1
         : _GEN_22 ? _slots_9_io_out_uop_prs1 : _slots_8_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_23
         ? _slots_10_io_out_uop_prs2
         : _GEN_22 ? _slots_9_io_out_uop_prs2 : _slots_8_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_23
         ? _slots_10_io_out_uop_prs3
         : _GEN_22 ? _slots_9_io_out_uop_prs3 : _slots_8_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_23
         ? _slots_10_io_out_uop_ppred
         : _GEN_22 ? _slots_9_io_out_uop_ppred : _slots_8_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_23
         ? _slots_10_io_out_uop_prs1_busy
         : _GEN_22 ? _slots_9_io_out_uop_prs1_busy : _slots_8_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_23
         ? _slots_10_io_out_uop_prs2_busy
         : _GEN_22 ? _slots_9_io_out_uop_prs2_busy : _slots_8_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_23
         ? _slots_10_io_out_uop_prs3_busy
         : _GEN_22 ? _slots_9_io_out_uop_prs3_busy : _slots_8_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_23
         ? _slots_10_io_out_uop_ppred_busy
         : _GEN_22 ? _slots_9_io_out_uop_ppred_busy : _slots_8_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_23
         ? _slots_10_io_out_uop_stale_pdst
         : _GEN_22 ? _slots_9_io_out_uop_stale_pdst : _slots_8_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_23
         ? _slots_10_io_out_uop_exception
         : _GEN_22 ? _slots_9_io_out_uop_exception : _slots_8_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_23
         ? _slots_10_io_out_uop_exc_cause
         : _GEN_22 ? _slots_9_io_out_uop_exc_cause : _slots_8_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_23
         ? _slots_10_io_out_uop_bypassable
         : _GEN_22 ? _slots_9_io_out_uop_bypassable : _slots_8_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_23
         ? _slots_10_io_out_uop_mem_cmd
         : _GEN_22 ? _slots_9_io_out_uop_mem_cmd : _slots_8_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_23
         ? _slots_10_io_out_uop_mem_size
         : _GEN_22 ? _slots_9_io_out_uop_mem_size : _slots_8_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_23
         ? _slots_10_io_out_uop_mem_signed
         : _GEN_22 ? _slots_9_io_out_uop_mem_signed : _slots_8_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_23
         ? _slots_10_io_out_uop_is_fence
         : _GEN_22 ? _slots_9_io_out_uop_is_fence : _slots_8_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_23
         ? _slots_10_io_out_uop_is_fencei
         : _GEN_22 ? _slots_9_io_out_uop_is_fencei : _slots_8_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_23
         ? _slots_10_io_out_uop_is_amo
         : _GEN_22 ? _slots_9_io_out_uop_is_amo : _slots_8_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_23
         ? _slots_10_io_out_uop_uses_ldq
         : _GEN_22 ? _slots_9_io_out_uop_uses_ldq : _slots_8_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_23
         ? _slots_10_io_out_uop_uses_stq
         : _GEN_22 ? _slots_9_io_out_uop_uses_stq : _slots_8_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_23
         ? _slots_10_io_out_uop_is_sys_pc2epc
         : _GEN_22
             ? _slots_9_io_out_uop_is_sys_pc2epc
             : _slots_8_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_23
         ? _slots_10_io_out_uop_is_unique
         : _GEN_22 ? _slots_9_io_out_uop_is_unique : _slots_8_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_23
         ? _slots_10_io_out_uop_flush_on_commit
         : _GEN_22
             ? _slots_9_io_out_uop_flush_on_commit
             : _slots_8_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_23
         ? _slots_10_io_out_uop_ldst_is_rs1
         : _GEN_22 ? _slots_9_io_out_uop_ldst_is_rs1 : _slots_8_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_23
         ? _slots_10_io_out_uop_ldst
         : _GEN_22 ? _slots_9_io_out_uop_ldst : _slots_8_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_23
         ? _slots_10_io_out_uop_lrs1
         : _GEN_22 ? _slots_9_io_out_uop_lrs1 : _slots_8_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_23
         ? _slots_10_io_out_uop_lrs2
         : _GEN_22 ? _slots_9_io_out_uop_lrs2 : _slots_8_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_23
         ? _slots_10_io_out_uop_lrs3
         : _GEN_22 ? _slots_9_io_out_uop_lrs3 : _slots_8_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_23
         ? _slots_10_io_out_uop_ldst_val
         : _GEN_22 ? _slots_9_io_out_uop_ldst_val : _slots_8_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_23
         ? _slots_10_io_out_uop_dst_rtype
         : _GEN_22 ? _slots_9_io_out_uop_dst_rtype : _slots_8_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_23
         ? _slots_10_io_out_uop_lrs1_rtype
         : _GEN_22 ? _slots_9_io_out_uop_lrs1_rtype : _slots_8_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_23
         ? _slots_10_io_out_uop_lrs2_rtype
         : _GEN_22 ? _slots_9_io_out_uop_lrs2_rtype : _slots_8_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_23
         ? _slots_10_io_out_uop_frs3_en
         : _GEN_22 ? _slots_9_io_out_uop_frs3_en : _slots_8_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_23
         ? _slots_10_io_out_uop_fp_val
         : _GEN_22 ? _slots_9_io_out_uop_fp_val : _slots_8_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_23
         ? _slots_10_io_out_uop_fp_single
         : _GEN_22 ? _slots_9_io_out_uop_fp_single : _slots_8_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_23
         ? _slots_10_io_out_uop_xcpt_pf_if
         : _GEN_22 ? _slots_9_io_out_uop_xcpt_pf_if : _slots_8_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_23
         ? _slots_10_io_out_uop_xcpt_ae_if
         : _GEN_22 ? _slots_9_io_out_uop_xcpt_ae_if : _slots_8_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_23
         ? _slots_10_io_out_uop_xcpt_ma_if
         : _GEN_22 ? _slots_9_io_out_uop_xcpt_ma_if : _slots_8_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_23
         ? _slots_10_io_out_uop_bp_debug_if
         : _GEN_22 ? _slots_9_io_out_uop_bp_debug_if : _slots_8_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_23
         ? _slots_10_io_out_uop_bp_xcpt_if
         : _GEN_22 ? _slots_9_io_out_uop_bp_xcpt_if : _slots_8_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_23
         ? _slots_10_io_out_uop_debug_fsrc
         : _GEN_22 ? _slots_9_io_out_uop_debug_fsrc : _slots_8_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_23
         ? _slots_10_io_out_uop_debug_tsrc
         : _GEN_22 ? _slots_9_io_out_uop_debug_tsrc : _slots_8_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_7_io_valid),
    .io_will_be_valid               (_slots_7_io_will_be_valid),
    .io_request                     (_slots_7_io_request),
    .io_out_uop_uopc                (_slots_7_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_7_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_7_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_7_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_7_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_7_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_7_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_7_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_7_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_7_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_7_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_7_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_7_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_7_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_7_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_7_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_7_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_7_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_7_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_7_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_7_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_7_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_7_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_7_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_7_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_7_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_7_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_7_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_7_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_7_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_7_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_7_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_7_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_7_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_7_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_7_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_7_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_7_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_7_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_7_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_7_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_7_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_7_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_7_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_7_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_7_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_7_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_7_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_7_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_7_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_7_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_7_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_7_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_7_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_7_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_7_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_7_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_7_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_7_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_7_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_7_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_7_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_7_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_7_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_7_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_7_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_7_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_7_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_7_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_7_io_uop_uopc),
    .io_uop_inst                    (_slots_7_io_uop_inst),
    .io_uop_debug_inst              (_slots_7_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_7_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_7_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_7_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_7_io_uop_fu_code),
    .io_uop_iw_state                (_slots_7_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_7_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_7_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_7_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_7_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_7_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_7_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_7_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_7_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_7_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_7_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_7_io_uop_pc_lob),
    .io_uop_taken                   (_slots_7_io_uop_taken),
    .io_uop_imm_packed              (_slots_7_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_7_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_7_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_7_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_7_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_7_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_7_io_uop_pdst),
    .io_uop_prs1                    (_slots_7_io_uop_prs1),
    .io_uop_prs2                    (_slots_7_io_uop_prs2),
    .io_uop_prs3                    (_slots_7_io_uop_prs3),
    .io_uop_ppred                   (_slots_7_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_7_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_7_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_7_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_7_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_7_io_uop_stale_pdst),
    .io_uop_exception               (_slots_7_io_uop_exception),
    .io_uop_exc_cause               (_slots_7_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_7_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_7_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_7_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_7_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_7_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_7_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_7_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_7_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_7_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_7_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_7_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_7_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_7_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_7_io_uop_ldst),
    .io_uop_lrs1                    (_slots_7_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_7_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_7_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_7_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_7_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_7_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_7_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_7_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_7_io_uop_fp_val),
    .io_uop_fp_single               (_slots_7_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_7_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_7_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_7_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_7_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_7_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_7_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_7_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_8 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_8_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_7),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_8_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_25
         ? _slots_11_io_out_uop_uopc
         : _GEN_24 ? _slots_10_io_out_uop_uopc : _slots_9_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_25
         ? _slots_11_io_out_uop_inst
         : _GEN_24 ? _slots_10_io_out_uop_inst : _slots_9_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_25
         ? _slots_11_io_out_uop_debug_inst
         : _GEN_24 ? _slots_10_io_out_uop_debug_inst : _slots_9_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_25
         ? _slots_11_io_out_uop_is_rvc
         : _GEN_24 ? _slots_10_io_out_uop_is_rvc : _slots_9_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_25
         ? _slots_11_io_out_uop_debug_pc
         : _GEN_24 ? _slots_10_io_out_uop_debug_pc : _slots_9_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_25
         ? _slots_11_io_out_uop_iq_type
         : _GEN_24 ? _slots_10_io_out_uop_iq_type : _slots_9_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_25
         ? _slots_11_io_out_uop_fu_code
         : _GEN_24 ? _slots_10_io_out_uop_fu_code : _slots_9_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_25
         ? _slots_11_io_out_uop_iw_state
         : _GEN_24 ? _slots_10_io_out_uop_iw_state : _slots_9_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_25
         ? _slots_11_io_out_uop_iw_p1_poisoned
         : _GEN_24
             ? _slots_10_io_out_uop_iw_p1_poisoned
             : _slots_9_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_25
         ? _slots_11_io_out_uop_iw_p2_poisoned
         : _GEN_24
             ? _slots_10_io_out_uop_iw_p2_poisoned
             : _slots_9_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_25
         ? _slots_11_io_out_uop_is_br
         : _GEN_24 ? _slots_10_io_out_uop_is_br : _slots_9_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_25
         ? _slots_11_io_out_uop_is_jalr
         : _GEN_24 ? _slots_10_io_out_uop_is_jalr : _slots_9_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_25
         ? _slots_11_io_out_uop_is_jal
         : _GEN_24 ? _slots_10_io_out_uop_is_jal : _slots_9_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_25
         ? _slots_11_io_out_uop_is_sfb
         : _GEN_24 ? _slots_10_io_out_uop_is_sfb : _slots_9_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_25
         ? _slots_11_io_out_uop_br_mask
         : _GEN_24 ? _slots_10_io_out_uop_br_mask : _slots_9_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_25
         ? _slots_11_io_out_uop_br_tag
         : _GEN_24 ? _slots_10_io_out_uop_br_tag : _slots_9_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_25
         ? _slots_11_io_out_uop_ftq_idx
         : _GEN_24 ? _slots_10_io_out_uop_ftq_idx : _slots_9_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_25
         ? _slots_11_io_out_uop_edge_inst
         : _GEN_24 ? _slots_10_io_out_uop_edge_inst : _slots_9_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_25
         ? _slots_11_io_out_uop_pc_lob
         : _GEN_24 ? _slots_10_io_out_uop_pc_lob : _slots_9_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_25
         ? _slots_11_io_out_uop_taken
         : _GEN_24 ? _slots_10_io_out_uop_taken : _slots_9_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_25
         ? _slots_11_io_out_uop_imm_packed
         : _GEN_24 ? _slots_10_io_out_uop_imm_packed : _slots_9_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_25
         ? _slots_11_io_out_uop_csr_addr
         : _GEN_24 ? _slots_10_io_out_uop_csr_addr : _slots_9_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_25
         ? _slots_11_io_out_uop_rob_idx
         : _GEN_24 ? _slots_10_io_out_uop_rob_idx : _slots_9_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_25
         ? _slots_11_io_out_uop_ldq_idx
         : _GEN_24 ? _slots_10_io_out_uop_ldq_idx : _slots_9_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_25
         ? _slots_11_io_out_uop_stq_idx
         : _GEN_24 ? _slots_10_io_out_uop_stq_idx : _slots_9_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_25
         ? _slots_11_io_out_uop_rxq_idx
         : _GEN_24 ? _slots_10_io_out_uop_rxq_idx : _slots_9_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_25
         ? _slots_11_io_out_uop_pdst
         : _GEN_24 ? _slots_10_io_out_uop_pdst : _slots_9_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_25
         ? _slots_11_io_out_uop_prs1
         : _GEN_24 ? _slots_10_io_out_uop_prs1 : _slots_9_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_25
         ? _slots_11_io_out_uop_prs2
         : _GEN_24 ? _slots_10_io_out_uop_prs2 : _slots_9_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_25
         ? _slots_11_io_out_uop_prs3
         : _GEN_24 ? _slots_10_io_out_uop_prs3 : _slots_9_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_25
         ? _slots_11_io_out_uop_ppred
         : _GEN_24 ? _slots_10_io_out_uop_ppred : _slots_9_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_25
         ? _slots_11_io_out_uop_prs1_busy
         : _GEN_24 ? _slots_10_io_out_uop_prs1_busy : _slots_9_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_25
         ? _slots_11_io_out_uop_prs2_busy
         : _GEN_24 ? _slots_10_io_out_uop_prs2_busy : _slots_9_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_25
         ? _slots_11_io_out_uop_prs3_busy
         : _GEN_24 ? _slots_10_io_out_uop_prs3_busy : _slots_9_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_25
         ? _slots_11_io_out_uop_ppred_busy
         : _GEN_24 ? _slots_10_io_out_uop_ppred_busy : _slots_9_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_25
         ? _slots_11_io_out_uop_stale_pdst
         : _GEN_24 ? _slots_10_io_out_uop_stale_pdst : _slots_9_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_25
         ? _slots_11_io_out_uop_exception
         : _GEN_24 ? _slots_10_io_out_uop_exception : _slots_9_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_25
         ? _slots_11_io_out_uop_exc_cause
         : _GEN_24 ? _slots_10_io_out_uop_exc_cause : _slots_9_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_25
         ? _slots_11_io_out_uop_bypassable
         : _GEN_24 ? _slots_10_io_out_uop_bypassable : _slots_9_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_25
         ? _slots_11_io_out_uop_mem_cmd
         : _GEN_24 ? _slots_10_io_out_uop_mem_cmd : _slots_9_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_25
         ? _slots_11_io_out_uop_mem_size
         : _GEN_24 ? _slots_10_io_out_uop_mem_size : _slots_9_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_25
         ? _slots_11_io_out_uop_mem_signed
         : _GEN_24 ? _slots_10_io_out_uop_mem_signed : _slots_9_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_25
         ? _slots_11_io_out_uop_is_fence
         : _GEN_24 ? _slots_10_io_out_uop_is_fence : _slots_9_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_25
         ? _slots_11_io_out_uop_is_fencei
         : _GEN_24 ? _slots_10_io_out_uop_is_fencei : _slots_9_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_25
         ? _slots_11_io_out_uop_is_amo
         : _GEN_24 ? _slots_10_io_out_uop_is_amo : _slots_9_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_25
         ? _slots_11_io_out_uop_uses_ldq
         : _GEN_24 ? _slots_10_io_out_uop_uses_ldq : _slots_9_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_25
         ? _slots_11_io_out_uop_uses_stq
         : _GEN_24 ? _slots_10_io_out_uop_uses_stq : _slots_9_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_25
         ? _slots_11_io_out_uop_is_sys_pc2epc
         : _GEN_24
             ? _slots_10_io_out_uop_is_sys_pc2epc
             : _slots_9_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_25
         ? _slots_11_io_out_uop_is_unique
         : _GEN_24 ? _slots_10_io_out_uop_is_unique : _slots_9_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_25
         ? _slots_11_io_out_uop_flush_on_commit
         : _GEN_24
             ? _slots_10_io_out_uop_flush_on_commit
             : _slots_9_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_25
         ? _slots_11_io_out_uop_ldst_is_rs1
         : _GEN_24 ? _slots_10_io_out_uop_ldst_is_rs1 : _slots_9_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_25
         ? _slots_11_io_out_uop_ldst
         : _GEN_24 ? _slots_10_io_out_uop_ldst : _slots_9_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_25
         ? _slots_11_io_out_uop_lrs1
         : _GEN_24 ? _slots_10_io_out_uop_lrs1 : _slots_9_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_25
         ? _slots_11_io_out_uop_lrs2
         : _GEN_24 ? _slots_10_io_out_uop_lrs2 : _slots_9_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_25
         ? _slots_11_io_out_uop_lrs3
         : _GEN_24 ? _slots_10_io_out_uop_lrs3 : _slots_9_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_25
         ? _slots_11_io_out_uop_ldst_val
         : _GEN_24 ? _slots_10_io_out_uop_ldst_val : _slots_9_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_25
         ? _slots_11_io_out_uop_dst_rtype
         : _GEN_24 ? _slots_10_io_out_uop_dst_rtype : _slots_9_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_25
         ? _slots_11_io_out_uop_lrs1_rtype
         : _GEN_24 ? _slots_10_io_out_uop_lrs1_rtype : _slots_9_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_25
         ? _slots_11_io_out_uop_lrs2_rtype
         : _GEN_24 ? _slots_10_io_out_uop_lrs2_rtype : _slots_9_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_25
         ? _slots_11_io_out_uop_frs3_en
         : _GEN_24 ? _slots_10_io_out_uop_frs3_en : _slots_9_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_25
         ? _slots_11_io_out_uop_fp_val
         : _GEN_24 ? _slots_10_io_out_uop_fp_val : _slots_9_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_25
         ? _slots_11_io_out_uop_fp_single
         : _GEN_24 ? _slots_10_io_out_uop_fp_single : _slots_9_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_25
         ? _slots_11_io_out_uop_xcpt_pf_if
         : _GEN_24 ? _slots_10_io_out_uop_xcpt_pf_if : _slots_9_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_25
         ? _slots_11_io_out_uop_xcpt_ae_if
         : _GEN_24 ? _slots_10_io_out_uop_xcpt_ae_if : _slots_9_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_25
         ? _slots_11_io_out_uop_xcpt_ma_if
         : _GEN_24 ? _slots_10_io_out_uop_xcpt_ma_if : _slots_9_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_25
         ? _slots_11_io_out_uop_bp_debug_if
         : _GEN_24 ? _slots_10_io_out_uop_bp_debug_if : _slots_9_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_25
         ? _slots_11_io_out_uop_bp_xcpt_if
         : _GEN_24 ? _slots_10_io_out_uop_bp_xcpt_if : _slots_9_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_25
         ? _slots_11_io_out_uop_debug_fsrc
         : _GEN_24 ? _slots_10_io_out_uop_debug_fsrc : _slots_9_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_25
         ? _slots_11_io_out_uop_debug_tsrc
         : _GEN_24 ? _slots_10_io_out_uop_debug_tsrc : _slots_9_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_8_io_valid),
    .io_will_be_valid               (_slots_8_io_will_be_valid),
    .io_request                     (_slots_8_io_request),
    .io_out_uop_uopc                (_slots_8_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_8_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_8_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_8_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_8_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_8_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_8_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_8_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_8_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_8_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_8_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_8_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_8_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_8_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_8_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_8_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_8_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_8_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_8_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_8_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_8_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_8_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_8_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_8_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_8_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_8_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_8_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_8_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_8_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_8_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_8_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_8_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_8_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_8_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_8_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_8_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_8_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_8_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_8_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_8_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_8_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_8_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_8_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_8_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_8_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_8_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_8_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_8_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_8_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_8_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_8_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_8_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_8_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_8_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_8_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_8_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_8_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_8_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_8_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_8_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_8_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_8_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_8_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_8_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_8_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_8_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_8_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_8_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_8_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_8_io_uop_uopc),
    .io_uop_inst                    (_slots_8_io_uop_inst),
    .io_uop_debug_inst              (_slots_8_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_8_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_8_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_8_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_8_io_uop_fu_code),
    .io_uop_iw_state                (_slots_8_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_8_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_8_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_8_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_8_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_8_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_8_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_8_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_8_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_8_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_8_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_8_io_uop_pc_lob),
    .io_uop_taken                   (_slots_8_io_uop_taken),
    .io_uop_imm_packed              (_slots_8_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_8_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_8_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_8_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_8_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_8_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_8_io_uop_pdst),
    .io_uop_prs1                    (_slots_8_io_uop_prs1),
    .io_uop_prs2                    (_slots_8_io_uop_prs2),
    .io_uop_prs3                    (_slots_8_io_uop_prs3),
    .io_uop_ppred                   (_slots_8_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_8_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_8_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_8_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_8_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_8_io_uop_stale_pdst),
    .io_uop_exception               (_slots_8_io_uop_exception),
    .io_uop_exc_cause               (_slots_8_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_8_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_8_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_8_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_8_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_8_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_8_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_8_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_8_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_8_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_8_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_8_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_8_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_8_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_8_io_uop_ldst),
    .io_uop_lrs1                    (_slots_8_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_8_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_8_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_8_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_8_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_8_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_8_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_8_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_8_io_uop_fp_val),
    .io_uop_fp_single               (_slots_8_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_8_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_8_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_8_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_8_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_8_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_8_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_8_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_9 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_9_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_8),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_9_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_27
         ? _slots_12_io_out_uop_uopc
         : _GEN_26 ? _slots_11_io_out_uop_uopc : _slots_10_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_27
         ? _slots_12_io_out_uop_inst
         : _GEN_26 ? _slots_11_io_out_uop_inst : _slots_10_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_27
         ? _slots_12_io_out_uop_debug_inst
         : _GEN_26 ? _slots_11_io_out_uop_debug_inst : _slots_10_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_27
         ? _slots_12_io_out_uop_is_rvc
         : _GEN_26 ? _slots_11_io_out_uop_is_rvc : _slots_10_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_27
         ? _slots_12_io_out_uop_debug_pc
         : _GEN_26 ? _slots_11_io_out_uop_debug_pc : _slots_10_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_27
         ? _slots_12_io_out_uop_iq_type
         : _GEN_26 ? _slots_11_io_out_uop_iq_type : _slots_10_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_27
         ? _slots_12_io_out_uop_fu_code
         : _GEN_26 ? _slots_11_io_out_uop_fu_code : _slots_10_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_27
         ? _slots_12_io_out_uop_iw_state
         : _GEN_26 ? _slots_11_io_out_uop_iw_state : _slots_10_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_27
         ? _slots_12_io_out_uop_iw_p1_poisoned
         : _GEN_26
             ? _slots_11_io_out_uop_iw_p1_poisoned
             : _slots_10_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_27
         ? _slots_12_io_out_uop_iw_p2_poisoned
         : _GEN_26
             ? _slots_11_io_out_uop_iw_p2_poisoned
             : _slots_10_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_27
         ? _slots_12_io_out_uop_is_br
         : _GEN_26 ? _slots_11_io_out_uop_is_br : _slots_10_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_27
         ? _slots_12_io_out_uop_is_jalr
         : _GEN_26 ? _slots_11_io_out_uop_is_jalr : _slots_10_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_27
         ? _slots_12_io_out_uop_is_jal
         : _GEN_26 ? _slots_11_io_out_uop_is_jal : _slots_10_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_27
         ? _slots_12_io_out_uop_is_sfb
         : _GEN_26 ? _slots_11_io_out_uop_is_sfb : _slots_10_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_27
         ? _slots_12_io_out_uop_br_mask
         : _GEN_26 ? _slots_11_io_out_uop_br_mask : _slots_10_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_27
         ? _slots_12_io_out_uop_br_tag
         : _GEN_26 ? _slots_11_io_out_uop_br_tag : _slots_10_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_27
         ? _slots_12_io_out_uop_ftq_idx
         : _GEN_26 ? _slots_11_io_out_uop_ftq_idx : _slots_10_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_27
         ? _slots_12_io_out_uop_edge_inst
         : _GEN_26 ? _slots_11_io_out_uop_edge_inst : _slots_10_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_27
         ? _slots_12_io_out_uop_pc_lob
         : _GEN_26 ? _slots_11_io_out_uop_pc_lob : _slots_10_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_27
         ? _slots_12_io_out_uop_taken
         : _GEN_26 ? _slots_11_io_out_uop_taken : _slots_10_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_27
         ? _slots_12_io_out_uop_imm_packed
         : _GEN_26 ? _slots_11_io_out_uop_imm_packed : _slots_10_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_27
         ? _slots_12_io_out_uop_csr_addr
         : _GEN_26 ? _slots_11_io_out_uop_csr_addr : _slots_10_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_27
         ? _slots_12_io_out_uop_rob_idx
         : _GEN_26 ? _slots_11_io_out_uop_rob_idx : _slots_10_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_27
         ? _slots_12_io_out_uop_ldq_idx
         : _GEN_26 ? _slots_11_io_out_uop_ldq_idx : _slots_10_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_27
         ? _slots_12_io_out_uop_stq_idx
         : _GEN_26 ? _slots_11_io_out_uop_stq_idx : _slots_10_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_27
         ? _slots_12_io_out_uop_rxq_idx
         : _GEN_26 ? _slots_11_io_out_uop_rxq_idx : _slots_10_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_27
         ? _slots_12_io_out_uop_pdst
         : _GEN_26 ? _slots_11_io_out_uop_pdst : _slots_10_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_27
         ? _slots_12_io_out_uop_prs1
         : _GEN_26 ? _slots_11_io_out_uop_prs1 : _slots_10_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_27
         ? _slots_12_io_out_uop_prs2
         : _GEN_26 ? _slots_11_io_out_uop_prs2 : _slots_10_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_27
         ? _slots_12_io_out_uop_prs3
         : _GEN_26 ? _slots_11_io_out_uop_prs3 : _slots_10_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_27
         ? _slots_12_io_out_uop_ppred
         : _GEN_26 ? _slots_11_io_out_uop_ppred : _slots_10_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_27
         ? _slots_12_io_out_uop_prs1_busy
         : _GEN_26 ? _slots_11_io_out_uop_prs1_busy : _slots_10_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_27
         ? _slots_12_io_out_uop_prs2_busy
         : _GEN_26 ? _slots_11_io_out_uop_prs2_busy : _slots_10_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_27
         ? _slots_12_io_out_uop_prs3_busy
         : _GEN_26 ? _slots_11_io_out_uop_prs3_busy : _slots_10_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_27
         ? _slots_12_io_out_uop_ppred_busy
         : _GEN_26 ? _slots_11_io_out_uop_ppred_busy : _slots_10_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_27
         ? _slots_12_io_out_uop_stale_pdst
         : _GEN_26 ? _slots_11_io_out_uop_stale_pdst : _slots_10_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_27
         ? _slots_12_io_out_uop_exception
         : _GEN_26 ? _slots_11_io_out_uop_exception : _slots_10_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_27
         ? _slots_12_io_out_uop_exc_cause
         : _GEN_26 ? _slots_11_io_out_uop_exc_cause : _slots_10_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_27
         ? _slots_12_io_out_uop_bypassable
         : _GEN_26 ? _slots_11_io_out_uop_bypassable : _slots_10_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_27
         ? _slots_12_io_out_uop_mem_cmd
         : _GEN_26 ? _slots_11_io_out_uop_mem_cmd : _slots_10_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_27
         ? _slots_12_io_out_uop_mem_size
         : _GEN_26 ? _slots_11_io_out_uop_mem_size : _slots_10_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_27
         ? _slots_12_io_out_uop_mem_signed
         : _GEN_26 ? _slots_11_io_out_uop_mem_signed : _slots_10_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_27
         ? _slots_12_io_out_uop_is_fence
         : _GEN_26 ? _slots_11_io_out_uop_is_fence : _slots_10_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_27
         ? _slots_12_io_out_uop_is_fencei
         : _GEN_26 ? _slots_11_io_out_uop_is_fencei : _slots_10_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_27
         ? _slots_12_io_out_uop_is_amo
         : _GEN_26 ? _slots_11_io_out_uop_is_amo : _slots_10_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_27
         ? _slots_12_io_out_uop_uses_ldq
         : _GEN_26 ? _slots_11_io_out_uop_uses_ldq : _slots_10_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_27
         ? _slots_12_io_out_uop_uses_stq
         : _GEN_26 ? _slots_11_io_out_uop_uses_stq : _slots_10_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_27
         ? _slots_12_io_out_uop_is_sys_pc2epc
         : _GEN_26
             ? _slots_11_io_out_uop_is_sys_pc2epc
             : _slots_10_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_27
         ? _slots_12_io_out_uop_is_unique
         : _GEN_26 ? _slots_11_io_out_uop_is_unique : _slots_10_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_27
         ? _slots_12_io_out_uop_flush_on_commit
         : _GEN_26
             ? _slots_11_io_out_uop_flush_on_commit
             : _slots_10_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_27
         ? _slots_12_io_out_uop_ldst_is_rs1
         : _GEN_26 ? _slots_11_io_out_uop_ldst_is_rs1 : _slots_10_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_27
         ? _slots_12_io_out_uop_ldst
         : _GEN_26 ? _slots_11_io_out_uop_ldst : _slots_10_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_27
         ? _slots_12_io_out_uop_lrs1
         : _GEN_26 ? _slots_11_io_out_uop_lrs1 : _slots_10_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_27
         ? _slots_12_io_out_uop_lrs2
         : _GEN_26 ? _slots_11_io_out_uop_lrs2 : _slots_10_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_27
         ? _slots_12_io_out_uop_lrs3
         : _GEN_26 ? _slots_11_io_out_uop_lrs3 : _slots_10_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_27
         ? _slots_12_io_out_uop_ldst_val
         : _GEN_26 ? _slots_11_io_out_uop_ldst_val : _slots_10_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_27
         ? _slots_12_io_out_uop_dst_rtype
         : _GEN_26 ? _slots_11_io_out_uop_dst_rtype : _slots_10_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_27
         ? _slots_12_io_out_uop_lrs1_rtype
         : _GEN_26 ? _slots_11_io_out_uop_lrs1_rtype : _slots_10_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_27
         ? _slots_12_io_out_uop_lrs2_rtype
         : _GEN_26 ? _slots_11_io_out_uop_lrs2_rtype : _slots_10_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_27
         ? _slots_12_io_out_uop_frs3_en
         : _GEN_26 ? _slots_11_io_out_uop_frs3_en : _slots_10_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_27
         ? _slots_12_io_out_uop_fp_val
         : _GEN_26 ? _slots_11_io_out_uop_fp_val : _slots_10_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_27
         ? _slots_12_io_out_uop_fp_single
         : _GEN_26 ? _slots_11_io_out_uop_fp_single : _slots_10_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_27
         ? _slots_12_io_out_uop_xcpt_pf_if
         : _GEN_26 ? _slots_11_io_out_uop_xcpt_pf_if : _slots_10_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_27
         ? _slots_12_io_out_uop_xcpt_ae_if
         : _GEN_26 ? _slots_11_io_out_uop_xcpt_ae_if : _slots_10_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_27
         ? _slots_12_io_out_uop_xcpt_ma_if
         : _GEN_26 ? _slots_11_io_out_uop_xcpt_ma_if : _slots_10_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_27
         ? _slots_12_io_out_uop_bp_debug_if
         : _GEN_26 ? _slots_11_io_out_uop_bp_debug_if : _slots_10_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_27
         ? _slots_12_io_out_uop_bp_xcpt_if
         : _GEN_26 ? _slots_11_io_out_uop_bp_xcpt_if : _slots_10_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_27
         ? _slots_12_io_out_uop_debug_fsrc
         : _GEN_26 ? _slots_11_io_out_uop_debug_fsrc : _slots_10_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_27
         ? _slots_12_io_out_uop_debug_tsrc
         : _GEN_26 ? _slots_11_io_out_uop_debug_tsrc : _slots_10_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_9_io_valid),
    .io_will_be_valid               (_slots_9_io_will_be_valid),
    .io_request                     (_slots_9_io_request),
    .io_out_uop_uopc                (_slots_9_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_9_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_9_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_9_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_9_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_9_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_9_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_9_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_9_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_9_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_9_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_9_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_9_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_9_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_9_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_9_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_9_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_9_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_9_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_9_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_9_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_9_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_9_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_9_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_9_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_9_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_9_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_9_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_9_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_9_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_9_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_9_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_9_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_9_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_9_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_9_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_9_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_9_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_9_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_9_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_9_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_9_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_9_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_9_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_9_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_9_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_9_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_9_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_9_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_9_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_9_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_9_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_9_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_9_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_9_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_9_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_9_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_9_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_9_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_9_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_9_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_9_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_9_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_9_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_9_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_9_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_9_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_9_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_9_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_9_io_uop_uopc),
    .io_uop_inst                    (_slots_9_io_uop_inst),
    .io_uop_debug_inst              (_slots_9_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_9_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_9_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_9_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_9_io_uop_fu_code),
    .io_uop_iw_state                (_slots_9_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_9_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_9_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_9_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_9_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_9_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_9_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_9_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_9_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_9_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_9_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_9_io_uop_pc_lob),
    .io_uop_taken                   (_slots_9_io_uop_taken),
    .io_uop_imm_packed              (_slots_9_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_9_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_9_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_9_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_9_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_9_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_9_io_uop_pdst),
    .io_uop_prs1                    (_slots_9_io_uop_prs1),
    .io_uop_prs2                    (_slots_9_io_uop_prs2),
    .io_uop_prs3                    (_slots_9_io_uop_prs3),
    .io_uop_ppred                   (_slots_9_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_9_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_9_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_9_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_9_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_9_io_uop_stale_pdst),
    .io_uop_exception               (_slots_9_io_uop_exception),
    .io_uop_exc_cause               (_slots_9_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_9_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_9_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_9_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_9_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_9_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_9_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_9_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_9_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_9_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_9_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_9_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_9_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_9_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_9_io_uop_ldst),
    .io_uop_lrs1                    (_slots_9_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_9_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_9_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_9_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_9_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_9_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_9_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_9_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_9_io_uop_fp_val),
    .io_uop_fp_single               (_slots_9_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_9_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_9_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_9_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_9_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_9_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_9_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_9_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_10 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_10_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_9),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_10_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_29
         ? _slots_13_io_out_uop_uopc
         : _GEN_28 ? _slots_12_io_out_uop_uopc : _slots_11_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_29
         ? _slots_13_io_out_uop_inst
         : _GEN_28 ? _slots_12_io_out_uop_inst : _slots_11_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_29
         ? _slots_13_io_out_uop_debug_inst
         : _GEN_28 ? _slots_12_io_out_uop_debug_inst : _slots_11_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_29
         ? _slots_13_io_out_uop_is_rvc
         : _GEN_28 ? _slots_12_io_out_uop_is_rvc : _slots_11_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_29
         ? _slots_13_io_out_uop_debug_pc
         : _GEN_28 ? _slots_12_io_out_uop_debug_pc : _slots_11_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_29
         ? _slots_13_io_out_uop_iq_type
         : _GEN_28 ? _slots_12_io_out_uop_iq_type : _slots_11_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_29
         ? _slots_13_io_out_uop_fu_code
         : _GEN_28 ? _slots_12_io_out_uop_fu_code : _slots_11_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_29
         ? _slots_13_io_out_uop_iw_state
         : _GEN_28 ? _slots_12_io_out_uop_iw_state : _slots_11_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_29
         ? _slots_13_io_out_uop_iw_p1_poisoned
         : _GEN_28
             ? _slots_12_io_out_uop_iw_p1_poisoned
             : _slots_11_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_29
         ? _slots_13_io_out_uop_iw_p2_poisoned
         : _GEN_28
             ? _slots_12_io_out_uop_iw_p2_poisoned
             : _slots_11_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_29
         ? _slots_13_io_out_uop_is_br
         : _GEN_28 ? _slots_12_io_out_uop_is_br : _slots_11_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_29
         ? _slots_13_io_out_uop_is_jalr
         : _GEN_28 ? _slots_12_io_out_uop_is_jalr : _slots_11_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_29
         ? _slots_13_io_out_uop_is_jal
         : _GEN_28 ? _slots_12_io_out_uop_is_jal : _slots_11_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_29
         ? _slots_13_io_out_uop_is_sfb
         : _GEN_28 ? _slots_12_io_out_uop_is_sfb : _slots_11_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_29
         ? _slots_13_io_out_uop_br_mask
         : _GEN_28 ? _slots_12_io_out_uop_br_mask : _slots_11_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_29
         ? _slots_13_io_out_uop_br_tag
         : _GEN_28 ? _slots_12_io_out_uop_br_tag : _slots_11_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_29
         ? _slots_13_io_out_uop_ftq_idx
         : _GEN_28 ? _slots_12_io_out_uop_ftq_idx : _slots_11_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_29
         ? _slots_13_io_out_uop_edge_inst
         : _GEN_28 ? _slots_12_io_out_uop_edge_inst : _slots_11_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_29
         ? _slots_13_io_out_uop_pc_lob
         : _GEN_28 ? _slots_12_io_out_uop_pc_lob : _slots_11_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_29
         ? _slots_13_io_out_uop_taken
         : _GEN_28 ? _slots_12_io_out_uop_taken : _slots_11_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_29
         ? _slots_13_io_out_uop_imm_packed
         : _GEN_28 ? _slots_12_io_out_uop_imm_packed : _slots_11_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_29
         ? _slots_13_io_out_uop_csr_addr
         : _GEN_28 ? _slots_12_io_out_uop_csr_addr : _slots_11_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_29
         ? _slots_13_io_out_uop_rob_idx
         : _GEN_28 ? _slots_12_io_out_uop_rob_idx : _slots_11_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_29
         ? _slots_13_io_out_uop_ldq_idx
         : _GEN_28 ? _slots_12_io_out_uop_ldq_idx : _slots_11_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_29
         ? _slots_13_io_out_uop_stq_idx
         : _GEN_28 ? _slots_12_io_out_uop_stq_idx : _slots_11_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_29
         ? _slots_13_io_out_uop_rxq_idx
         : _GEN_28 ? _slots_12_io_out_uop_rxq_idx : _slots_11_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_29
         ? _slots_13_io_out_uop_pdst
         : _GEN_28 ? _slots_12_io_out_uop_pdst : _slots_11_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_29
         ? _slots_13_io_out_uop_prs1
         : _GEN_28 ? _slots_12_io_out_uop_prs1 : _slots_11_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_29
         ? _slots_13_io_out_uop_prs2
         : _GEN_28 ? _slots_12_io_out_uop_prs2 : _slots_11_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_29
         ? _slots_13_io_out_uop_prs3
         : _GEN_28 ? _slots_12_io_out_uop_prs3 : _slots_11_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_29
         ? _slots_13_io_out_uop_ppred
         : _GEN_28 ? _slots_12_io_out_uop_ppred : _slots_11_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_29
         ? _slots_13_io_out_uop_prs1_busy
         : _GEN_28 ? _slots_12_io_out_uop_prs1_busy : _slots_11_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_29
         ? _slots_13_io_out_uop_prs2_busy
         : _GEN_28 ? _slots_12_io_out_uop_prs2_busy : _slots_11_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_29
         ? _slots_13_io_out_uop_prs3_busy
         : _GEN_28 ? _slots_12_io_out_uop_prs3_busy : _slots_11_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_29
         ? _slots_13_io_out_uop_ppred_busy
         : _GEN_28 ? _slots_12_io_out_uop_ppred_busy : _slots_11_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_29
         ? _slots_13_io_out_uop_stale_pdst
         : _GEN_28 ? _slots_12_io_out_uop_stale_pdst : _slots_11_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_29
         ? _slots_13_io_out_uop_exception
         : _GEN_28 ? _slots_12_io_out_uop_exception : _slots_11_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_29
         ? _slots_13_io_out_uop_exc_cause
         : _GEN_28 ? _slots_12_io_out_uop_exc_cause : _slots_11_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_29
         ? _slots_13_io_out_uop_bypassable
         : _GEN_28 ? _slots_12_io_out_uop_bypassable : _slots_11_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_29
         ? _slots_13_io_out_uop_mem_cmd
         : _GEN_28 ? _slots_12_io_out_uop_mem_cmd : _slots_11_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_29
         ? _slots_13_io_out_uop_mem_size
         : _GEN_28 ? _slots_12_io_out_uop_mem_size : _slots_11_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_29
         ? _slots_13_io_out_uop_mem_signed
         : _GEN_28 ? _slots_12_io_out_uop_mem_signed : _slots_11_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_29
         ? _slots_13_io_out_uop_is_fence
         : _GEN_28 ? _slots_12_io_out_uop_is_fence : _slots_11_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_29
         ? _slots_13_io_out_uop_is_fencei
         : _GEN_28 ? _slots_12_io_out_uop_is_fencei : _slots_11_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_29
         ? _slots_13_io_out_uop_is_amo
         : _GEN_28 ? _slots_12_io_out_uop_is_amo : _slots_11_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_29
         ? _slots_13_io_out_uop_uses_ldq
         : _GEN_28 ? _slots_12_io_out_uop_uses_ldq : _slots_11_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_29
         ? _slots_13_io_out_uop_uses_stq
         : _GEN_28 ? _slots_12_io_out_uop_uses_stq : _slots_11_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_29
         ? _slots_13_io_out_uop_is_sys_pc2epc
         : _GEN_28
             ? _slots_12_io_out_uop_is_sys_pc2epc
             : _slots_11_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_29
         ? _slots_13_io_out_uop_is_unique
         : _GEN_28 ? _slots_12_io_out_uop_is_unique : _slots_11_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_29
         ? _slots_13_io_out_uop_flush_on_commit
         : _GEN_28
             ? _slots_12_io_out_uop_flush_on_commit
             : _slots_11_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_29
         ? _slots_13_io_out_uop_ldst_is_rs1
         : _GEN_28 ? _slots_12_io_out_uop_ldst_is_rs1 : _slots_11_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_29
         ? _slots_13_io_out_uop_ldst
         : _GEN_28 ? _slots_12_io_out_uop_ldst : _slots_11_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_29
         ? _slots_13_io_out_uop_lrs1
         : _GEN_28 ? _slots_12_io_out_uop_lrs1 : _slots_11_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_29
         ? _slots_13_io_out_uop_lrs2
         : _GEN_28 ? _slots_12_io_out_uop_lrs2 : _slots_11_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_29
         ? _slots_13_io_out_uop_lrs3
         : _GEN_28 ? _slots_12_io_out_uop_lrs3 : _slots_11_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_29
         ? _slots_13_io_out_uop_ldst_val
         : _GEN_28 ? _slots_12_io_out_uop_ldst_val : _slots_11_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_29
         ? _slots_13_io_out_uop_dst_rtype
         : _GEN_28 ? _slots_12_io_out_uop_dst_rtype : _slots_11_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_29
         ? _slots_13_io_out_uop_lrs1_rtype
         : _GEN_28 ? _slots_12_io_out_uop_lrs1_rtype : _slots_11_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_29
         ? _slots_13_io_out_uop_lrs2_rtype
         : _GEN_28 ? _slots_12_io_out_uop_lrs2_rtype : _slots_11_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_29
         ? _slots_13_io_out_uop_frs3_en
         : _GEN_28 ? _slots_12_io_out_uop_frs3_en : _slots_11_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_29
         ? _slots_13_io_out_uop_fp_val
         : _GEN_28 ? _slots_12_io_out_uop_fp_val : _slots_11_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_29
         ? _slots_13_io_out_uop_fp_single
         : _GEN_28 ? _slots_12_io_out_uop_fp_single : _slots_11_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_29
         ? _slots_13_io_out_uop_xcpt_pf_if
         : _GEN_28 ? _slots_12_io_out_uop_xcpt_pf_if : _slots_11_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_29
         ? _slots_13_io_out_uop_xcpt_ae_if
         : _GEN_28 ? _slots_12_io_out_uop_xcpt_ae_if : _slots_11_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_29
         ? _slots_13_io_out_uop_xcpt_ma_if
         : _GEN_28 ? _slots_12_io_out_uop_xcpt_ma_if : _slots_11_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_29
         ? _slots_13_io_out_uop_bp_debug_if
         : _GEN_28 ? _slots_12_io_out_uop_bp_debug_if : _slots_11_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_29
         ? _slots_13_io_out_uop_bp_xcpt_if
         : _GEN_28 ? _slots_12_io_out_uop_bp_xcpt_if : _slots_11_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_29
         ? _slots_13_io_out_uop_debug_fsrc
         : _GEN_28 ? _slots_12_io_out_uop_debug_fsrc : _slots_11_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_29
         ? _slots_13_io_out_uop_debug_tsrc
         : _GEN_28 ? _slots_12_io_out_uop_debug_tsrc : _slots_11_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_10_io_valid),
    .io_will_be_valid               (_slots_10_io_will_be_valid),
    .io_request                     (_slots_10_io_request),
    .io_out_uop_uopc                (_slots_10_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_10_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_10_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_10_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_10_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_10_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_10_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_10_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_10_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_10_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_10_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_10_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_10_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_10_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_10_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_10_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_10_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_10_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_10_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_10_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_10_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_10_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_10_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_10_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_10_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_10_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_10_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_10_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_10_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_10_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_10_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_10_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_10_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_10_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_10_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_10_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_10_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_10_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_10_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_10_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_10_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_10_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_10_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_10_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_10_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_10_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_10_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_10_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_10_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_10_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_10_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_10_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_10_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_10_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_10_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_10_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_10_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_10_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_10_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_10_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_10_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_10_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_10_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_10_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_10_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_10_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_10_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_10_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_10_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_10_io_uop_uopc),
    .io_uop_inst                    (_slots_10_io_uop_inst),
    .io_uop_debug_inst              (_slots_10_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_10_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_10_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_10_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_10_io_uop_fu_code),
    .io_uop_iw_state                (_slots_10_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_10_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_10_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_10_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_10_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_10_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_10_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_10_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_10_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_10_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_10_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_10_io_uop_pc_lob),
    .io_uop_taken                   (_slots_10_io_uop_taken),
    .io_uop_imm_packed              (_slots_10_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_10_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_10_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_10_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_10_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_10_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_10_io_uop_pdst),
    .io_uop_prs1                    (_slots_10_io_uop_prs1),
    .io_uop_prs2                    (_slots_10_io_uop_prs2),
    .io_uop_prs3                    (_slots_10_io_uop_prs3),
    .io_uop_ppred                   (_slots_10_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_10_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_10_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_10_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_10_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_10_io_uop_stale_pdst),
    .io_uop_exception               (_slots_10_io_uop_exception),
    .io_uop_exc_cause               (_slots_10_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_10_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_10_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_10_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_10_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_10_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_10_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_10_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_10_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_10_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_10_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_10_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_10_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_10_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_10_io_uop_ldst),
    .io_uop_lrs1                    (_slots_10_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_10_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_10_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_10_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_10_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_10_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_10_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_10_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_10_io_uop_fp_val),
    .io_uop_fp_single               (_slots_10_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_10_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_10_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_10_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_10_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_10_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_10_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_10_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_11 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_11_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_10),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_11_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_31
         ? _slots_14_io_out_uop_uopc
         : _GEN_30 ? _slots_13_io_out_uop_uopc : _slots_12_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_31
         ? _slots_14_io_out_uop_inst
         : _GEN_30 ? _slots_13_io_out_uop_inst : _slots_12_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_31
         ? _slots_14_io_out_uop_debug_inst
         : _GEN_30 ? _slots_13_io_out_uop_debug_inst : _slots_12_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_31
         ? _slots_14_io_out_uop_is_rvc
         : _GEN_30 ? _slots_13_io_out_uop_is_rvc : _slots_12_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_31
         ? _slots_14_io_out_uop_debug_pc
         : _GEN_30 ? _slots_13_io_out_uop_debug_pc : _slots_12_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_31
         ? _slots_14_io_out_uop_iq_type
         : _GEN_30 ? _slots_13_io_out_uop_iq_type : _slots_12_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_31
         ? _slots_14_io_out_uop_fu_code
         : _GEN_30 ? _slots_13_io_out_uop_fu_code : _slots_12_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_31
         ? _slots_14_io_out_uop_iw_state
         : _GEN_30 ? _slots_13_io_out_uop_iw_state : _slots_12_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_31
         ? _slots_14_io_out_uop_iw_p1_poisoned
         : _GEN_30
             ? _slots_13_io_out_uop_iw_p1_poisoned
             : _slots_12_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_31
         ? _slots_14_io_out_uop_iw_p2_poisoned
         : _GEN_30
             ? _slots_13_io_out_uop_iw_p2_poisoned
             : _slots_12_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_31
         ? _slots_14_io_out_uop_is_br
         : _GEN_30 ? _slots_13_io_out_uop_is_br : _slots_12_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_31
         ? _slots_14_io_out_uop_is_jalr
         : _GEN_30 ? _slots_13_io_out_uop_is_jalr : _slots_12_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_31
         ? _slots_14_io_out_uop_is_jal
         : _GEN_30 ? _slots_13_io_out_uop_is_jal : _slots_12_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_31
         ? _slots_14_io_out_uop_is_sfb
         : _GEN_30 ? _slots_13_io_out_uop_is_sfb : _slots_12_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_31
         ? _slots_14_io_out_uop_br_mask
         : _GEN_30 ? _slots_13_io_out_uop_br_mask : _slots_12_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_31
         ? _slots_14_io_out_uop_br_tag
         : _GEN_30 ? _slots_13_io_out_uop_br_tag : _slots_12_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_31
         ? _slots_14_io_out_uop_ftq_idx
         : _GEN_30 ? _slots_13_io_out_uop_ftq_idx : _slots_12_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_31
         ? _slots_14_io_out_uop_edge_inst
         : _GEN_30 ? _slots_13_io_out_uop_edge_inst : _slots_12_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_31
         ? _slots_14_io_out_uop_pc_lob
         : _GEN_30 ? _slots_13_io_out_uop_pc_lob : _slots_12_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_31
         ? _slots_14_io_out_uop_taken
         : _GEN_30 ? _slots_13_io_out_uop_taken : _slots_12_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_31
         ? _slots_14_io_out_uop_imm_packed
         : _GEN_30 ? _slots_13_io_out_uop_imm_packed : _slots_12_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_31
         ? _slots_14_io_out_uop_csr_addr
         : _GEN_30 ? _slots_13_io_out_uop_csr_addr : _slots_12_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_31
         ? _slots_14_io_out_uop_rob_idx
         : _GEN_30 ? _slots_13_io_out_uop_rob_idx : _slots_12_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_31
         ? _slots_14_io_out_uop_ldq_idx
         : _GEN_30 ? _slots_13_io_out_uop_ldq_idx : _slots_12_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_31
         ? _slots_14_io_out_uop_stq_idx
         : _GEN_30 ? _slots_13_io_out_uop_stq_idx : _slots_12_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_31
         ? _slots_14_io_out_uop_rxq_idx
         : _GEN_30 ? _slots_13_io_out_uop_rxq_idx : _slots_12_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_31
         ? _slots_14_io_out_uop_pdst
         : _GEN_30 ? _slots_13_io_out_uop_pdst : _slots_12_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_31
         ? _slots_14_io_out_uop_prs1
         : _GEN_30 ? _slots_13_io_out_uop_prs1 : _slots_12_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_31
         ? _slots_14_io_out_uop_prs2
         : _GEN_30 ? _slots_13_io_out_uop_prs2 : _slots_12_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_31
         ? _slots_14_io_out_uop_prs3
         : _GEN_30 ? _slots_13_io_out_uop_prs3 : _slots_12_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_31
         ? _slots_14_io_out_uop_ppred
         : _GEN_30 ? _slots_13_io_out_uop_ppred : _slots_12_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_31
         ? _slots_14_io_out_uop_prs1_busy
         : _GEN_30 ? _slots_13_io_out_uop_prs1_busy : _slots_12_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_31
         ? _slots_14_io_out_uop_prs2_busy
         : _GEN_30 ? _slots_13_io_out_uop_prs2_busy : _slots_12_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_31
         ? _slots_14_io_out_uop_prs3_busy
         : _GEN_30 ? _slots_13_io_out_uop_prs3_busy : _slots_12_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_31
         ? _slots_14_io_out_uop_ppred_busy
         : _GEN_30 ? _slots_13_io_out_uop_ppred_busy : _slots_12_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_31
         ? _slots_14_io_out_uop_stale_pdst
         : _GEN_30 ? _slots_13_io_out_uop_stale_pdst : _slots_12_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_31
         ? _slots_14_io_out_uop_exception
         : _GEN_30 ? _slots_13_io_out_uop_exception : _slots_12_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_31
         ? _slots_14_io_out_uop_exc_cause
         : _GEN_30 ? _slots_13_io_out_uop_exc_cause : _slots_12_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_31
         ? _slots_14_io_out_uop_bypassable
         : _GEN_30 ? _slots_13_io_out_uop_bypassable : _slots_12_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_31
         ? _slots_14_io_out_uop_mem_cmd
         : _GEN_30 ? _slots_13_io_out_uop_mem_cmd : _slots_12_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_31
         ? _slots_14_io_out_uop_mem_size
         : _GEN_30 ? _slots_13_io_out_uop_mem_size : _slots_12_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_31
         ? _slots_14_io_out_uop_mem_signed
         : _GEN_30 ? _slots_13_io_out_uop_mem_signed : _slots_12_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_31
         ? _slots_14_io_out_uop_is_fence
         : _GEN_30 ? _slots_13_io_out_uop_is_fence : _slots_12_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_31
         ? _slots_14_io_out_uop_is_fencei
         : _GEN_30 ? _slots_13_io_out_uop_is_fencei : _slots_12_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_31
         ? _slots_14_io_out_uop_is_amo
         : _GEN_30 ? _slots_13_io_out_uop_is_amo : _slots_12_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_31
         ? _slots_14_io_out_uop_uses_ldq
         : _GEN_30 ? _slots_13_io_out_uop_uses_ldq : _slots_12_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_31
         ? _slots_14_io_out_uop_uses_stq
         : _GEN_30 ? _slots_13_io_out_uop_uses_stq : _slots_12_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_31
         ? _slots_14_io_out_uop_is_sys_pc2epc
         : _GEN_30
             ? _slots_13_io_out_uop_is_sys_pc2epc
             : _slots_12_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_31
         ? _slots_14_io_out_uop_is_unique
         : _GEN_30 ? _slots_13_io_out_uop_is_unique : _slots_12_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_31
         ? _slots_14_io_out_uop_flush_on_commit
         : _GEN_30
             ? _slots_13_io_out_uop_flush_on_commit
             : _slots_12_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_31
         ? _slots_14_io_out_uop_ldst_is_rs1
         : _GEN_30 ? _slots_13_io_out_uop_ldst_is_rs1 : _slots_12_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_31
         ? _slots_14_io_out_uop_ldst
         : _GEN_30 ? _slots_13_io_out_uop_ldst : _slots_12_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_31
         ? _slots_14_io_out_uop_lrs1
         : _GEN_30 ? _slots_13_io_out_uop_lrs1 : _slots_12_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_31
         ? _slots_14_io_out_uop_lrs2
         : _GEN_30 ? _slots_13_io_out_uop_lrs2 : _slots_12_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_31
         ? _slots_14_io_out_uop_lrs3
         : _GEN_30 ? _slots_13_io_out_uop_lrs3 : _slots_12_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_31
         ? _slots_14_io_out_uop_ldst_val
         : _GEN_30 ? _slots_13_io_out_uop_ldst_val : _slots_12_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_31
         ? _slots_14_io_out_uop_dst_rtype
         : _GEN_30 ? _slots_13_io_out_uop_dst_rtype : _slots_12_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_31
         ? _slots_14_io_out_uop_lrs1_rtype
         : _GEN_30 ? _slots_13_io_out_uop_lrs1_rtype : _slots_12_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_31
         ? _slots_14_io_out_uop_lrs2_rtype
         : _GEN_30 ? _slots_13_io_out_uop_lrs2_rtype : _slots_12_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_31
         ? _slots_14_io_out_uop_frs3_en
         : _GEN_30 ? _slots_13_io_out_uop_frs3_en : _slots_12_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_31
         ? _slots_14_io_out_uop_fp_val
         : _GEN_30 ? _slots_13_io_out_uop_fp_val : _slots_12_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_31
         ? _slots_14_io_out_uop_fp_single
         : _GEN_30 ? _slots_13_io_out_uop_fp_single : _slots_12_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_31
         ? _slots_14_io_out_uop_xcpt_pf_if
         : _GEN_30 ? _slots_13_io_out_uop_xcpt_pf_if : _slots_12_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_31
         ? _slots_14_io_out_uop_xcpt_ae_if
         : _GEN_30 ? _slots_13_io_out_uop_xcpt_ae_if : _slots_12_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_31
         ? _slots_14_io_out_uop_xcpt_ma_if
         : _GEN_30 ? _slots_13_io_out_uop_xcpt_ma_if : _slots_12_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_31
         ? _slots_14_io_out_uop_bp_debug_if
         : _GEN_30 ? _slots_13_io_out_uop_bp_debug_if : _slots_12_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_31
         ? _slots_14_io_out_uop_bp_xcpt_if
         : _GEN_30 ? _slots_13_io_out_uop_bp_xcpt_if : _slots_12_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_31
         ? _slots_14_io_out_uop_debug_fsrc
         : _GEN_30 ? _slots_13_io_out_uop_debug_fsrc : _slots_12_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_31
         ? _slots_14_io_out_uop_debug_tsrc
         : _GEN_30 ? _slots_13_io_out_uop_debug_tsrc : _slots_12_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_11_io_valid),
    .io_will_be_valid               (_slots_11_io_will_be_valid),
    .io_request                     (_slots_11_io_request),
    .io_out_uop_uopc                (_slots_11_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_11_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_11_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_11_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_11_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_11_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_11_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_11_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_11_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_11_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_11_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_11_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_11_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_11_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_11_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_11_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_11_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_11_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_11_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_11_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_11_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_11_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_11_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_11_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_11_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_11_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_11_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_11_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_11_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_11_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_11_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_11_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_11_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_11_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_11_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_11_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_11_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_11_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_11_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_11_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_11_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_11_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_11_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_11_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_11_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_11_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_11_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_11_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_11_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_11_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_11_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_11_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_11_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_11_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_11_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_11_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_11_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_11_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_11_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_11_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_11_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_11_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_11_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_11_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_11_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_11_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_11_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_11_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_11_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_11_io_uop_uopc),
    .io_uop_inst                    (_slots_11_io_uop_inst),
    .io_uop_debug_inst              (_slots_11_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_11_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_11_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_11_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_11_io_uop_fu_code),
    .io_uop_iw_state                (_slots_11_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_11_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_11_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_11_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_11_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_11_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_11_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_11_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_11_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_11_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_11_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_11_io_uop_pc_lob),
    .io_uop_taken                   (_slots_11_io_uop_taken),
    .io_uop_imm_packed              (_slots_11_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_11_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_11_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_11_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_11_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_11_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_11_io_uop_pdst),
    .io_uop_prs1                    (_slots_11_io_uop_prs1),
    .io_uop_prs2                    (_slots_11_io_uop_prs2),
    .io_uop_prs3                    (_slots_11_io_uop_prs3),
    .io_uop_ppred                   (_slots_11_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_11_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_11_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_11_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_11_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_11_io_uop_stale_pdst),
    .io_uop_exception               (_slots_11_io_uop_exception),
    .io_uop_exc_cause               (_slots_11_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_11_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_11_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_11_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_11_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_11_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_11_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_11_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_11_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_11_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_11_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_11_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_11_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_11_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_11_io_uop_ldst),
    .io_uop_lrs1                    (_slots_11_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_11_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_11_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_11_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_11_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_11_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_11_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_11_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_11_io_uop_fp_val),
    .io_uop_fp_single               (_slots_11_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_11_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_11_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_11_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_11_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_11_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_11_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_11_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_12 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_12_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_11),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_12_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_33
         ? _slots_15_io_out_uop_uopc
         : _GEN_32 ? _slots_14_io_out_uop_uopc : _slots_13_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_33
         ? _slots_15_io_out_uop_inst
         : _GEN_32 ? _slots_14_io_out_uop_inst : _slots_13_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_33
         ? _slots_15_io_out_uop_debug_inst
         : _GEN_32 ? _slots_14_io_out_uop_debug_inst : _slots_13_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_33
         ? _slots_15_io_out_uop_is_rvc
         : _GEN_32 ? _slots_14_io_out_uop_is_rvc : _slots_13_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_33
         ? _slots_15_io_out_uop_debug_pc
         : _GEN_32 ? _slots_14_io_out_uop_debug_pc : _slots_13_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_33
         ? _slots_15_io_out_uop_iq_type
         : _GEN_32 ? _slots_14_io_out_uop_iq_type : _slots_13_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_33
         ? _slots_15_io_out_uop_fu_code
         : _GEN_32 ? _slots_14_io_out_uop_fu_code : _slots_13_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_33
         ? _slots_15_io_out_uop_iw_state
         : _GEN_32 ? _slots_14_io_out_uop_iw_state : _slots_13_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_33
         ? _slots_15_io_out_uop_iw_p1_poisoned
         : _GEN_32
             ? _slots_14_io_out_uop_iw_p1_poisoned
             : _slots_13_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_33
         ? _slots_15_io_out_uop_iw_p2_poisoned
         : _GEN_32
             ? _slots_14_io_out_uop_iw_p2_poisoned
             : _slots_13_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_33
         ? _slots_15_io_out_uop_is_br
         : _GEN_32 ? _slots_14_io_out_uop_is_br : _slots_13_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_33
         ? _slots_15_io_out_uop_is_jalr
         : _GEN_32 ? _slots_14_io_out_uop_is_jalr : _slots_13_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_33
         ? _slots_15_io_out_uop_is_jal
         : _GEN_32 ? _slots_14_io_out_uop_is_jal : _slots_13_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_33
         ? _slots_15_io_out_uop_is_sfb
         : _GEN_32 ? _slots_14_io_out_uop_is_sfb : _slots_13_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_33
         ? _slots_15_io_out_uop_br_mask
         : _GEN_32 ? _slots_14_io_out_uop_br_mask : _slots_13_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_33
         ? _slots_15_io_out_uop_br_tag
         : _GEN_32 ? _slots_14_io_out_uop_br_tag : _slots_13_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_33
         ? _slots_15_io_out_uop_ftq_idx
         : _GEN_32 ? _slots_14_io_out_uop_ftq_idx : _slots_13_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_33
         ? _slots_15_io_out_uop_edge_inst
         : _GEN_32 ? _slots_14_io_out_uop_edge_inst : _slots_13_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_33
         ? _slots_15_io_out_uop_pc_lob
         : _GEN_32 ? _slots_14_io_out_uop_pc_lob : _slots_13_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_33
         ? _slots_15_io_out_uop_taken
         : _GEN_32 ? _slots_14_io_out_uop_taken : _slots_13_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_33
         ? _slots_15_io_out_uop_imm_packed
         : _GEN_32 ? _slots_14_io_out_uop_imm_packed : _slots_13_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_33
         ? _slots_15_io_out_uop_csr_addr
         : _GEN_32 ? _slots_14_io_out_uop_csr_addr : _slots_13_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_33
         ? _slots_15_io_out_uop_rob_idx
         : _GEN_32 ? _slots_14_io_out_uop_rob_idx : _slots_13_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_33
         ? _slots_15_io_out_uop_ldq_idx
         : _GEN_32 ? _slots_14_io_out_uop_ldq_idx : _slots_13_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_33
         ? _slots_15_io_out_uop_stq_idx
         : _GEN_32 ? _slots_14_io_out_uop_stq_idx : _slots_13_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_33
         ? _slots_15_io_out_uop_rxq_idx
         : _GEN_32 ? _slots_14_io_out_uop_rxq_idx : _slots_13_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_33
         ? _slots_15_io_out_uop_pdst
         : _GEN_32 ? _slots_14_io_out_uop_pdst : _slots_13_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_33
         ? _slots_15_io_out_uop_prs1
         : _GEN_32 ? _slots_14_io_out_uop_prs1 : _slots_13_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_33
         ? _slots_15_io_out_uop_prs2
         : _GEN_32 ? _slots_14_io_out_uop_prs2 : _slots_13_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_33
         ? _slots_15_io_out_uop_prs3
         : _GEN_32 ? _slots_14_io_out_uop_prs3 : _slots_13_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_33
         ? _slots_15_io_out_uop_ppred
         : _GEN_32 ? _slots_14_io_out_uop_ppred : _slots_13_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_33
         ? _slots_15_io_out_uop_prs1_busy
         : _GEN_32 ? _slots_14_io_out_uop_prs1_busy : _slots_13_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_33
         ? _slots_15_io_out_uop_prs2_busy
         : _GEN_32 ? _slots_14_io_out_uop_prs2_busy : _slots_13_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_33
         ? _slots_15_io_out_uop_prs3_busy
         : _GEN_32 ? _slots_14_io_out_uop_prs3_busy : _slots_13_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_33
         ? _slots_15_io_out_uop_ppred_busy
         : _GEN_32 ? _slots_14_io_out_uop_ppred_busy : _slots_13_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_33
         ? _slots_15_io_out_uop_stale_pdst
         : _GEN_32 ? _slots_14_io_out_uop_stale_pdst : _slots_13_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_33
         ? _slots_15_io_out_uop_exception
         : _GEN_32 ? _slots_14_io_out_uop_exception : _slots_13_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_33
         ? _slots_15_io_out_uop_exc_cause
         : _GEN_32 ? _slots_14_io_out_uop_exc_cause : _slots_13_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_33
         ? _slots_15_io_out_uop_bypassable
         : _GEN_32 ? _slots_14_io_out_uop_bypassable : _slots_13_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_33
         ? _slots_15_io_out_uop_mem_cmd
         : _GEN_32 ? _slots_14_io_out_uop_mem_cmd : _slots_13_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_33
         ? _slots_15_io_out_uop_mem_size
         : _GEN_32 ? _slots_14_io_out_uop_mem_size : _slots_13_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_33
         ? _slots_15_io_out_uop_mem_signed
         : _GEN_32 ? _slots_14_io_out_uop_mem_signed : _slots_13_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_33
         ? _slots_15_io_out_uop_is_fence
         : _GEN_32 ? _slots_14_io_out_uop_is_fence : _slots_13_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_33
         ? _slots_15_io_out_uop_is_fencei
         : _GEN_32 ? _slots_14_io_out_uop_is_fencei : _slots_13_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_33
         ? _slots_15_io_out_uop_is_amo
         : _GEN_32 ? _slots_14_io_out_uop_is_amo : _slots_13_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_33
         ? _slots_15_io_out_uop_uses_ldq
         : _GEN_32 ? _slots_14_io_out_uop_uses_ldq : _slots_13_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_33
         ? _slots_15_io_out_uop_uses_stq
         : _GEN_32 ? _slots_14_io_out_uop_uses_stq : _slots_13_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_33
         ? _slots_15_io_out_uop_is_sys_pc2epc
         : _GEN_32
             ? _slots_14_io_out_uop_is_sys_pc2epc
             : _slots_13_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_33
         ? _slots_15_io_out_uop_is_unique
         : _GEN_32 ? _slots_14_io_out_uop_is_unique : _slots_13_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_33
         ? _slots_15_io_out_uop_flush_on_commit
         : _GEN_32
             ? _slots_14_io_out_uop_flush_on_commit
             : _slots_13_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_33
         ? _slots_15_io_out_uop_ldst_is_rs1
         : _GEN_32 ? _slots_14_io_out_uop_ldst_is_rs1 : _slots_13_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_33
         ? _slots_15_io_out_uop_ldst
         : _GEN_32 ? _slots_14_io_out_uop_ldst : _slots_13_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_33
         ? _slots_15_io_out_uop_lrs1
         : _GEN_32 ? _slots_14_io_out_uop_lrs1 : _slots_13_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_33
         ? _slots_15_io_out_uop_lrs2
         : _GEN_32 ? _slots_14_io_out_uop_lrs2 : _slots_13_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_33
         ? _slots_15_io_out_uop_lrs3
         : _GEN_32 ? _slots_14_io_out_uop_lrs3 : _slots_13_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_33
         ? _slots_15_io_out_uop_ldst_val
         : _GEN_32 ? _slots_14_io_out_uop_ldst_val : _slots_13_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_33
         ? _slots_15_io_out_uop_dst_rtype
         : _GEN_32 ? _slots_14_io_out_uop_dst_rtype : _slots_13_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_33
         ? _slots_15_io_out_uop_lrs1_rtype
         : _GEN_32 ? _slots_14_io_out_uop_lrs1_rtype : _slots_13_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_33
         ? _slots_15_io_out_uop_lrs2_rtype
         : _GEN_32 ? _slots_14_io_out_uop_lrs2_rtype : _slots_13_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_33
         ? _slots_15_io_out_uop_frs3_en
         : _GEN_32 ? _slots_14_io_out_uop_frs3_en : _slots_13_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_33
         ? _slots_15_io_out_uop_fp_val
         : _GEN_32 ? _slots_14_io_out_uop_fp_val : _slots_13_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_33
         ? _slots_15_io_out_uop_fp_single
         : _GEN_32 ? _slots_14_io_out_uop_fp_single : _slots_13_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_33
         ? _slots_15_io_out_uop_xcpt_pf_if
         : _GEN_32 ? _slots_14_io_out_uop_xcpt_pf_if : _slots_13_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_33
         ? _slots_15_io_out_uop_xcpt_ae_if
         : _GEN_32 ? _slots_14_io_out_uop_xcpt_ae_if : _slots_13_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_33
         ? _slots_15_io_out_uop_xcpt_ma_if
         : _GEN_32 ? _slots_14_io_out_uop_xcpt_ma_if : _slots_13_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_33
         ? _slots_15_io_out_uop_bp_debug_if
         : _GEN_32 ? _slots_14_io_out_uop_bp_debug_if : _slots_13_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_33
         ? _slots_15_io_out_uop_bp_xcpt_if
         : _GEN_32 ? _slots_14_io_out_uop_bp_xcpt_if : _slots_13_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_33
         ? _slots_15_io_out_uop_debug_fsrc
         : _GEN_32 ? _slots_14_io_out_uop_debug_fsrc : _slots_13_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_33
         ? _slots_15_io_out_uop_debug_tsrc
         : _GEN_32 ? _slots_14_io_out_uop_debug_tsrc : _slots_13_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_12_io_valid),
    .io_will_be_valid               (_slots_12_io_will_be_valid),
    .io_request                     (_slots_12_io_request),
    .io_out_uop_uopc                (_slots_12_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_12_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_12_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_12_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_12_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_12_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_12_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_12_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_12_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_12_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_12_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_12_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_12_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_12_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_12_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_12_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_12_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_12_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_12_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_12_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_12_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_12_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_12_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_12_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_12_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_12_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_12_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_12_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_12_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_12_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_12_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_12_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_12_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_12_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_12_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_12_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_12_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_12_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_12_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_12_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_12_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_12_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_12_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_12_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_12_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_12_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_12_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_12_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_12_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_12_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_12_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_12_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_12_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_12_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_12_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_12_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_12_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_12_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_12_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_12_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_12_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_12_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_12_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_12_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_12_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_12_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_12_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_12_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_12_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_12_io_uop_uopc),
    .io_uop_inst                    (_slots_12_io_uop_inst),
    .io_uop_debug_inst              (_slots_12_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_12_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_12_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_12_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_12_io_uop_fu_code),
    .io_uop_iw_state                (_slots_12_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_12_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_12_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_12_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_12_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_12_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_12_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_12_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_12_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_12_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_12_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_12_io_uop_pc_lob),
    .io_uop_taken                   (_slots_12_io_uop_taken),
    .io_uop_imm_packed              (_slots_12_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_12_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_12_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_12_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_12_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_12_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_12_io_uop_pdst),
    .io_uop_prs1                    (_slots_12_io_uop_prs1),
    .io_uop_prs2                    (_slots_12_io_uop_prs2),
    .io_uop_prs3                    (_slots_12_io_uop_prs3),
    .io_uop_ppred                   (_slots_12_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_12_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_12_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_12_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_12_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_12_io_uop_stale_pdst),
    .io_uop_exception               (_slots_12_io_uop_exception),
    .io_uop_exc_cause               (_slots_12_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_12_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_12_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_12_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_12_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_12_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_12_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_12_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_12_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_12_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_12_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_12_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_12_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_12_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_12_io_uop_ldst),
    .io_uop_lrs1                    (_slots_12_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_12_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_12_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_12_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_12_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_12_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_12_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_12_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_12_io_uop_fp_val),
    .io_uop_fp_single               (_slots_12_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_12_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_12_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_12_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_12_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_12_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_12_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_12_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_13 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_13_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_12),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_13_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_35
         ? _slots_16_io_out_uop_uopc
         : _GEN_34 ? _slots_15_io_out_uop_uopc : _slots_14_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_35
         ? _slots_16_io_out_uop_inst
         : _GEN_34 ? _slots_15_io_out_uop_inst : _slots_14_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_35
         ? _slots_16_io_out_uop_debug_inst
         : _GEN_34 ? _slots_15_io_out_uop_debug_inst : _slots_14_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_35
         ? _slots_16_io_out_uop_is_rvc
         : _GEN_34 ? _slots_15_io_out_uop_is_rvc : _slots_14_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_35
         ? _slots_16_io_out_uop_debug_pc
         : _GEN_34 ? _slots_15_io_out_uop_debug_pc : _slots_14_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_35
         ? _slots_16_io_out_uop_iq_type
         : _GEN_34 ? _slots_15_io_out_uop_iq_type : _slots_14_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_35
         ? _slots_16_io_out_uop_fu_code
         : _GEN_34 ? _slots_15_io_out_uop_fu_code : _slots_14_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_35
         ? _slots_16_io_out_uop_iw_state
         : _GEN_34 ? _slots_15_io_out_uop_iw_state : _slots_14_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_35
         ? _slots_16_io_out_uop_iw_p1_poisoned
         : _GEN_34
             ? _slots_15_io_out_uop_iw_p1_poisoned
             : _slots_14_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_35
         ? _slots_16_io_out_uop_iw_p2_poisoned
         : _GEN_34
             ? _slots_15_io_out_uop_iw_p2_poisoned
             : _slots_14_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_35
         ? _slots_16_io_out_uop_is_br
         : _GEN_34 ? _slots_15_io_out_uop_is_br : _slots_14_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_35
         ? _slots_16_io_out_uop_is_jalr
         : _GEN_34 ? _slots_15_io_out_uop_is_jalr : _slots_14_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_35
         ? _slots_16_io_out_uop_is_jal
         : _GEN_34 ? _slots_15_io_out_uop_is_jal : _slots_14_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_35
         ? _slots_16_io_out_uop_is_sfb
         : _GEN_34 ? _slots_15_io_out_uop_is_sfb : _slots_14_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_35
         ? _slots_16_io_out_uop_br_mask
         : _GEN_34 ? _slots_15_io_out_uop_br_mask : _slots_14_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_35
         ? _slots_16_io_out_uop_br_tag
         : _GEN_34 ? _slots_15_io_out_uop_br_tag : _slots_14_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_35
         ? _slots_16_io_out_uop_ftq_idx
         : _GEN_34 ? _slots_15_io_out_uop_ftq_idx : _slots_14_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_35
         ? _slots_16_io_out_uop_edge_inst
         : _GEN_34 ? _slots_15_io_out_uop_edge_inst : _slots_14_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_35
         ? _slots_16_io_out_uop_pc_lob
         : _GEN_34 ? _slots_15_io_out_uop_pc_lob : _slots_14_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_35
         ? _slots_16_io_out_uop_taken
         : _GEN_34 ? _slots_15_io_out_uop_taken : _slots_14_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_35
         ? _slots_16_io_out_uop_imm_packed
         : _GEN_34 ? _slots_15_io_out_uop_imm_packed : _slots_14_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_35
         ? _slots_16_io_out_uop_csr_addr
         : _GEN_34 ? _slots_15_io_out_uop_csr_addr : _slots_14_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_35
         ? _slots_16_io_out_uop_rob_idx
         : _GEN_34 ? _slots_15_io_out_uop_rob_idx : _slots_14_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_35
         ? _slots_16_io_out_uop_ldq_idx
         : _GEN_34 ? _slots_15_io_out_uop_ldq_idx : _slots_14_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_35
         ? _slots_16_io_out_uop_stq_idx
         : _GEN_34 ? _slots_15_io_out_uop_stq_idx : _slots_14_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_35
         ? _slots_16_io_out_uop_rxq_idx
         : _GEN_34 ? _slots_15_io_out_uop_rxq_idx : _slots_14_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_35
         ? _slots_16_io_out_uop_pdst
         : _GEN_34 ? _slots_15_io_out_uop_pdst : _slots_14_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_35
         ? _slots_16_io_out_uop_prs1
         : _GEN_34 ? _slots_15_io_out_uop_prs1 : _slots_14_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_35
         ? _slots_16_io_out_uop_prs2
         : _GEN_34 ? _slots_15_io_out_uop_prs2 : _slots_14_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_35
         ? _slots_16_io_out_uop_prs3
         : _GEN_34 ? _slots_15_io_out_uop_prs3 : _slots_14_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_35
         ? _slots_16_io_out_uop_ppred
         : _GEN_34 ? _slots_15_io_out_uop_ppred : _slots_14_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_35
         ? _slots_16_io_out_uop_prs1_busy
         : _GEN_34 ? _slots_15_io_out_uop_prs1_busy : _slots_14_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_35
         ? _slots_16_io_out_uop_prs2_busy
         : _GEN_34 ? _slots_15_io_out_uop_prs2_busy : _slots_14_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_35
         ? _slots_16_io_out_uop_prs3_busy
         : _GEN_34 ? _slots_15_io_out_uop_prs3_busy : _slots_14_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_35
         ? _slots_16_io_out_uop_ppred_busy
         : _GEN_34 ? _slots_15_io_out_uop_ppred_busy : _slots_14_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_35
         ? _slots_16_io_out_uop_stale_pdst
         : _GEN_34 ? _slots_15_io_out_uop_stale_pdst : _slots_14_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_35
         ? _slots_16_io_out_uop_exception
         : _GEN_34 ? _slots_15_io_out_uop_exception : _slots_14_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_35
         ? _slots_16_io_out_uop_exc_cause
         : _GEN_34 ? _slots_15_io_out_uop_exc_cause : _slots_14_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_35
         ? _slots_16_io_out_uop_bypassable
         : _GEN_34 ? _slots_15_io_out_uop_bypassable : _slots_14_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_35
         ? _slots_16_io_out_uop_mem_cmd
         : _GEN_34 ? _slots_15_io_out_uop_mem_cmd : _slots_14_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_35
         ? _slots_16_io_out_uop_mem_size
         : _GEN_34 ? _slots_15_io_out_uop_mem_size : _slots_14_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_35
         ? _slots_16_io_out_uop_mem_signed
         : _GEN_34 ? _slots_15_io_out_uop_mem_signed : _slots_14_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_35
         ? _slots_16_io_out_uop_is_fence
         : _GEN_34 ? _slots_15_io_out_uop_is_fence : _slots_14_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_35
         ? _slots_16_io_out_uop_is_fencei
         : _GEN_34 ? _slots_15_io_out_uop_is_fencei : _slots_14_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_35
         ? _slots_16_io_out_uop_is_amo
         : _GEN_34 ? _slots_15_io_out_uop_is_amo : _slots_14_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_35
         ? _slots_16_io_out_uop_uses_ldq
         : _GEN_34 ? _slots_15_io_out_uop_uses_ldq : _slots_14_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_35
         ? _slots_16_io_out_uop_uses_stq
         : _GEN_34 ? _slots_15_io_out_uop_uses_stq : _slots_14_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_35
         ? _slots_16_io_out_uop_is_sys_pc2epc
         : _GEN_34
             ? _slots_15_io_out_uop_is_sys_pc2epc
             : _slots_14_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_35
         ? _slots_16_io_out_uop_is_unique
         : _GEN_34 ? _slots_15_io_out_uop_is_unique : _slots_14_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_35
         ? _slots_16_io_out_uop_flush_on_commit
         : _GEN_34
             ? _slots_15_io_out_uop_flush_on_commit
             : _slots_14_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_35
         ? _slots_16_io_out_uop_ldst_is_rs1
         : _GEN_34 ? _slots_15_io_out_uop_ldst_is_rs1 : _slots_14_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_35
         ? _slots_16_io_out_uop_ldst
         : _GEN_34 ? _slots_15_io_out_uop_ldst : _slots_14_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_35
         ? _slots_16_io_out_uop_lrs1
         : _GEN_34 ? _slots_15_io_out_uop_lrs1 : _slots_14_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_35
         ? _slots_16_io_out_uop_lrs2
         : _GEN_34 ? _slots_15_io_out_uop_lrs2 : _slots_14_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_35
         ? _slots_16_io_out_uop_lrs3
         : _GEN_34 ? _slots_15_io_out_uop_lrs3 : _slots_14_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_35
         ? _slots_16_io_out_uop_ldst_val
         : _GEN_34 ? _slots_15_io_out_uop_ldst_val : _slots_14_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_35
         ? _slots_16_io_out_uop_dst_rtype
         : _GEN_34 ? _slots_15_io_out_uop_dst_rtype : _slots_14_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_35
         ? _slots_16_io_out_uop_lrs1_rtype
         : _GEN_34 ? _slots_15_io_out_uop_lrs1_rtype : _slots_14_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_35
         ? _slots_16_io_out_uop_lrs2_rtype
         : _GEN_34 ? _slots_15_io_out_uop_lrs2_rtype : _slots_14_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_35
         ? _slots_16_io_out_uop_frs3_en
         : _GEN_34 ? _slots_15_io_out_uop_frs3_en : _slots_14_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_35
         ? _slots_16_io_out_uop_fp_val
         : _GEN_34 ? _slots_15_io_out_uop_fp_val : _slots_14_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_35
         ? _slots_16_io_out_uop_fp_single
         : _GEN_34 ? _slots_15_io_out_uop_fp_single : _slots_14_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_35
         ? _slots_16_io_out_uop_xcpt_pf_if
         : _GEN_34 ? _slots_15_io_out_uop_xcpt_pf_if : _slots_14_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_35
         ? _slots_16_io_out_uop_xcpt_ae_if
         : _GEN_34 ? _slots_15_io_out_uop_xcpt_ae_if : _slots_14_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_35
         ? _slots_16_io_out_uop_xcpt_ma_if
         : _GEN_34 ? _slots_15_io_out_uop_xcpt_ma_if : _slots_14_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_35
         ? _slots_16_io_out_uop_bp_debug_if
         : _GEN_34 ? _slots_15_io_out_uop_bp_debug_if : _slots_14_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_35
         ? _slots_16_io_out_uop_bp_xcpt_if
         : _GEN_34 ? _slots_15_io_out_uop_bp_xcpt_if : _slots_14_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_35
         ? _slots_16_io_out_uop_debug_fsrc
         : _GEN_34 ? _slots_15_io_out_uop_debug_fsrc : _slots_14_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_35
         ? _slots_16_io_out_uop_debug_tsrc
         : _GEN_34 ? _slots_15_io_out_uop_debug_tsrc : _slots_14_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_13_io_valid),
    .io_will_be_valid               (_slots_13_io_will_be_valid),
    .io_request                     (_slots_13_io_request),
    .io_out_uop_uopc                (_slots_13_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_13_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_13_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_13_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_13_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_13_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_13_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_13_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_13_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_13_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_13_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_13_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_13_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_13_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_13_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_13_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_13_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_13_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_13_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_13_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_13_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_13_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_13_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_13_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_13_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_13_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_13_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_13_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_13_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_13_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_13_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_13_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_13_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_13_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_13_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_13_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_13_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_13_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_13_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_13_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_13_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_13_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_13_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_13_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_13_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_13_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_13_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_13_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_13_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_13_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_13_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_13_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_13_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_13_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_13_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_13_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_13_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_13_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_13_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_13_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_13_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_13_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_13_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_13_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_13_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_13_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_13_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_13_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_13_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_13_io_uop_uopc),
    .io_uop_inst                    (_slots_13_io_uop_inst),
    .io_uop_debug_inst              (_slots_13_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_13_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_13_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_13_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_13_io_uop_fu_code),
    .io_uop_iw_state                (_slots_13_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_13_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_13_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_13_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_13_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_13_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_13_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_13_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_13_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_13_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_13_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_13_io_uop_pc_lob),
    .io_uop_taken                   (_slots_13_io_uop_taken),
    .io_uop_imm_packed              (_slots_13_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_13_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_13_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_13_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_13_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_13_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_13_io_uop_pdst),
    .io_uop_prs1                    (_slots_13_io_uop_prs1),
    .io_uop_prs2                    (_slots_13_io_uop_prs2),
    .io_uop_prs3                    (_slots_13_io_uop_prs3),
    .io_uop_ppred                   (_slots_13_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_13_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_13_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_13_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_13_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_13_io_uop_stale_pdst),
    .io_uop_exception               (_slots_13_io_uop_exception),
    .io_uop_exc_cause               (_slots_13_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_13_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_13_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_13_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_13_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_13_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_13_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_13_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_13_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_13_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_13_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_13_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_13_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_13_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_13_io_uop_ldst),
    .io_uop_lrs1                    (_slots_13_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_13_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_13_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_13_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_13_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_13_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_13_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_13_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_13_io_uop_fp_val),
    .io_uop_fp_single               (_slots_13_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_13_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_13_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_13_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_13_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_13_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_13_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_13_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_14 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_14_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_13),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_14_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_37
         ? _slots_17_io_out_uop_uopc
         : _GEN_36 ? _slots_16_io_out_uop_uopc : _slots_15_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_37
         ? _slots_17_io_out_uop_inst
         : _GEN_36 ? _slots_16_io_out_uop_inst : _slots_15_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_37
         ? _slots_17_io_out_uop_debug_inst
         : _GEN_36 ? _slots_16_io_out_uop_debug_inst : _slots_15_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_37
         ? _slots_17_io_out_uop_is_rvc
         : _GEN_36 ? _slots_16_io_out_uop_is_rvc : _slots_15_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_37
         ? _slots_17_io_out_uop_debug_pc
         : _GEN_36 ? _slots_16_io_out_uop_debug_pc : _slots_15_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_37
         ? _slots_17_io_out_uop_iq_type
         : _GEN_36 ? _slots_16_io_out_uop_iq_type : _slots_15_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_37
         ? _slots_17_io_out_uop_fu_code
         : _GEN_36 ? _slots_16_io_out_uop_fu_code : _slots_15_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_37
         ? _slots_17_io_out_uop_iw_state
         : _GEN_36 ? _slots_16_io_out_uop_iw_state : _slots_15_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_37
         ? _slots_17_io_out_uop_iw_p1_poisoned
         : _GEN_36
             ? _slots_16_io_out_uop_iw_p1_poisoned
             : _slots_15_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_37
         ? _slots_17_io_out_uop_iw_p2_poisoned
         : _GEN_36
             ? _slots_16_io_out_uop_iw_p2_poisoned
             : _slots_15_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_37
         ? _slots_17_io_out_uop_is_br
         : _GEN_36 ? _slots_16_io_out_uop_is_br : _slots_15_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_37
         ? _slots_17_io_out_uop_is_jalr
         : _GEN_36 ? _slots_16_io_out_uop_is_jalr : _slots_15_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_37
         ? _slots_17_io_out_uop_is_jal
         : _GEN_36 ? _slots_16_io_out_uop_is_jal : _slots_15_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_37
         ? _slots_17_io_out_uop_is_sfb
         : _GEN_36 ? _slots_16_io_out_uop_is_sfb : _slots_15_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_37
         ? _slots_17_io_out_uop_br_mask
         : _GEN_36 ? _slots_16_io_out_uop_br_mask : _slots_15_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_37
         ? _slots_17_io_out_uop_br_tag
         : _GEN_36 ? _slots_16_io_out_uop_br_tag : _slots_15_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_37
         ? _slots_17_io_out_uop_ftq_idx
         : _GEN_36 ? _slots_16_io_out_uop_ftq_idx : _slots_15_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_37
         ? _slots_17_io_out_uop_edge_inst
         : _GEN_36 ? _slots_16_io_out_uop_edge_inst : _slots_15_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_37
         ? _slots_17_io_out_uop_pc_lob
         : _GEN_36 ? _slots_16_io_out_uop_pc_lob : _slots_15_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_37
         ? _slots_17_io_out_uop_taken
         : _GEN_36 ? _slots_16_io_out_uop_taken : _slots_15_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_37
         ? _slots_17_io_out_uop_imm_packed
         : _GEN_36 ? _slots_16_io_out_uop_imm_packed : _slots_15_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_37
         ? _slots_17_io_out_uop_csr_addr
         : _GEN_36 ? _slots_16_io_out_uop_csr_addr : _slots_15_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_37
         ? _slots_17_io_out_uop_rob_idx
         : _GEN_36 ? _slots_16_io_out_uop_rob_idx : _slots_15_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_37
         ? _slots_17_io_out_uop_ldq_idx
         : _GEN_36 ? _slots_16_io_out_uop_ldq_idx : _slots_15_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_37
         ? _slots_17_io_out_uop_stq_idx
         : _GEN_36 ? _slots_16_io_out_uop_stq_idx : _slots_15_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_37
         ? _slots_17_io_out_uop_rxq_idx
         : _GEN_36 ? _slots_16_io_out_uop_rxq_idx : _slots_15_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_37
         ? _slots_17_io_out_uop_pdst
         : _GEN_36 ? _slots_16_io_out_uop_pdst : _slots_15_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_37
         ? _slots_17_io_out_uop_prs1
         : _GEN_36 ? _slots_16_io_out_uop_prs1 : _slots_15_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_37
         ? _slots_17_io_out_uop_prs2
         : _GEN_36 ? _slots_16_io_out_uop_prs2 : _slots_15_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_37
         ? _slots_17_io_out_uop_prs3
         : _GEN_36 ? _slots_16_io_out_uop_prs3 : _slots_15_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_37
         ? _slots_17_io_out_uop_ppred
         : _GEN_36 ? _slots_16_io_out_uop_ppred : _slots_15_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_37
         ? _slots_17_io_out_uop_prs1_busy
         : _GEN_36 ? _slots_16_io_out_uop_prs1_busy : _slots_15_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_37
         ? _slots_17_io_out_uop_prs2_busy
         : _GEN_36 ? _slots_16_io_out_uop_prs2_busy : _slots_15_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_37
         ? _slots_17_io_out_uop_prs3_busy
         : _GEN_36 ? _slots_16_io_out_uop_prs3_busy : _slots_15_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_37
         ? _slots_17_io_out_uop_ppred_busy
         : _GEN_36 ? _slots_16_io_out_uop_ppred_busy : _slots_15_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_37
         ? _slots_17_io_out_uop_stale_pdst
         : _GEN_36 ? _slots_16_io_out_uop_stale_pdst : _slots_15_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_37
         ? _slots_17_io_out_uop_exception
         : _GEN_36 ? _slots_16_io_out_uop_exception : _slots_15_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_37
         ? _slots_17_io_out_uop_exc_cause
         : _GEN_36 ? _slots_16_io_out_uop_exc_cause : _slots_15_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_37
         ? _slots_17_io_out_uop_bypassable
         : _GEN_36 ? _slots_16_io_out_uop_bypassable : _slots_15_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_37
         ? _slots_17_io_out_uop_mem_cmd
         : _GEN_36 ? _slots_16_io_out_uop_mem_cmd : _slots_15_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_37
         ? _slots_17_io_out_uop_mem_size
         : _GEN_36 ? _slots_16_io_out_uop_mem_size : _slots_15_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_37
         ? _slots_17_io_out_uop_mem_signed
         : _GEN_36 ? _slots_16_io_out_uop_mem_signed : _slots_15_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_37
         ? _slots_17_io_out_uop_is_fence
         : _GEN_36 ? _slots_16_io_out_uop_is_fence : _slots_15_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_37
         ? _slots_17_io_out_uop_is_fencei
         : _GEN_36 ? _slots_16_io_out_uop_is_fencei : _slots_15_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_37
         ? _slots_17_io_out_uop_is_amo
         : _GEN_36 ? _slots_16_io_out_uop_is_amo : _slots_15_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_37
         ? _slots_17_io_out_uop_uses_ldq
         : _GEN_36 ? _slots_16_io_out_uop_uses_ldq : _slots_15_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_37
         ? _slots_17_io_out_uop_uses_stq
         : _GEN_36 ? _slots_16_io_out_uop_uses_stq : _slots_15_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_37
         ? _slots_17_io_out_uop_is_sys_pc2epc
         : _GEN_36
             ? _slots_16_io_out_uop_is_sys_pc2epc
             : _slots_15_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_37
         ? _slots_17_io_out_uop_is_unique
         : _GEN_36 ? _slots_16_io_out_uop_is_unique : _slots_15_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_37
         ? _slots_17_io_out_uop_flush_on_commit
         : _GEN_36
             ? _slots_16_io_out_uop_flush_on_commit
             : _slots_15_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_37
         ? _slots_17_io_out_uop_ldst_is_rs1
         : _GEN_36 ? _slots_16_io_out_uop_ldst_is_rs1 : _slots_15_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_37
         ? _slots_17_io_out_uop_ldst
         : _GEN_36 ? _slots_16_io_out_uop_ldst : _slots_15_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_37
         ? _slots_17_io_out_uop_lrs1
         : _GEN_36 ? _slots_16_io_out_uop_lrs1 : _slots_15_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_37
         ? _slots_17_io_out_uop_lrs2
         : _GEN_36 ? _slots_16_io_out_uop_lrs2 : _slots_15_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_37
         ? _slots_17_io_out_uop_lrs3
         : _GEN_36 ? _slots_16_io_out_uop_lrs3 : _slots_15_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_37
         ? _slots_17_io_out_uop_ldst_val
         : _GEN_36 ? _slots_16_io_out_uop_ldst_val : _slots_15_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_37
         ? _slots_17_io_out_uop_dst_rtype
         : _GEN_36 ? _slots_16_io_out_uop_dst_rtype : _slots_15_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_37
         ? _slots_17_io_out_uop_lrs1_rtype
         : _GEN_36 ? _slots_16_io_out_uop_lrs1_rtype : _slots_15_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_37
         ? _slots_17_io_out_uop_lrs2_rtype
         : _GEN_36 ? _slots_16_io_out_uop_lrs2_rtype : _slots_15_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_37
         ? _slots_17_io_out_uop_frs3_en
         : _GEN_36 ? _slots_16_io_out_uop_frs3_en : _slots_15_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_37
         ? _slots_17_io_out_uop_fp_val
         : _GEN_36 ? _slots_16_io_out_uop_fp_val : _slots_15_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_37
         ? _slots_17_io_out_uop_fp_single
         : _GEN_36 ? _slots_16_io_out_uop_fp_single : _slots_15_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_37
         ? _slots_17_io_out_uop_xcpt_pf_if
         : _GEN_36 ? _slots_16_io_out_uop_xcpt_pf_if : _slots_15_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_37
         ? _slots_17_io_out_uop_xcpt_ae_if
         : _GEN_36 ? _slots_16_io_out_uop_xcpt_ae_if : _slots_15_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_37
         ? _slots_17_io_out_uop_xcpt_ma_if
         : _GEN_36 ? _slots_16_io_out_uop_xcpt_ma_if : _slots_15_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_37
         ? _slots_17_io_out_uop_bp_debug_if
         : _GEN_36 ? _slots_16_io_out_uop_bp_debug_if : _slots_15_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_37
         ? _slots_17_io_out_uop_bp_xcpt_if
         : _GEN_36 ? _slots_16_io_out_uop_bp_xcpt_if : _slots_15_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_37
         ? _slots_17_io_out_uop_debug_fsrc
         : _GEN_36 ? _slots_16_io_out_uop_debug_fsrc : _slots_15_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_37
         ? _slots_17_io_out_uop_debug_tsrc
         : _GEN_36 ? _slots_16_io_out_uop_debug_tsrc : _slots_15_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_14_io_valid),
    .io_will_be_valid               (_slots_14_io_will_be_valid),
    .io_request                     (_slots_14_io_request),
    .io_out_uop_uopc                (_slots_14_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_14_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_14_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_14_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_14_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_14_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_14_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_14_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_14_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_14_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_14_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_14_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_14_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_14_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_14_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_14_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_14_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_14_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_14_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_14_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_14_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_14_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_14_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_14_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_14_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_14_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_14_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_14_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_14_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_14_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_14_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_14_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_14_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_14_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_14_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_14_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_14_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_14_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_14_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_14_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_14_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_14_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_14_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_14_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_14_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_14_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_14_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_14_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_14_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_14_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_14_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_14_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_14_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_14_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_14_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_14_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_14_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_14_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_14_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_14_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_14_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_14_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_14_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_14_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_14_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_14_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_14_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_14_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_14_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_14_io_uop_uopc),
    .io_uop_inst                    (_slots_14_io_uop_inst),
    .io_uop_debug_inst              (_slots_14_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_14_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_14_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_14_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_14_io_uop_fu_code),
    .io_uop_iw_state                (_slots_14_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_14_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_14_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_14_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_14_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_14_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_14_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_14_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_14_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_14_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_14_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_14_io_uop_pc_lob),
    .io_uop_taken                   (_slots_14_io_uop_taken),
    .io_uop_imm_packed              (_slots_14_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_14_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_14_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_14_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_14_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_14_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_14_io_uop_pdst),
    .io_uop_prs1                    (_slots_14_io_uop_prs1),
    .io_uop_prs2                    (_slots_14_io_uop_prs2),
    .io_uop_prs3                    (_slots_14_io_uop_prs3),
    .io_uop_ppred                   (_slots_14_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_14_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_14_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_14_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_14_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_14_io_uop_stale_pdst),
    .io_uop_exception               (_slots_14_io_uop_exception),
    .io_uop_exc_cause               (_slots_14_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_14_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_14_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_14_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_14_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_14_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_14_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_14_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_14_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_14_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_14_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_14_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_14_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_14_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_14_io_uop_ldst),
    .io_uop_lrs1                    (_slots_14_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_14_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_14_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_14_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_14_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_14_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_14_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_14_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_14_io_uop_fp_val),
    .io_uop_fp_single               (_slots_14_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_14_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_14_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_14_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_14_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_14_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_14_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_14_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_15 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_15_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_14),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_15_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_39
         ? _slots_18_io_out_uop_uopc
         : _GEN_38 ? _slots_17_io_out_uop_uopc : _slots_16_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_39
         ? _slots_18_io_out_uop_inst
         : _GEN_38 ? _slots_17_io_out_uop_inst : _slots_16_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_39
         ? _slots_18_io_out_uop_debug_inst
         : _GEN_38 ? _slots_17_io_out_uop_debug_inst : _slots_16_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_39
         ? _slots_18_io_out_uop_is_rvc
         : _GEN_38 ? _slots_17_io_out_uop_is_rvc : _slots_16_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_39
         ? _slots_18_io_out_uop_debug_pc
         : _GEN_38 ? _slots_17_io_out_uop_debug_pc : _slots_16_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_39
         ? _slots_18_io_out_uop_iq_type
         : _GEN_38 ? _slots_17_io_out_uop_iq_type : _slots_16_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_39
         ? _slots_18_io_out_uop_fu_code
         : _GEN_38 ? _slots_17_io_out_uop_fu_code : _slots_16_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_39
         ? _slots_18_io_out_uop_iw_state
         : _GEN_38 ? _slots_17_io_out_uop_iw_state : _slots_16_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_39
         ? _slots_18_io_out_uop_iw_p1_poisoned
         : _GEN_38
             ? _slots_17_io_out_uop_iw_p1_poisoned
             : _slots_16_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_39
         ? _slots_18_io_out_uop_iw_p2_poisoned
         : _GEN_38
             ? _slots_17_io_out_uop_iw_p2_poisoned
             : _slots_16_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_39
         ? _slots_18_io_out_uop_is_br
         : _GEN_38 ? _slots_17_io_out_uop_is_br : _slots_16_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_39
         ? _slots_18_io_out_uop_is_jalr
         : _GEN_38 ? _slots_17_io_out_uop_is_jalr : _slots_16_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_39
         ? _slots_18_io_out_uop_is_jal
         : _GEN_38 ? _slots_17_io_out_uop_is_jal : _slots_16_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_39
         ? _slots_18_io_out_uop_is_sfb
         : _GEN_38 ? _slots_17_io_out_uop_is_sfb : _slots_16_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_39
         ? _slots_18_io_out_uop_br_mask
         : _GEN_38 ? _slots_17_io_out_uop_br_mask : _slots_16_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_39
         ? _slots_18_io_out_uop_br_tag
         : _GEN_38 ? _slots_17_io_out_uop_br_tag : _slots_16_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_39
         ? _slots_18_io_out_uop_ftq_idx
         : _GEN_38 ? _slots_17_io_out_uop_ftq_idx : _slots_16_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_39
         ? _slots_18_io_out_uop_edge_inst
         : _GEN_38 ? _slots_17_io_out_uop_edge_inst : _slots_16_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_39
         ? _slots_18_io_out_uop_pc_lob
         : _GEN_38 ? _slots_17_io_out_uop_pc_lob : _slots_16_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_39
         ? _slots_18_io_out_uop_taken
         : _GEN_38 ? _slots_17_io_out_uop_taken : _slots_16_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_39
         ? _slots_18_io_out_uop_imm_packed
         : _GEN_38 ? _slots_17_io_out_uop_imm_packed : _slots_16_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_39
         ? _slots_18_io_out_uop_csr_addr
         : _GEN_38 ? _slots_17_io_out_uop_csr_addr : _slots_16_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_39
         ? _slots_18_io_out_uop_rob_idx
         : _GEN_38 ? _slots_17_io_out_uop_rob_idx : _slots_16_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_39
         ? _slots_18_io_out_uop_ldq_idx
         : _GEN_38 ? _slots_17_io_out_uop_ldq_idx : _slots_16_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_39
         ? _slots_18_io_out_uop_stq_idx
         : _GEN_38 ? _slots_17_io_out_uop_stq_idx : _slots_16_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_39
         ? _slots_18_io_out_uop_rxq_idx
         : _GEN_38 ? _slots_17_io_out_uop_rxq_idx : _slots_16_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_39
         ? _slots_18_io_out_uop_pdst
         : _GEN_38 ? _slots_17_io_out_uop_pdst : _slots_16_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_39
         ? _slots_18_io_out_uop_prs1
         : _GEN_38 ? _slots_17_io_out_uop_prs1 : _slots_16_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_39
         ? _slots_18_io_out_uop_prs2
         : _GEN_38 ? _slots_17_io_out_uop_prs2 : _slots_16_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_39
         ? _slots_18_io_out_uop_prs3
         : _GEN_38 ? _slots_17_io_out_uop_prs3 : _slots_16_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_39
         ? _slots_18_io_out_uop_ppred
         : _GEN_38 ? _slots_17_io_out_uop_ppred : _slots_16_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_39
         ? _slots_18_io_out_uop_prs1_busy
         : _GEN_38 ? _slots_17_io_out_uop_prs1_busy : _slots_16_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_39
         ? _slots_18_io_out_uop_prs2_busy
         : _GEN_38 ? _slots_17_io_out_uop_prs2_busy : _slots_16_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_39
         ? _slots_18_io_out_uop_prs3_busy
         : _GEN_38 ? _slots_17_io_out_uop_prs3_busy : _slots_16_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_39
         ? _slots_18_io_out_uop_ppred_busy
         : _GEN_38 ? _slots_17_io_out_uop_ppred_busy : _slots_16_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_39
         ? _slots_18_io_out_uop_stale_pdst
         : _GEN_38 ? _slots_17_io_out_uop_stale_pdst : _slots_16_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_39
         ? _slots_18_io_out_uop_exception
         : _GEN_38 ? _slots_17_io_out_uop_exception : _slots_16_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_39
         ? _slots_18_io_out_uop_exc_cause
         : _GEN_38 ? _slots_17_io_out_uop_exc_cause : _slots_16_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_39
         ? _slots_18_io_out_uop_bypassable
         : _GEN_38 ? _slots_17_io_out_uop_bypassable : _slots_16_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_39
         ? _slots_18_io_out_uop_mem_cmd
         : _GEN_38 ? _slots_17_io_out_uop_mem_cmd : _slots_16_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_39
         ? _slots_18_io_out_uop_mem_size
         : _GEN_38 ? _slots_17_io_out_uop_mem_size : _slots_16_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_39
         ? _slots_18_io_out_uop_mem_signed
         : _GEN_38 ? _slots_17_io_out_uop_mem_signed : _slots_16_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_39
         ? _slots_18_io_out_uop_is_fence
         : _GEN_38 ? _slots_17_io_out_uop_is_fence : _slots_16_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_39
         ? _slots_18_io_out_uop_is_fencei
         : _GEN_38 ? _slots_17_io_out_uop_is_fencei : _slots_16_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_39
         ? _slots_18_io_out_uop_is_amo
         : _GEN_38 ? _slots_17_io_out_uop_is_amo : _slots_16_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_39
         ? _slots_18_io_out_uop_uses_ldq
         : _GEN_38 ? _slots_17_io_out_uop_uses_ldq : _slots_16_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_39
         ? _slots_18_io_out_uop_uses_stq
         : _GEN_38 ? _slots_17_io_out_uop_uses_stq : _slots_16_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_39
         ? _slots_18_io_out_uop_is_sys_pc2epc
         : _GEN_38
             ? _slots_17_io_out_uop_is_sys_pc2epc
             : _slots_16_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_39
         ? _slots_18_io_out_uop_is_unique
         : _GEN_38 ? _slots_17_io_out_uop_is_unique : _slots_16_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_39
         ? _slots_18_io_out_uop_flush_on_commit
         : _GEN_38
             ? _slots_17_io_out_uop_flush_on_commit
             : _slots_16_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_39
         ? _slots_18_io_out_uop_ldst_is_rs1
         : _GEN_38 ? _slots_17_io_out_uop_ldst_is_rs1 : _slots_16_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_39
         ? _slots_18_io_out_uop_ldst
         : _GEN_38 ? _slots_17_io_out_uop_ldst : _slots_16_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_39
         ? _slots_18_io_out_uop_lrs1
         : _GEN_38 ? _slots_17_io_out_uop_lrs1 : _slots_16_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_39
         ? _slots_18_io_out_uop_lrs2
         : _GEN_38 ? _slots_17_io_out_uop_lrs2 : _slots_16_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_39
         ? _slots_18_io_out_uop_lrs3
         : _GEN_38 ? _slots_17_io_out_uop_lrs3 : _slots_16_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_39
         ? _slots_18_io_out_uop_ldst_val
         : _GEN_38 ? _slots_17_io_out_uop_ldst_val : _slots_16_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_39
         ? _slots_18_io_out_uop_dst_rtype
         : _GEN_38 ? _slots_17_io_out_uop_dst_rtype : _slots_16_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_39
         ? _slots_18_io_out_uop_lrs1_rtype
         : _GEN_38 ? _slots_17_io_out_uop_lrs1_rtype : _slots_16_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_39
         ? _slots_18_io_out_uop_lrs2_rtype
         : _GEN_38 ? _slots_17_io_out_uop_lrs2_rtype : _slots_16_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_39
         ? _slots_18_io_out_uop_frs3_en
         : _GEN_38 ? _slots_17_io_out_uop_frs3_en : _slots_16_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_39
         ? _slots_18_io_out_uop_fp_val
         : _GEN_38 ? _slots_17_io_out_uop_fp_val : _slots_16_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_39
         ? _slots_18_io_out_uop_fp_single
         : _GEN_38 ? _slots_17_io_out_uop_fp_single : _slots_16_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_39
         ? _slots_18_io_out_uop_xcpt_pf_if
         : _GEN_38 ? _slots_17_io_out_uop_xcpt_pf_if : _slots_16_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_39
         ? _slots_18_io_out_uop_xcpt_ae_if
         : _GEN_38 ? _slots_17_io_out_uop_xcpt_ae_if : _slots_16_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_39
         ? _slots_18_io_out_uop_xcpt_ma_if
         : _GEN_38 ? _slots_17_io_out_uop_xcpt_ma_if : _slots_16_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_39
         ? _slots_18_io_out_uop_bp_debug_if
         : _GEN_38 ? _slots_17_io_out_uop_bp_debug_if : _slots_16_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_39
         ? _slots_18_io_out_uop_bp_xcpt_if
         : _GEN_38 ? _slots_17_io_out_uop_bp_xcpt_if : _slots_16_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_39
         ? _slots_18_io_out_uop_debug_fsrc
         : _GEN_38 ? _slots_17_io_out_uop_debug_fsrc : _slots_16_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_39
         ? _slots_18_io_out_uop_debug_tsrc
         : _GEN_38 ? _slots_17_io_out_uop_debug_tsrc : _slots_16_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_15_io_valid),
    .io_will_be_valid               (_slots_15_io_will_be_valid),
    .io_request                     (_slots_15_io_request),
    .io_out_uop_uopc                (_slots_15_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_15_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_15_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_15_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_15_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_15_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_15_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_15_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_15_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_15_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_15_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_15_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_15_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_15_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_15_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_15_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_15_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_15_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_15_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_15_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_15_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_15_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_15_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_15_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_15_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_15_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_15_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_15_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_15_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_15_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_15_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_15_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_15_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_15_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_15_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_15_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_15_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_15_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_15_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_15_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_15_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_15_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_15_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_15_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_15_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_15_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_15_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_15_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_15_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_15_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_15_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_15_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_15_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_15_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_15_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_15_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_15_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_15_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_15_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_15_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_15_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_15_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_15_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_15_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_15_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_15_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_15_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_15_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_15_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_15_io_uop_uopc),
    .io_uop_inst                    (_slots_15_io_uop_inst),
    .io_uop_debug_inst              (_slots_15_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_15_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_15_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_15_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_15_io_uop_fu_code),
    .io_uop_iw_state                (_slots_15_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_15_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_15_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_15_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_15_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_15_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_15_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_15_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_15_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_15_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_15_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_15_io_uop_pc_lob),
    .io_uop_taken                   (_slots_15_io_uop_taken),
    .io_uop_imm_packed              (_slots_15_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_15_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_15_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_15_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_15_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_15_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_15_io_uop_pdst),
    .io_uop_prs1                    (_slots_15_io_uop_prs1),
    .io_uop_prs2                    (_slots_15_io_uop_prs2),
    .io_uop_prs3                    (_slots_15_io_uop_prs3),
    .io_uop_ppred                   (_slots_15_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_15_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_15_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_15_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_15_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_15_io_uop_stale_pdst),
    .io_uop_exception               (_slots_15_io_uop_exception),
    .io_uop_exc_cause               (_slots_15_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_15_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_15_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_15_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_15_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_15_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_15_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_15_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_15_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_15_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_15_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_15_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_15_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_15_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_15_io_uop_ldst),
    .io_uop_lrs1                    (_slots_15_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_15_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_15_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_15_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_15_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_15_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_15_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_15_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_15_io_uop_fp_val),
    .io_uop_fp_single               (_slots_15_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_15_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_15_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_15_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_15_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_15_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_15_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_15_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_16 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_16_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_15),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_16_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_41
         ? _slots_19_io_out_uop_uopc
         : _GEN_40 ? _slots_18_io_out_uop_uopc : _slots_17_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_41
         ? _slots_19_io_out_uop_inst
         : _GEN_40 ? _slots_18_io_out_uop_inst : _slots_17_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_41
         ? _slots_19_io_out_uop_debug_inst
         : _GEN_40 ? _slots_18_io_out_uop_debug_inst : _slots_17_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_41
         ? _slots_19_io_out_uop_is_rvc
         : _GEN_40 ? _slots_18_io_out_uop_is_rvc : _slots_17_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_41
         ? _slots_19_io_out_uop_debug_pc
         : _GEN_40 ? _slots_18_io_out_uop_debug_pc : _slots_17_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_41
         ? _slots_19_io_out_uop_iq_type
         : _GEN_40 ? _slots_18_io_out_uop_iq_type : _slots_17_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_41
         ? _slots_19_io_out_uop_fu_code
         : _GEN_40 ? _slots_18_io_out_uop_fu_code : _slots_17_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_41
         ? _slots_19_io_out_uop_iw_state
         : _GEN_40 ? _slots_18_io_out_uop_iw_state : _slots_17_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_41
         ? _slots_19_io_out_uop_iw_p1_poisoned
         : _GEN_40
             ? _slots_18_io_out_uop_iw_p1_poisoned
             : _slots_17_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_41
         ? _slots_19_io_out_uop_iw_p2_poisoned
         : _GEN_40
             ? _slots_18_io_out_uop_iw_p2_poisoned
             : _slots_17_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_41
         ? _slots_19_io_out_uop_is_br
         : _GEN_40 ? _slots_18_io_out_uop_is_br : _slots_17_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_41
         ? _slots_19_io_out_uop_is_jalr
         : _GEN_40 ? _slots_18_io_out_uop_is_jalr : _slots_17_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_41
         ? _slots_19_io_out_uop_is_jal
         : _GEN_40 ? _slots_18_io_out_uop_is_jal : _slots_17_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_41
         ? _slots_19_io_out_uop_is_sfb
         : _GEN_40 ? _slots_18_io_out_uop_is_sfb : _slots_17_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_41
         ? _slots_19_io_out_uop_br_mask
         : _GEN_40 ? _slots_18_io_out_uop_br_mask : _slots_17_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_41
         ? _slots_19_io_out_uop_br_tag
         : _GEN_40 ? _slots_18_io_out_uop_br_tag : _slots_17_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_41
         ? _slots_19_io_out_uop_ftq_idx
         : _GEN_40 ? _slots_18_io_out_uop_ftq_idx : _slots_17_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_41
         ? _slots_19_io_out_uop_edge_inst
         : _GEN_40 ? _slots_18_io_out_uop_edge_inst : _slots_17_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_41
         ? _slots_19_io_out_uop_pc_lob
         : _GEN_40 ? _slots_18_io_out_uop_pc_lob : _slots_17_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_41
         ? _slots_19_io_out_uop_taken
         : _GEN_40 ? _slots_18_io_out_uop_taken : _slots_17_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_41
         ? _slots_19_io_out_uop_imm_packed
         : _GEN_40 ? _slots_18_io_out_uop_imm_packed : _slots_17_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_41
         ? _slots_19_io_out_uop_csr_addr
         : _GEN_40 ? _slots_18_io_out_uop_csr_addr : _slots_17_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_41
         ? _slots_19_io_out_uop_rob_idx
         : _GEN_40 ? _slots_18_io_out_uop_rob_idx : _slots_17_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_41
         ? _slots_19_io_out_uop_ldq_idx
         : _GEN_40 ? _slots_18_io_out_uop_ldq_idx : _slots_17_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_41
         ? _slots_19_io_out_uop_stq_idx
         : _GEN_40 ? _slots_18_io_out_uop_stq_idx : _slots_17_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_41
         ? _slots_19_io_out_uop_rxq_idx
         : _GEN_40 ? _slots_18_io_out_uop_rxq_idx : _slots_17_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_41
         ? _slots_19_io_out_uop_pdst
         : _GEN_40 ? _slots_18_io_out_uop_pdst : _slots_17_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_41
         ? _slots_19_io_out_uop_prs1
         : _GEN_40 ? _slots_18_io_out_uop_prs1 : _slots_17_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_41
         ? _slots_19_io_out_uop_prs2
         : _GEN_40 ? _slots_18_io_out_uop_prs2 : _slots_17_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_41
         ? _slots_19_io_out_uop_prs3
         : _GEN_40 ? _slots_18_io_out_uop_prs3 : _slots_17_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_41
         ? _slots_19_io_out_uop_ppred
         : _GEN_40 ? _slots_18_io_out_uop_ppred : _slots_17_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_41
         ? _slots_19_io_out_uop_prs1_busy
         : _GEN_40 ? _slots_18_io_out_uop_prs1_busy : _slots_17_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_41
         ? _slots_19_io_out_uop_prs2_busy
         : _GEN_40 ? _slots_18_io_out_uop_prs2_busy : _slots_17_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_41
         ? _slots_19_io_out_uop_prs3_busy
         : _GEN_40 ? _slots_18_io_out_uop_prs3_busy : _slots_17_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_41
         ? _slots_19_io_out_uop_ppred_busy
         : _GEN_40 ? _slots_18_io_out_uop_ppred_busy : _slots_17_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_41
         ? _slots_19_io_out_uop_stale_pdst
         : _GEN_40 ? _slots_18_io_out_uop_stale_pdst : _slots_17_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_41
         ? _slots_19_io_out_uop_exception
         : _GEN_40 ? _slots_18_io_out_uop_exception : _slots_17_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_41
         ? _slots_19_io_out_uop_exc_cause
         : _GEN_40 ? _slots_18_io_out_uop_exc_cause : _slots_17_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_41
         ? _slots_19_io_out_uop_bypassable
         : _GEN_40 ? _slots_18_io_out_uop_bypassable : _slots_17_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_41
         ? _slots_19_io_out_uop_mem_cmd
         : _GEN_40 ? _slots_18_io_out_uop_mem_cmd : _slots_17_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_41
         ? _slots_19_io_out_uop_mem_size
         : _GEN_40 ? _slots_18_io_out_uop_mem_size : _slots_17_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_41
         ? _slots_19_io_out_uop_mem_signed
         : _GEN_40 ? _slots_18_io_out_uop_mem_signed : _slots_17_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_41
         ? _slots_19_io_out_uop_is_fence
         : _GEN_40 ? _slots_18_io_out_uop_is_fence : _slots_17_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_41
         ? _slots_19_io_out_uop_is_fencei
         : _GEN_40 ? _slots_18_io_out_uop_is_fencei : _slots_17_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_41
         ? _slots_19_io_out_uop_is_amo
         : _GEN_40 ? _slots_18_io_out_uop_is_amo : _slots_17_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_41
         ? _slots_19_io_out_uop_uses_ldq
         : _GEN_40 ? _slots_18_io_out_uop_uses_ldq : _slots_17_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_41
         ? _slots_19_io_out_uop_uses_stq
         : _GEN_40 ? _slots_18_io_out_uop_uses_stq : _slots_17_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_41
         ? _slots_19_io_out_uop_is_sys_pc2epc
         : _GEN_40
             ? _slots_18_io_out_uop_is_sys_pc2epc
             : _slots_17_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_41
         ? _slots_19_io_out_uop_is_unique
         : _GEN_40 ? _slots_18_io_out_uop_is_unique : _slots_17_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_41
         ? _slots_19_io_out_uop_flush_on_commit
         : _GEN_40
             ? _slots_18_io_out_uop_flush_on_commit
             : _slots_17_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_41
         ? _slots_19_io_out_uop_ldst_is_rs1
         : _GEN_40 ? _slots_18_io_out_uop_ldst_is_rs1 : _slots_17_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_41
         ? _slots_19_io_out_uop_ldst
         : _GEN_40 ? _slots_18_io_out_uop_ldst : _slots_17_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_41
         ? _slots_19_io_out_uop_lrs1
         : _GEN_40 ? _slots_18_io_out_uop_lrs1 : _slots_17_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_41
         ? _slots_19_io_out_uop_lrs2
         : _GEN_40 ? _slots_18_io_out_uop_lrs2 : _slots_17_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_41
         ? _slots_19_io_out_uop_lrs3
         : _GEN_40 ? _slots_18_io_out_uop_lrs3 : _slots_17_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_41
         ? _slots_19_io_out_uop_ldst_val
         : _GEN_40 ? _slots_18_io_out_uop_ldst_val : _slots_17_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_41
         ? _slots_19_io_out_uop_dst_rtype
         : _GEN_40 ? _slots_18_io_out_uop_dst_rtype : _slots_17_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_41
         ? _slots_19_io_out_uop_lrs1_rtype
         : _GEN_40 ? _slots_18_io_out_uop_lrs1_rtype : _slots_17_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_41
         ? _slots_19_io_out_uop_lrs2_rtype
         : _GEN_40 ? _slots_18_io_out_uop_lrs2_rtype : _slots_17_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_41
         ? _slots_19_io_out_uop_frs3_en
         : _GEN_40 ? _slots_18_io_out_uop_frs3_en : _slots_17_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_41
         ? _slots_19_io_out_uop_fp_val
         : _GEN_40 ? _slots_18_io_out_uop_fp_val : _slots_17_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_41
         ? _slots_19_io_out_uop_fp_single
         : _GEN_40 ? _slots_18_io_out_uop_fp_single : _slots_17_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_41
         ? _slots_19_io_out_uop_xcpt_pf_if
         : _GEN_40 ? _slots_18_io_out_uop_xcpt_pf_if : _slots_17_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_41
         ? _slots_19_io_out_uop_xcpt_ae_if
         : _GEN_40 ? _slots_18_io_out_uop_xcpt_ae_if : _slots_17_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_41
         ? _slots_19_io_out_uop_xcpt_ma_if
         : _GEN_40 ? _slots_18_io_out_uop_xcpt_ma_if : _slots_17_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_41
         ? _slots_19_io_out_uop_bp_debug_if
         : _GEN_40 ? _slots_18_io_out_uop_bp_debug_if : _slots_17_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_41
         ? _slots_19_io_out_uop_bp_xcpt_if
         : _GEN_40 ? _slots_18_io_out_uop_bp_xcpt_if : _slots_17_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_41
         ? _slots_19_io_out_uop_debug_fsrc
         : _GEN_40 ? _slots_18_io_out_uop_debug_fsrc : _slots_17_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_41
         ? _slots_19_io_out_uop_debug_tsrc
         : _GEN_40 ? _slots_18_io_out_uop_debug_tsrc : _slots_17_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_16_io_valid),
    .io_will_be_valid               (_slots_16_io_will_be_valid),
    .io_request                     (_slots_16_io_request),
    .io_out_uop_uopc                (_slots_16_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_16_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_16_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_16_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_16_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_16_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_16_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_16_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_16_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_16_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_16_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_16_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_16_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_16_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_16_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_16_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_16_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_16_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_16_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_16_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_16_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_16_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_16_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_16_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_16_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_16_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_16_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_16_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_16_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_16_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_16_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_16_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_16_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_16_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_16_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_16_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_16_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_16_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_16_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_16_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_16_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_16_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_16_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_16_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_16_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_16_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_16_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_16_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_16_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_16_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_16_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_16_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_16_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_16_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_16_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_16_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_16_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_16_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_16_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_16_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_16_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_16_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_16_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_16_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_16_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_16_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_16_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_16_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_16_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_16_io_uop_uopc),
    .io_uop_inst                    (_slots_16_io_uop_inst),
    .io_uop_debug_inst              (_slots_16_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_16_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_16_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_16_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_16_io_uop_fu_code),
    .io_uop_iw_state                (_slots_16_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_16_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_16_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_16_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_16_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_16_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_16_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_16_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_16_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_16_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_16_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_16_io_uop_pc_lob),
    .io_uop_taken                   (_slots_16_io_uop_taken),
    .io_uop_imm_packed              (_slots_16_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_16_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_16_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_16_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_16_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_16_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_16_io_uop_pdst),
    .io_uop_prs1                    (_slots_16_io_uop_prs1),
    .io_uop_prs2                    (_slots_16_io_uop_prs2),
    .io_uop_prs3                    (_slots_16_io_uop_prs3),
    .io_uop_ppred                   (_slots_16_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_16_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_16_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_16_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_16_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_16_io_uop_stale_pdst),
    .io_uop_exception               (_slots_16_io_uop_exception),
    .io_uop_exc_cause               (_slots_16_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_16_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_16_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_16_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_16_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_16_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_16_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_16_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_16_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_16_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_16_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_16_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_16_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_16_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_16_io_uop_ldst),
    .io_uop_lrs1                    (_slots_16_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_16_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_16_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_16_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_16_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_16_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_16_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_16_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_16_io_uop_fp_val),
    .io_uop_fp_single               (_slots_16_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_16_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_16_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_16_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_16_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_16_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_16_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_16_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_17 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_17_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_16),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_17_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_43
         ? _slots_20_io_out_uop_uopc
         : _GEN_42 ? _slots_19_io_out_uop_uopc : _slots_18_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_43
         ? _slots_20_io_out_uop_inst
         : _GEN_42 ? _slots_19_io_out_uop_inst : _slots_18_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_43
         ? _slots_20_io_out_uop_debug_inst
         : _GEN_42 ? _slots_19_io_out_uop_debug_inst : _slots_18_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_43
         ? _slots_20_io_out_uop_is_rvc
         : _GEN_42 ? _slots_19_io_out_uop_is_rvc : _slots_18_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_43
         ? _slots_20_io_out_uop_debug_pc
         : _GEN_42 ? _slots_19_io_out_uop_debug_pc : _slots_18_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_43
         ? _slots_20_io_out_uop_iq_type
         : _GEN_42 ? _slots_19_io_out_uop_iq_type : _slots_18_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_43
         ? _slots_20_io_out_uop_fu_code
         : _GEN_42 ? _slots_19_io_out_uop_fu_code : _slots_18_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_43
         ? _slots_20_io_out_uop_iw_state
         : _GEN_42 ? _slots_19_io_out_uop_iw_state : _slots_18_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_43
         ? _slots_20_io_out_uop_iw_p1_poisoned
         : _GEN_42
             ? _slots_19_io_out_uop_iw_p1_poisoned
             : _slots_18_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_43
         ? _slots_20_io_out_uop_iw_p2_poisoned
         : _GEN_42
             ? _slots_19_io_out_uop_iw_p2_poisoned
             : _slots_18_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_43
         ? _slots_20_io_out_uop_is_br
         : _GEN_42 ? _slots_19_io_out_uop_is_br : _slots_18_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_43
         ? _slots_20_io_out_uop_is_jalr
         : _GEN_42 ? _slots_19_io_out_uop_is_jalr : _slots_18_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_43
         ? _slots_20_io_out_uop_is_jal
         : _GEN_42 ? _slots_19_io_out_uop_is_jal : _slots_18_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_43
         ? _slots_20_io_out_uop_is_sfb
         : _GEN_42 ? _slots_19_io_out_uop_is_sfb : _slots_18_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_43
         ? _slots_20_io_out_uop_br_mask
         : _GEN_42 ? _slots_19_io_out_uop_br_mask : _slots_18_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_43
         ? _slots_20_io_out_uop_br_tag
         : _GEN_42 ? _slots_19_io_out_uop_br_tag : _slots_18_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_43
         ? _slots_20_io_out_uop_ftq_idx
         : _GEN_42 ? _slots_19_io_out_uop_ftq_idx : _slots_18_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_43
         ? _slots_20_io_out_uop_edge_inst
         : _GEN_42 ? _slots_19_io_out_uop_edge_inst : _slots_18_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_43
         ? _slots_20_io_out_uop_pc_lob
         : _GEN_42 ? _slots_19_io_out_uop_pc_lob : _slots_18_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_43
         ? _slots_20_io_out_uop_taken
         : _GEN_42 ? _slots_19_io_out_uop_taken : _slots_18_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_43
         ? _slots_20_io_out_uop_imm_packed
         : _GEN_42 ? _slots_19_io_out_uop_imm_packed : _slots_18_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_43
         ? _slots_20_io_out_uop_csr_addr
         : _GEN_42 ? _slots_19_io_out_uop_csr_addr : _slots_18_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_43
         ? _slots_20_io_out_uop_rob_idx
         : _GEN_42 ? _slots_19_io_out_uop_rob_idx : _slots_18_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_43
         ? _slots_20_io_out_uop_ldq_idx
         : _GEN_42 ? _slots_19_io_out_uop_ldq_idx : _slots_18_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_43
         ? _slots_20_io_out_uop_stq_idx
         : _GEN_42 ? _slots_19_io_out_uop_stq_idx : _slots_18_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_43
         ? _slots_20_io_out_uop_rxq_idx
         : _GEN_42 ? _slots_19_io_out_uop_rxq_idx : _slots_18_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_43
         ? _slots_20_io_out_uop_pdst
         : _GEN_42 ? _slots_19_io_out_uop_pdst : _slots_18_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_43
         ? _slots_20_io_out_uop_prs1
         : _GEN_42 ? _slots_19_io_out_uop_prs1 : _slots_18_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_43
         ? _slots_20_io_out_uop_prs2
         : _GEN_42 ? _slots_19_io_out_uop_prs2 : _slots_18_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_43
         ? _slots_20_io_out_uop_prs3
         : _GEN_42 ? _slots_19_io_out_uop_prs3 : _slots_18_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_43
         ? _slots_20_io_out_uop_ppred
         : _GEN_42 ? _slots_19_io_out_uop_ppred : _slots_18_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_43
         ? _slots_20_io_out_uop_prs1_busy
         : _GEN_42 ? _slots_19_io_out_uop_prs1_busy : _slots_18_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_43
         ? _slots_20_io_out_uop_prs2_busy
         : _GEN_42 ? _slots_19_io_out_uop_prs2_busy : _slots_18_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_43
         ? _slots_20_io_out_uop_prs3_busy
         : _GEN_42 ? _slots_19_io_out_uop_prs3_busy : _slots_18_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_43
         ? _slots_20_io_out_uop_ppred_busy
         : _GEN_42 ? _slots_19_io_out_uop_ppred_busy : _slots_18_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_43
         ? _slots_20_io_out_uop_stale_pdst
         : _GEN_42 ? _slots_19_io_out_uop_stale_pdst : _slots_18_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_43
         ? _slots_20_io_out_uop_exception
         : _GEN_42 ? _slots_19_io_out_uop_exception : _slots_18_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_43
         ? _slots_20_io_out_uop_exc_cause
         : _GEN_42 ? _slots_19_io_out_uop_exc_cause : _slots_18_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_43
         ? _slots_20_io_out_uop_bypassable
         : _GEN_42 ? _slots_19_io_out_uop_bypassable : _slots_18_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_43
         ? _slots_20_io_out_uop_mem_cmd
         : _GEN_42 ? _slots_19_io_out_uop_mem_cmd : _slots_18_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_43
         ? _slots_20_io_out_uop_mem_size
         : _GEN_42 ? _slots_19_io_out_uop_mem_size : _slots_18_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_43
         ? _slots_20_io_out_uop_mem_signed
         : _GEN_42 ? _slots_19_io_out_uop_mem_signed : _slots_18_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_43
         ? _slots_20_io_out_uop_is_fence
         : _GEN_42 ? _slots_19_io_out_uop_is_fence : _slots_18_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_43
         ? _slots_20_io_out_uop_is_fencei
         : _GEN_42 ? _slots_19_io_out_uop_is_fencei : _slots_18_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_43
         ? _slots_20_io_out_uop_is_amo
         : _GEN_42 ? _slots_19_io_out_uop_is_amo : _slots_18_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_43
         ? _slots_20_io_out_uop_uses_ldq
         : _GEN_42 ? _slots_19_io_out_uop_uses_ldq : _slots_18_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_43
         ? _slots_20_io_out_uop_uses_stq
         : _GEN_42 ? _slots_19_io_out_uop_uses_stq : _slots_18_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_43
         ? _slots_20_io_out_uop_is_sys_pc2epc
         : _GEN_42
             ? _slots_19_io_out_uop_is_sys_pc2epc
             : _slots_18_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_43
         ? _slots_20_io_out_uop_is_unique
         : _GEN_42 ? _slots_19_io_out_uop_is_unique : _slots_18_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_43
         ? _slots_20_io_out_uop_flush_on_commit
         : _GEN_42
             ? _slots_19_io_out_uop_flush_on_commit
             : _slots_18_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_43
         ? _slots_20_io_out_uop_ldst_is_rs1
         : _GEN_42 ? _slots_19_io_out_uop_ldst_is_rs1 : _slots_18_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_43
         ? _slots_20_io_out_uop_ldst
         : _GEN_42 ? _slots_19_io_out_uop_ldst : _slots_18_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_43
         ? _slots_20_io_out_uop_lrs1
         : _GEN_42 ? _slots_19_io_out_uop_lrs1 : _slots_18_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_43
         ? _slots_20_io_out_uop_lrs2
         : _GEN_42 ? _slots_19_io_out_uop_lrs2 : _slots_18_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_43
         ? _slots_20_io_out_uop_lrs3
         : _GEN_42 ? _slots_19_io_out_uop_lrs3 : _slots_18_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_43
         ? _slots_20_io_out_uop_ldst_val
         : _GEN_42 ? _slots_19_io_out_uop_ldst_val : _slots_18_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_43
         ? _slots_20_io_out_uop_dst_rtype
         : _GEN_42 ? _slots_19_io_out_uop_dst_rtype : _slots_18_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_43
         ? _slots_20_io_out_uop_lrs1_rtype
         : _GEN_42 ? _slots_19_io_out_uop_lrs1_rtype : _slots_18_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_43
         ? _slots_20_io_out_uop_lrs2_rtype
         : _GEN_42 ? _slots_19_io_out_uop_lrs2_rtype : _slots_18_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_43
         ? _slots_20_io_out_uop_frs3_en
         : _GEN_42 ? _slots_19_io_out_uop_frs3_en : _slots_18_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_43
         ? _slots_20_io_out_uop_fp_val
         : _GEN_42 ? _slots_19_io_out_uop_fp_val : _slots_18_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_43
         ? _slots_20_io_out_uop_fp_single
         : _GEN_42 ? _slots_19_io_out_uop_fp_single : _slots_18_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_43
         ? _slots_20_io_out_uop_xcpt_pf_if
         : _GEN_42 ? _slots_19_io_out_uop_xcpt_pf_if : _slots_18_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_43
         ? _slots_20_io_out_uop_xcpt_ae_if
         : _GEN_42 ? _slots_19_io_out_uop_xcpt_ae_if : _slots_18_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_43
         ? _slots_20_io_out_uop_xcpt_ma_if
         : _GEN_42 ? _slots_19_io_out_uop_xcpt_ma_if : _slots_18_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_43
         ? _slots_20_io_out_uop_bp_debug_if
         : _GEN_42 ? _slots_19_io_out_uop_bp_debug_if : _slots_18_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_43
         ? _slots_20_io_out_uop_bp_xcpt_if
         : _GEN_42 ? _slots_19_io_out_uop_bp_xcpt_if : _slots_18_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_43
         ? _slots_20_io_out_uop_debug_fsrc
         : _GEN_42 ? _slots_19_io_out_uop_debug_fsrc : _slots_18_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_43
         ? _slots_20_io_out_uop_debug_tsrc
         : _GEN_42 ? _slots_19_io_out_uop_debug_tsrc : _slots_18_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_17_io_valid),
    .io_will_be_valid               (_slots_17_io_will_be_valid),
    .io_request                     (_slots_17_io_request),
    .io_out_uop_uopc                (_slots_17_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_17_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_17_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_17_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_17_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_17_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_17_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_17_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_17_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_17_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_17_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_17_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_17_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_17_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_17_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_17_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_17_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_17_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_17_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_17_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_17_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_17_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_17_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_17_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_17_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_17_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_17_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_17_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_17_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_17_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_17_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_17_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_17_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_17_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_17_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_17_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_17_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_17_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_17_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_17_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_17_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_17_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_17_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_17_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_17_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_17_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_17_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_17_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_17_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_17_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_17_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_17_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_17_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_17_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_17_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_17_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_17_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_17_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_17_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_17_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_17_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_17_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_17_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_17_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_17_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_17_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_17_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_17_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_17_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_17_io_uop_uopc),
    .io_uop_inst                    (_slots_17_io_uop_inst),
    .io_uop_debug_inst              (_slots_17_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_17_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_17_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_17_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_17_io_uop_fu_code),
    .io_uop_iw_state                (_slots_17_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_17_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_17_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_17_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_17_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_17_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_17_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_17_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_17_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_17_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_17_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_17_io_uop_pc_lob),
    .io_uop_taken                   (_slots_17_io_uop_taken),
    .io_uop_imm_packed              (_slots_17_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_17_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_17_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_17_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_17_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_17_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_17_io_uop_pdst),
    .io_uop_prs1                    (_slots_17_io_uop_prs1),
    .io_uop_prs2                    (_slots_17_io_uop_prs2),
    .io_uop_prs3                    (_slots_17_io_uop_prs3),
    .io_uop_ppred                   (_slots_17_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_17_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_17_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_17_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_17_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_17_io_uop_stale_pdst),
    .io_uop_exception               (_slots_17_io_uop_exception),
    .io_uop_exc_cause               (_slots_17_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_17_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_17_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_17_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_17_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_17_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_17_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_17_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_17_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_17_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_17_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_17_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_17_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_17_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_17_io_uop_ldst),
    .io_uop_lrs1                    (_slots_17_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_17_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_17_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_17_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_17_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_17_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_17_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_17_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_17_io_uop_fp_val),
    .io_uop_fp_single               (_slots_17_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_17_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_17_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_17_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_17_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_17_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_17_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_17_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_18 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_18_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_17),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_18_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_45
         ? _slots_21_io_out_uop_uopc
         : _GEN_44 ? _slots_20_io_out_uop_uopc : _slots_19_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_45
         ? _slots_21_io_out_uop_inst
         : _GEN_44 ? _slots_20_io_out_uop_inst : _slots_19_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_45
         ? _slots_21_io_out_uop_debug_inst
         : _GEN_44 ? _slots_20_io_out_uop_debug_inst : _slots_19_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_45
         ? _slots_21_io_out_uop_is_rvc
         : _GEN_44 ? _slots_20_io_out_uop_is_rvc : _slots_19_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_45
         ? _slots_21_io_out_uop_debug_pc
         : _GEN_44 ? _slots_20_io_out_uop_debug_pc : _slots_19_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_45
         ? _slots_21_io_out_uop_iq_type
         : _GEN_44 ? _slots_20_io_out_uop_iq_type : _slots_19_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_45
         ? _slots_21_io_out_uop_fu_code
         : _GEN_44 ? _slots_20_io_out_uop_fu_code : _slots_19_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_45
         ? _slots_21_io_out_uop_iw_state
         : _GEN_44 ? _slots_20_io_out_uop_iw_state : _slots_19_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_45
         ? _slots_21_io_out_uop_iw_p1_poisoned
         : _GEN_44
             ? _slots_20_io_out_uop_iw_p1_poisoned
             : _slots_19_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_45
         ? _slots_21_io_out_uop_iw_p2_poisoned
         : _GEN_44
             ? _slots_20_io_out_uop_iw_p2_poisoned
             : _slots_19_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_45
         ? _slots_21_io_out_uop_is_br
         : _GEN_44 ? _slots_20_io_out_uop_is_br : _slots_19_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_45
         ? _slots_21_io_out_uop_is_jalr
         : _GEN_44 ? _slots_20_io_out_uop_is_jalr : _slots_19_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_45
         ? _slots_21_io_out_uop_is_jal
         : _GEN_44 ? _slots_20_io_out_uop_is_jal : _slots_19_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_45
         ? _slots_21_io_out_uop_is_sfb
         : _GEN_44 ? _slots_20_io_out_uop_is_sfb : _slots_19_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_45
         ? _slots_21_io_out_uop_br_mask
         : _GEN_44 ? _slots_20_io_out_uop_br_mask : _slots_19_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_45
         ? _slots_21_io_out_uop_br_tag
         : _GEN_44 ? _slots_20_io_out_uop_br_tag : _slots_19_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_45
         ? _slots_21_io_out_uop_ftq_idx
         : _GEN_44 ? _slots_20_io_out_uop_ftq_idx : _slots_19_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_45
         ? _slots_21_io_out_uop_edge_inst
         : _GEN_44 ? _slots_20_io_out_uop_edge_inst : _slots_19_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_45
         ? _slots_21_io_out_uop_pc_lob
         : _GEN_44 ? _slots_20_io_out_uop_pc_lob : _slots_19_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_45
         ? _slots_21_io_out_uop_taken
         : _GEN_44 ? _slots_20_io_out_uop_taken : _slots_19_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_45
         ? _slots_21_io_out_uop_imm_packed
         : _GEN_44 ? _slots_20_io_out_uop_imm_packed : _slots_19_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_45
         ? _slots_21_io_out_uop_csr_addr
         : _GEN_44 ? _slots_20_io_out_uop_csr_addr : _slots_19_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_45
         ? _slots_21_io_out_uop_rob_idx
         : _GEN_44 ? _slots_20_io_out_uop_rob_idx : _slots_19_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_45
         ? _slots_21_io_out_uop_ldq_idx
         : _GEN_44 ? _slots_20_io_out_uop_ldq_idx : _slots_19_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_45
         ? _slots_21_io_out_uop_stq_idx
         : _GEN_44 ? _slots_20_io_out_uop_stq_idx : _slots_19_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_45
         ? _slots_21_io_out_uop_rxq_idx
         : _GEN_44 ? _slots_20_io_out_uop_rxq_idx : _slots_19_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_45
         ? _slots_21_io_out_uop_pdst
         : _GEN_44 ? _slots_20_io_out_uop_pdst : _slots_19_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_45
         ? _slots_21_io_out_uop_prs1
         : _GEN_44 ? _slots_20_io_out_uop_prs1 : _slots_19_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_45
         ? _slots_21_io_out_uop_prs2
         : _GEN_44 ? _slots_20_io_out_uop_prs2 : _slots_19_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_45
         ? _slots_21_io_out_uop_prs3
         : _GEN_44 ? _slots_20_io_out_uop_prs3 : _slots_19_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_45
         ? _slots_21_io_out_uop_ppred
         : _GEN_44 ? _slots_20_io_out_uop_ppred : _slots_19_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_45
         ? _slots_21_io_out_uop_prs1_busy
         : _GEN_44 ? _slots_20_io_out_uop_prs1_busy : _slots_19_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_45
         ? _slots_21_io_out_uop_prs2_busy
         : _GEN_44 ? _slots_20_io_out_uop_prs2_busy : _slots_19_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_45
         ? _slots_21_io_out_uop_prs3_busy
         : _GEN_44 ? _slots_20_io_out_uop_prs3_busy : _slots_19_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_45
         ? _slots_21_io_out_uop_ppred_busy
         : _GEN_44 ? _slots_20_io_out_uop_ppred_busy : _slots_19_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_45
         ? _slots_21_io_out_uop_stale_pdst
         : _GEN_44 ? _slots_20_io_out_uop_stale_pdst : _slots_19_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_45
         ? _slots_21_io_out_uop_exception
         : _GEN_44 ? _slots_20_io_out_uop_exception : _slots_19_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_45
         ? _slots_21_io_out_uop_exc_cause
         : _GEN_44 ? _slots_20_io_out_uop_exc_cause : _slots_19_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_45
         ? _slots_21_io_out_uop_bypassable
         : _GEN_44 ? _slots_20_io_out_uop_bypassable : _slots_19_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_45
         ? _slots_21_io_out_uop_mem_cmd
         : _GEN_44 ? _slots_20_io_out_uop_mem_cmd : _slots_19_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_45
         ? _slots_21_io_out_uop_mem_size
         : _GEN_44 ? _slots_20_io_out_uop_mem_size : _slots_19_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_45
         ? _slots_21_io_out_uop_mem_signed
         : _GEN_44 ? _slots_20_io_out_uop_mem_signed : _slots_19_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_45
         ? _slots_21_io_out_uop_is_fence
         : _GEN_44 ? _slots_20_io_out_uop_is_fence : _slots_19_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_45
         ? _slots_21_io_out_uop_is_fencei
         : _GEN_44 ? _slots_20_io_out_uop_is_fencei : _slots_19_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_45
         ? _slots_21_io_out_uop_is_amo
         : _GEN_44 ? _slots_20_io_out_uop_is_amo : _slots_19_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_45
         ? _slots_21_io_out_uop_uses_ldq
         : _GEN_44 ? _slots_20_io_out_uop_uses_ldq : _slots_19_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_45
         ? _slots_21_io_out_uop_uses_stq
         : _GEN_44 ? _slots_20_io_out_uop_uses_stq : _slots_19_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_45
         ? _slots_21_io_out_uop_is_sys_pc2epc
         : _GEN_44
             ? _slots_20_io_out_uop_is_sys_pc2epc
             : _slots_19_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_45
         ? _slots_21_io_out_uop_is_unique
         : _GEN_44 ? _slots_20_io_out_uop_is_unique : _slots_19_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_45
         ? _slots_21_io_out_uop_flush_on_commit
         : _GEN_44
             ? _slots_20_io_out_uop_flush_on_commit
             : _slots_19_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_45
         ? _slots_21_io_out_uop_ldst_is_rs1
         : _GEN_44 ? _slots_20_io_out_uop_ldst_is_rs1 : _slots_19_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_45
         ? _slots_21_io_out_uop_ldst
         : _GEN_44 ? _slots_20_io_out_uop_ldst : _slots_19_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_45
         ? _slots_21_io_out_uop_lrs1
         : _GEN_44 ? _slots_20_io_out_uop_lrs1 : _slots_19_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_45
         ? _slots_21_io_out_uop_lrs2
         : _GEN_44 ? _slots_20_io_out_uop_lrs2 : _slots_19_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_45
         ? _slots_21_io_out_uop_lrs3
         : _GEN_44 ? _slots_20_io_out_uop_lrs3 : _slots_19_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_45
         ? _slots_21_io_out_uop_ldst_val
         : _GEN_44 ? _slots_20_io_out_uop_ldst_val : _slots_19_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_45
         ? _slots_21_io_out_uop_dst_rtype
         : _GEN_44 ? _slots_20_io_out_uop_dst_rtype : _slots_19_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_45
         ? _slots_21_io_out_uop_lrs1_rtype
         : _GEN_44 ? _slots_20_io_out_uop_lrs1_rtype : _slots_19_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_45
         ? _slots_21_io_out_uop_lrs2_rtype
         : _GEN_44 ? _slots_20_io_out_uop_lrs2_rtype : _slots_19_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_45
         ? _slots_21_io_out_uop_frs3_en
         : _GEN_44 ? _slots_20_io_out_uop_frs3_en : _slots_19_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_45
         ? _slots_21_io_out_uop_fp_val
         : _GEN_44 ? _slots_20_io_out_uop_fp_val : _slots_19_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_45
         ? _slots_21_io_out_uop_fp_single
         : _GEN_44 ? _slots_20_io_out_uop_fp_single : _slots_19_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_45
         ? _slots_21_io_out_uop_xcpt_pf_if
         : _GEN_44 ? _slots_20_io_out_uop_xcpt_pf_if : _slots_19_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_45
         ? _slots_21_io_out_uop_xcpt_ae_if
         : _GEN_44 ? _slots_20_io_out_uop_xcpt_ae_if : _slots_19_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_45
         ? _slots_21_io_out_uop_xcpt_ma_if
         : _GEN_44 ? _slots_20_io_out_uop_xcpt_ma_if : _slots_19_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_45
         ? _slots_21_io_out_uop_bp_debug_if
         : _GEN_44 ? _slots_20_io_out_uop_bp_debug_if : _slots_19_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_45
         ? _slots_21_io_out_uop_bp_xcpt_if
         : _GEN_44 ? _slots_20_io_out_uop_bp_xcpt_if : _slots_19_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_45
         ? _slots_21_io_out_uop_debug_fsrc
         : _GEN_44 ? _slots_20_io_out_uop_debug_fsrc : _slots_19_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_45
         ? _slots_21_io_out_uop_debug_tsrc
         : _GEN_44 ? _slots_20_io_out_uop_debug_tsrc : _slots_19_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_18_io_valid),
    .io_will_be_valid               (_slots_18_io_will_be_valid),
    .io_request                     (_slots_18_io_request),
    .io_out_uop_uopc                (_slots_18_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_18_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_18_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_18_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_18_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_18_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_18_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_18_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_18_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_18_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_18_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_18_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_18_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_18_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_18_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_18_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_18_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_18_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_18_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_18_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_18_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_18_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_18_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_18_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_18_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_18_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_18_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_18_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_18_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_18_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_18_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_18_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_18_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_18_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_18_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_18_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_18_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_18_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_18_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_18_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_18_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_18_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_18_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_18_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_18_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_18_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_18_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_18_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_18_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_18_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_18_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_18_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_18_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_18_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_18_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_18_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_18_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_18_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_18_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_18_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_18_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_18_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_18_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_18_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_18_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_18_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_18_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_18_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_18_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_18_io_uop_uopc),
    .io_uop_inst                    (_slots_18_io_uop_inst),
    .io_uop_debug_inst              (_slots_18_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_18_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_18_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_18_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_18_io_uop_fu_code),
    .io_uop_iw_state                (_slots_18_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_18_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_18_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_18_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_18_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_18_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_18_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_18_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_18_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_18_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_18_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_18_io_uop_pc_lob),
    .io_uop_taken                   (_slots_18_io_uop_taken),
    .io_uop_imm_packed              (_slots_18_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_18_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_18_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_18_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_18_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_18_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_18_io_uop_pdst),
    .io_uop_prs1                    (_slots_18_io_uop_prs1),
    .io_uop_prs2                    (_slots_18_io_uop_prs2),
    .io_uop_prs3                    (_slots_18_io_uop_prs3),
    .io_uop_ppred                   (_slots_18_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_18_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_18_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_18_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_18_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_18_io_uop_stale_pdst),
    .io_uop_exception               (_slots_18_io_uop_exception),
    .io_uop_exc_cause               (_slots_18_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_18_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_18_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_18_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_18_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_18_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_18_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_18_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_18_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_18_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_18_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_18_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_18_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_18_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_18_io_uop_ldst),
    .io_uop_lrs1                    (_slots_18_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_18_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_18_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_18_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_18_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_18_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_18_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_18_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_18_io_uop_fp_val),
    .io_uop_fp_single               (_slots_18_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_18_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_18_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_18_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_18_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_18_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_18_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_18_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_19 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_19_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_18),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_19_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_47
         ? _slots_22_io_out_uop_uopc
         : _GEN_46 ? _slots_21_io_out_uop_uopc : _slots_20_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_47
         ? _slots_22_io_out_uop_inst
         : _GEN_46 ? _slots_21_io_out_uop_inst : _slots_20_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_47
         ? _slots_22_io_out_uop_debug_inst
         : _GEN_46 ? _slots_21_io_out_uop_debug_inst : _slots_20_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_47
         ? _slots_22_io_out_uop_is_rvc
         : _GEN_46 ? _slots_21_io_out_uop_is_rvc : _slots_20_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_47
         ? _slots_22_io_out_uop_debug_pc
         : _GEN_46 ? _slots_21_io_out_uop_debug_pc : _slots_20_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_47
         ? _slots_22_io_out_uop_iq_type
         : _GEN_46 ? _slots_21_io_out_uop_iq_type : _slots_20_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_47
         ? _slots_22_io_out_uop_fu_code
         : _GEN_46 ? _slots_21_io_out_uop_fu_code : _slots_20_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_47
         ? _slots_22_io_out_uop_iw_state
         : _GEN_46 ? _slots_21_io_out_uop_iw_state : _slots_20_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_47
         ? _slots_22_io_out_uop_iw_p1_poisoned
         : _GEN_46
             ? _slots_21_io_out_uop_iw_p1_poisoned
             : _slots_20_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_47
         ? _slots_22_io_out_uop_iw_p2_poisoned
         : _GEN_46
             ? _slots_21_io_out_uop_iw_p2_poisoned
             : _slots_20_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_47
         ? _slots_22_io_out_uop_is_br
         : _GEN_46 ? _slots_21_io_out_uop_is_br : _slots_20_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_47
         ? _slots_22_io_out_uop_is_jalr
         : _GEN_46 ? _slots_21_io_out_uop_is_jalr : _slots_20_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_47
         ? _slots_22_io_out_uop_is_jal
         : _GEN_46 ? _slots_21_io_out_uop_is_jal : _slots_20_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_47
         ? _slots_22_io_out_uop_is_sfb
         : _GEN_46 ? _slots_21_io_out_uop_is_sfb : _slots_20_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_47
         ? _slots_22_io_out_uop_br_mask
         : _GEN_46 ? _slots_21_io_out_uop_br_mask : _slots_20_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_47
         ? _slots_22_io_out_uop_br_tag
         : _GEN_46 ? _slots_21_io_out_uop_br_tag : _slots_20_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_47
         ? _slots_22_io_out_uop_ftq_idx
         : _GEN_46 ? _slots_21_io_out_uop_ftq_idx : _slots_20_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_47
         ? _slots_22_io_out_uop_edge_inst
         : _GEN_46 ? _slots_21_io_out_uop_edge_inst : _slots_20_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_47
         ? _slots_22_io_out_uop_pc_lob
         : _GEN_46 ? _slots_21_io_out_uop_pc_lob : _slots_20_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_47
         ? _slots_22_io_out_uop_taken
         : _GEN_46 ? _slots_21_io_out_uop_taken : _slots_20_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_47
         ? _slots_22_io_out_uop_imm_packed
         : _GEN_46 ? _slots_21_io_out_uop_imm_packed : _slots_20_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_47
         ? _slots_22_io_out_uop_csr_addr
         : _GEN_46 ? _slots_21_io_out_uop_csr_addr : _slots_20_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_47
         ? _slots_22_io_out_uop_rob_idx
         : _GEN_46 ? _slots_21_io_out_uop_rob_idx : _slots_20_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_47
         ? _slots_22_io_out_uop_ldq_idx
         : _GEN_46 ? _slots_21_io_out_uop_ldq_idx : _slots_20_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_47
         ? _slots_22_io_out_uop_stq_idx
         : _GEN_46 ? _slots_21_io_out_uop_stq_idx : _slots_20_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_47
         ? _slots_22_io_out_uop_rxq_idx
         : _GEN_46 ? _slots_21_io_out_uop_rxq_idx : _slots_20_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_47
         ? _slots_22_io_out_uop_pdst
         : _GEN_46 ? _slots_21_io_out_uop_pdst : _slots_20_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_47
         ? _slots_22_io_out_uop_prs1
         : _GEN_46 ? _slots_21_io_out_uop_prs1 : _slots_20_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_47
         ? _slots_22_io_out_uop_prs2
         : _GEN_46 ? _slots_21_io_out_uop_prs2 : _slots_20_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_47
         ? _slots_22_io_out_uop_prs3
         : _GEN_46 ? _slots_21_io_out_uop_prs3 : _slots_20_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_47
         ? _slots_22_io_out_uop_ppred
         : _GEN_46 ? _slots_21_io_out_uop_ppred : _slots_20_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_47
         ? _slots_22_io_out_uop_prs1_busy
         : _GEN_46 ? _slots_21_io_out_uop_prs1_busy : _slots_20_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_47
         ? _slots_22_io_out_uop_prs2_busy
         : _GEN_46 ? _slots_21_io_out_uop_prs2_busy : _slots_20_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_47
         ? _slots_22_io_out_uop_prs3_busy
         : _GEN_46 ? _slots_21_io_out_uop_prs3_busy : _slots_20_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_47
         ? _slots_22_io_out_uop_ppred_busy
         : _GEN_46 ? _slots_21_io_out_uop_ppred_busy : _slots_20_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_47
         ? _slots_22_io_out_uop_stale_pdst
         : _GEN_46 ? _slots_21_io_out_uop_stale_pdst : _slots_20_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_47
         ? _slots_22_io_out_uop_exception
         : _GEN_46 ? _slots_21_io_out_uop_exception : _slots_20_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_47
         ? _slots_22_io_out_uop_exc_cause
         : _GEN_46 ? _slots_21_io_out_uop_exc_cause : _slots_20_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_47
         ? _slots_22_io_out_uop_bypassable
         : _GEN_46 ? _slots_21_io_out_uop_bypassable : _slots_20_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_47
         ? _slots_22_io_out_uop_mem_cmd
         : _GEN_46 ? _slots_21_io_out_uop_mem_cmd : _slots_20_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_47
         ? _slots_22_io_out_uop_mem_size
         : _GEN_46 ? _slots_21_io_out_uop_mem_size : _slots_20_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_47
         ? _slots_22_io_out_uop_mem_signed
         : _GEN_46 ? _slots_21_io_out_uop_mem_signed : _slots_20_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_47
         ? _slots_22_io_out_uop_is_fence
         : _GEN_46 ? _slots_21_io_out_uop_is_fence : _slots_20_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_47
         ? _slots_22_io_out_uop_is_fencei
         : _GEN_46 ? _slots_21_io_out_uop_is_fencei : _slots_20_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_47
         ? _slots_22_io_out_uop_is_amo
         : _GEN_46 ? _slots_21_io_out_uop_is_amo : _slots_20_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_47
         ? _slots_22_io_out_uop_uses_ldq
         : _GEN_46 ? _slots_21_io_out_uop_uses_ldq : _slots_20_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_47
         ? _slots_22_io_out_uop_uses_stq
         : _GEN_46 ? _slots_21_io_out_uop_uses_stq : _slots_20_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_47
         ? _slots_22_io_out_uop_is_sys_pc2epc
         : _GEN_46
             ? _slots_21_io_out_uop_is_sys_pc2epc
             : _slots_20_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_47
         ? _slots_22_io_out_uop_is_unique
         : _GEN_46 ? _slots_21_io_out_uop_is_unique : _slots_20_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_47
         ? _slots_22_io_out_uop_flush_on_commit
         : _GEN_46
             ? _slots_21_io_out_uop_flush_on_commit
             : _slots_20_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_47
         ? _slots_22_io_out_uop_ldst_is_rs1
         : _GEN_46 ? _slots_21_io_out_uop_ldst_is_rs1 : _slots_20_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_47
         ? _slots_22_io_out_uop_ldst
         : _GEN_46 ? _slots_21_io_out_uop_ldst : _slots_20_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_47
         ? _slots_22_io_out_uop_lrs1
         : _GEN_46 ? _slots_21_io_out_uop_lrs1 : _slots_20_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_47
         ? _slots_22_io_out_uop_lrs2
         : _GEN_46 ? _slots_21_io_out_uop_lrs2 : _slots_20_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_47
         ? _slots_22_io_out_uop_lrs3
         : _GEN_46 ? _slots_21_io_out_uop_lrs3 : _slots_20_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_47
         ? _slots_22_io_out_uop_ldst_val
         : _GEN_46 ? _slots_21_io_out_uop_ldst_val : _slots_20_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_47
         ? _slots_22_io_out_uop_dst_rtype
         : _GEN_46 ? _slots_21_io_out_uop_dst_rtype : _slots_20_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_47
         ? _slots_22_io_out_uop_lrs1_rtype
         : _GEN_46 ? _slots_21_io_out_uop_lrs1_rtype : _slots_20_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_47
         ? _slots_22_io_out_uop_lrs2_rtype
         : _GEN_46 ? _slots_21_io_out_uop_lrs2_rtype : _slots_20_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_47
         ? _slots_22_io_out_uop_frs3_en
         : _GEN_46 ? _slots_21_io_out_uop_frs3_en : _slots_20_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_47
         ? _slots_22_io_out_uop_fp_val
         : _GEN_46 ? _slots_21_io_out_uop_fp_val : _slots_20_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_47
         ? _slots_22_io_out_uop_fp_single
         : _GEN_46 ? _slots_21_io_out_uop_fp_single : _slots_20_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_47
         ? _slots_22_io_out_uop_xcpt_pf_if
         : _GEN_46 ? _slots_21_io_out_uop_xcpt_pf_if : _slots_20_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_47
         ? _slots_22_io_out_uop_xcpt_ae_if
         : _GEN_46 ? _slots_21_io_out_uop_xcpt_ae_if : _slots_20_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_47
         ? _slots_22_io_out_uop_xcpt_ma_if
         : _GEN_46 ? _slots_21_io_out_uop_xcpt_ma_if : _slots_20_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_47
         ? _slots_22_io_out_uop_bp_debug_if
         : _GEN_46 ? _slots_21_io_out_uop_bp_debug_if : _slots_20_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_47
         ? _slots_22_io_out_uop_bp_xcpt_if
         : _GEN_46 ? _slots_21_io_out_uop_bp_xcpt_if : _slots_20_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_47
         ? _slots_22_io_out_uop_debug_fsrc
         : _GEN_46 ? _slots_21_io_out_uop_debug_fsrc : _slots_20_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_47
         ? _slots_22_io_out_uop_debug_tsrc
         : _GEN_46 ? _slots_21_io_out_uop_debug_tsrc : _slots_20_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_19_io_valid),
    .io_will_be_valid               (_slots_19_io_will_be_valid),
    .io_request                     (_slots_19_io_request),
    .io_out_uop_uopc                (_slots_19_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_19_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_19_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_19_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_19_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_19_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_19_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_19_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_19_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_19_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_19_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_19_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_19_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_19_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_19_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_19_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_19_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_19_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_19_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_19_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_19_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_19_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_19_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_19_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_19_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_19_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_19_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_19_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_19_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_19_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_19_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_19_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_19_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_19_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_19_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_19_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_19_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_19_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_19_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_19_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_19_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_19_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_19_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_19_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_19_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_19_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_19_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_19_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_19_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_19_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_19_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_19_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_19_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_19_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_19_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_19_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_19_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_19_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_19_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_19_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_19_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_19_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_19_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_19_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_19_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_19_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_19_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_19_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_19_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_19_io_uop_uopc),
    .io_uop_inst                    (_slots_19_io_uop_inst),
    .io_uop_debug_inst              (_slots_19_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_19_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_19_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_19_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_19_io_uop_fu_code),
    .io_uop_iw_state                (_slots_19_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_19_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_19_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_19_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_19_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_19_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_19_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_19_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_19_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_19_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_19_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_19_io_uop_pc_lob),
    .io_uop_taken                   (_slots_19_io_uop_taken),
    .io_uop_imm_packed              (_slots_19_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_19_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_19_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_19_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_19_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_19_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_19_io_uop_pdst),
    .io_uop_prs1                    (_slots_19_io_uop_prs1),
    .io_uop_prs2                    (_slots_19_io_uop_prs2),
    .io_uop_prs3                    (_slots_19_io_uop_prs3),
    .io_uop_ppred                   (_slots_19_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_19_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_19_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_19_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_19_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_19_io_uop_stale_pdst),
    .io_uop_exception               (_slots_19_io_uop_exception),
    .io_uop_exc_cause               (_slots_19_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_19_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_19_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_19_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_19_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_19_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_19_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_19_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_19_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_19_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_19_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_19_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_19_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_19_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_19_io_uop_ldst),
    .io_uop_lrs1                    (_slots_19_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_19_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_19_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_19_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_19_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_19_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_19_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_19_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_19_io_uop_fp_val),
    .io_uop_fp_single               (_slots_19_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_19_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_19_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_19_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_19_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_19_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_19_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_19_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_20 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_20_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_19),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_20_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_49
         ? _slots_23_io_out_uop_uopc
         : _GEN_48 ? _slots_22_io_out_uop_uopc : _slots_21_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_49
         ? _slots_23_io_out_uop_inst
         : _GEN_48 ? _slots_22_io_out_uop_inst : _slots_21_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_49
         ? _slots_23_io_out_uop_debug_inst
         : _GEN_48 ? _slots_22_io_out_uop_debug_inst : _slots_21_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_49
         ? _slots_23_io_out_uop_is_rvc
         : _GEN_48 ? _slots_22_io_out_uop_is_rvc : _slots_21_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_49
         ? _slots_23_io_out_uop_debug_pc
         : _GEN_48 ? _slots_22_io_out_uop_debug_pc : _slots_21_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_49
         ? _slots_23_io_out_uop_iq_type
         : _GEN_48 ? _slots_22_io_out_uop_iq_type : _slots_21_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_49
         ? _slots_23_io_out_uop_fu_code
         : _GEN_48 ? _slots_22_io_out_uop_fu_code : _slots_21_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_49
         ? _slots_23_io_out_uop_iw_state
         : _GEN_48 ? _slots_22_io_out_uop_iw_state : _slots_21_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_49
         ? _slots_23_io_out_uop_iw_p1_poisoned
         : _GEN_48
             ? _slots_22_io_out_uop_iw_p1_poisoned
             : _slots_21_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_49
         ? _slots_23_io_out_uop_iw_p2_poisoned
         : _GEN_48
             ? _slots_22_io_out_uop_iw_p2_poisoned
             : _slots_21_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_49
         ? _slots_23_io_out_uop_is_br
         : _GEN_48 ? _slots_22_io_out_uop_is_br : _slots_21_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_49
         ? _slots_23_io_out_uop_is_jalr
         : _GEN_48 ? _slots_22_io_out_uop_is_jalr : _slots_21_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_49
         ? _slots_23_io_out_uop_is_jal
         : _GEN_48 ? _slots_22_io_out_uop_is_jal : _slots_21_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_49
         ? _slots_23_io_out_uop_is_sfb
         : _GEN_48 ? _slots_22_io_out_uop_is_sfb : _slots_21_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_49
         ? _slots_23_io_out_uop_br_mask
         : _GEN_48 ? _slots_22_io_out_uop_br_mask : _slots_21_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_49
         ? _slots_23_io_out_uop_br_tag
         : _GEN_48 ? _slots_22_io_out_uop_br_tag : _slots_21_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_49
         ? _slots_23_io_out_uop_ftq_idx
         : _GEN_48 ? _slots_22_io_out_uop_ftq_idx : _slots_21_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_49
         ? _slots_23_io_out_uop_edge_inst
         : _GEN_48 ? _slots_22_io_out_uop_edge_inst : _slots_21_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_49
         ? _slots_23_io_out_uop_pc_lob
         : _GEN_48 ? _slots_22_io_out_uop_pc_lob : _slots_21_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_49
         ? _slots_23_io_out_uop_taken
         : _GEN_48 ? _slots_22_io_out_uop_taken : _slots_21_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_49
         ? _slots_23_io_out_uop_imm_packed
         : _GEN_48 ? _slots_22_io_out_uop_imm_packed : _slots_21_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_49
         ? _slots_23_io_out_uop_csr_addr
         : _GEN_48 ? _slots_22_io_out_uop_csr_addr : _slots_21_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_49
         ? _slots_23_io_out_uop_rob_idx
         : _GEN_48 ? _slots_22_io_out_uop_rob_idx : _slots_21_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_49
         ? _slots_23_io_out_uop_ldq_idx
         : _GEN_48 ? _slots_22_io_out_uop_ldq_idx : _slots_21_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_49
         ? _slots_23_io_out_uop_stq_idx
         : _GEN_48 ? _slots_22_io_out_uop_stq_idx : _slots_21_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_49
         ? _slots_23_io_out_uop_rxq_idx
         : _GEN_48 ? _slots_22_io_out_uop_rxq_idx : _slots_21_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_49
         ? _slots_23_io_out_uop_pdst
         : _GEN_48 ? _slots_22_io_out_uop_pdst : _slots_21_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_49
         ? _slots_23_io_out_uop_prs1
         : _GEN_48 ? _slots_22_io_out_uop_prs1 : _slots_21_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_49
         ? _slots_23_io_out_uop_prs2
         : _GEN_48 ? _slots_22_io_out_uop_prs2 : _slots_21_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_49
         ? _slots_23_io_out_uop_prs3
         : _GEN_48 ? _slots_22_io_out_uop_prs3 : _slots_21_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_49
         ? _slots_23_io_out_uop_ppred
         : _GEN_48 ? _slots_22_io_out_uop_ppred : _slots_21_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_49
         ? _slots_23_io_out_uop_prs1_busy
         : _GEN_48 ? _slots_22_io_out_uop_prs1_busy : _slots_21_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_49
         ? _slots_23_io_out_uop_prs2_busy
         : _GEN_48 ? _slots_22_io_out_uop_prs2_busy : _slots_21_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_49
         ? _slots_23_io_out_uop_prs3_busy
         : _GEN_48 ? _slots_22_io_out_uop_prs3_busy : _slots_21_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_49
         ? _slots_23_io_out_uop_ppred_busy
         : _GEN_48 ? _slots_22_io_out_uop_ppred_busy : _slots_21_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_49
         ? _slots_23_io_out_uop_stale_pdst
         : _GEN_48 ? _slots_22_io_out_uop_stale_pdst : _slots_21_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_49
         ? _slots_23_io_out_uop_exception
         : _GEN_48 ? _slots_22_io_out_uop_exception : _slots_21_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_49
         ? _slots_23_io_out_uop_exc_cause
         : _GEN_48 ? _slots_22_io_out_uop_exc_cause : _slots_21_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_49
         ? _slots_23_io_out_uop_bypassable
         : _GEN_48 ? _slots_22_io_out_uop_bypassable : _slots_21_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_49
         ? _slots_23_io_out_uop_mem_cmd
         : _GEN_48 ? _slots_22_io_out_uop_mem_cmd : _slots_21_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_49
         ? _slots_23_io_out_uop_mem_size
         : _GEN_48 ? _slots_22_io_out_uop_mem_size : _slots_21_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_49
         ? _slots_23_io_out_uop_mem_signed
         : _GEN_48 ? _slots_22_io_out_uop_mem_signed : _slots_21_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_49
         ? _slots_23_io_out_uop_is_fence
         : _GEN_48 ? _slots_22_io_out_uop_is_fence : _slots_21_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_49
         ? _slots_23_io_out_uop_is_fencei
         : _GEN_48 ? _slots_22_io_out_uop_is_fencei : _slots_21_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_49
         ? _slots_23_io_out_uop_is_amo
         : _GEN_48 ? _slots_22_io_out_uop_is_amo : _slots_21_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_49
         ? _slots_23_io_out_uop_uses_ldq
         : _GEN_48 ? _slots_22_io_out_uop_uses_ldq : _slots_21_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_49
         ? _slots_23_io_out_uop_uses_stq
         : _GEN_48 ? _slots_22_io_out_uop_uses_stq : _slots_21_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_49
         ? _slots_23_io_out_uop_is_sys_pc2epc
         : _GEN_48
             ? _slots_22_io_out_uop_is_sys_pc2epc
             : _slots_21_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_49
         ? _slots_23_io_out_uop_is_unique
         : _GEN_48 ? _slots_22_io_out_uop_is_unique : _slots_21_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_49
         ? _slots_23_io_out_uop_flush_on_commit
         : _GEN_48
             ? _slots_22_io_out_uop_flush_on_commit
             : _slots_21_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_49
         ? _slots_23_io_out_uop_ldst_is_rs1
         : _GEN_48 ? _slots_22_io_out_uop_ldst_is_rs1 : _slots_21_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_49
         ? _slots_23_io_out_uop_ldst
         : _GEN_48 ? _slots_22_io_out_uop_ldst : _slots_21_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_49
         ? _slots_23_io_out_uop_lrs1
         : _GEN_48 ? _slots_22_io_out_uop_lrs1 : _slots_21_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_49
         ? _slots_23_io_out_uop_lrs2
         : _GEN_48 ? _slots_22_io_out_uop_lrs2 : _slots_21_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_49
         ? _slots_23_io_out_uop_lrs3
         : _GEN_48 ? _slots_22_io_out_uop_lrs3 : _slots_21_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_49
         ? _slots_23_io_out_uop_ldst_val
         : _GEN_48 ? _slots_22_io_out_uop_ldst_val : _slots_21_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_49
         ? _slots_23_io_out_uop_dst_rtype
         : _GEN_48 ? _slots_22_io_out_uop_dst_rtype : _slots_21_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_49
         ? _slots_23_io_out_uop_lrs1_rtype
         : _GEN_48 ? _slots_22_io_out_uop_lrs1_rtype : _slots_21_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_49
         ? _slots_23_io_out_uop_lrs2_rtype
         : _GEN_48 ? _slots_22_io_out_uop_lrs2_rtype : _slots_21_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_49
         ? _slots_23_io_out_uop_frs3_en
         : _GEN_48 ? _slots_22_io_out_uop_frs3_en : _slots_21_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_49
         ? _slots_23_io_out_uop_fp_val
         : _GEN_48 ? _slots_22_io_out_uop_fp_val : _slots_21_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_49
         ? _slots_23_io_out_uop_fp_single
         : _GEN_48 ? _slots_22_io_out_uop_fp_single : _slots_21_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_49
         ? _slots_23_io_out_uop_xcpt_pf_if
         : _GEN_48 ? _slots_22_io_out_uop_xcpt_pf_if : _slots_21_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_49
         ? _slots_23_io_out_uop_xcpt_ae_if
         : _GEN_48 ? _slots_22_io_out_uop_xcpt_ae_if : _slots_21_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_49
         ? _slots_23_io_out_uop_xcpt_ma_if
         : _GEN_48 ? _slots_22_io_out_uop_xcpt_ma_if : _slots_21_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_49
         ? _slots_23_io_out_uop_bp_debug_if
         : _GEN_48 ? _slots_22_io_out_uop_bp_debug_if : _slots_21_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_49
         ? _slots_23_io_out_uop_bp_xcpt_if
         : _GEN_48 ? _slots_22_io_out_uop_bp_xcpt_if : _slots_21_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_49
         ? _slots_23_io_out_uop_debug_fsrc
         : _GEN_48 ? _slots_22_io_out_uop_debug_fsrc : _slots_21_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_49
         ? _slots_23_io_out_uop_debug_tsrc
         : _GEN_48 ? _slots_22_io_out_uop_debug_tsrc : _slots_21_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_20_io_valid),
    .io_will_be_valid               (_slots_20_io_will_be_valid),
    .io_request                     (_slots_20_io_request),
    .io_out_uop_uopc                (_slots_20_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_20_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_20_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_20_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_20_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_20_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_20_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_20_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_20_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_20_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_20_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_20_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_20_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_20_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_20_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_20_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_20_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_20_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_20_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_20_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_20_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_20_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_20_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_20_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_20_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_20_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_20_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_20_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_20_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_20_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_20_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_20_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_20_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_20_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_20_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_20_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_20_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_20_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_20_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_20_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_20_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_20_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_20_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_20_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_20_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_20_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_20_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_20_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_20_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_20_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_20_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_20_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_20_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_20_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_20_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_20_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_20_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_20_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_20_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_20_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_20_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_20_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_20_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_20_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_20_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_20_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_20_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_20_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_20_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_20_io_uop_uopc),
    .io_uop_inst                    (_slots_20_io_uop_inst),
    .io_uop_debug_inst              (_slots_20_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_20_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_20_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_20_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_20_io_uop_fu_code),
    .io_uop_iw_state                (_slots_20_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_20_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_20_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_20_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_20_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_20_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_20_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_20_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_20_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_20_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_20_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_20_io_uop_pc_lob),
    .io_uop_taken                   (_slots_20_io_uop_taken),
    .io_uop_imm_packed              (_slots_20_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_20_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_20_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_20_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_20_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_20_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_20_io_uop_pdst),
    .io_uop_prs1                    (_slots_20_io_uop_prs1),
    .io_uop_prs2                    (_slots_20_io_uop_prs2),
    .io_uop_prs3                    (_slots_20_io_uop_prs3),
    .io_uop_ppred                   (_slots_20_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_20_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_20_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_20_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_20_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_20_io_uop_stale_pdst),
    .io_uop_exception               (_slots_20_io_uop_exception),
    .io_uop_exc_cause               (_slots_20_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_20_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_20_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_20_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_20_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_20_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_20_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_20_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_20_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_20_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_20_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_20_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_20_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_20_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_20_io_uop_ldst),
    .io_uop_lrs1                    (_slots_20_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_20_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_20_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_20_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_20_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_20_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_20_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_20_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_20_io_uop_fp_val),
    .io_uop_fp_single               (_slots_20_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_20_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_20_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_20_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_20_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_20_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_20_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_20_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_21 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_21_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_20),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_21_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_51
         ? _slots_24_io_out_uop_uopc
         : _GEN_50 ? _slots_23_io_out_uop_uopc : _slots_22_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_51
         ? _slots_24_io_out_uop_inst
         : _GEN_50 ? _slots_23_io_out_uop_inst : _slots_22_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_51
         ? _slots_24_io_out_uop_debug_inst
         : _GEN_50 ? _slots_23_io_out_uop_debug_inst : _slots_22_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_51
         ? _slots_24_io_out_uop_is_rvc
         : _GEN_50 ? _slots_23_io_out_uop_is_rvc : _slots_22_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_51
         ? _slots_24_io_out_uop_debug_pc
         : _GEN_50 ? _slots_23_io_out_uop_debug_pc : _slots_22_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_51
         ? _slots_24_io_out_uop_iq_type
         : _GEN_50 ? _slots_23_io_out_uop_iq_type : _slots_22_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_51
         ? _slots_24_io_out_uop_fu_code
         : _GEN_50 ? _slots_23_io_out_uop_fu_code : _slots_22_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_51
         ? _slots_24_io_out_uop_iw_state
         : _GEN_50 ? _slots_23_io_out_uop_iw_state : _slots_22_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_51
         ? _slots_24_io_out_uop_iw_p1_poisoned
         : _GEN_50
             ? _slots_23_io_out_uop_iw_p1_poisoned
             : _slots_22_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_51
         ? _slots_24_io_out_uop_iw_p2_poisoned
         : _GEN_50
             ? _slots_23_io_out_uop_iw_p2_poisoned
             : _slots_22_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_51
         ? _slots_24_io_out_uop_is_br
         : _GEN_50 ? _slots_23_io_out_uop_is_br : _slots_22_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_51
         ? _slots_24_io_out_uop_is_jalr
         : _GEN_50 ? _slots_23_io_out_uop_is_jalr : _slots_22_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_51
         ? _slots_24_io_out_uop_is_jal
         : _GEN_50 ? _slots_23_io_out_uop_is_jal : _slots_22_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_51
         ? _slots_24_io_out_uop_is_sfb
         : _GEN_50 ? _slots_23_io_out_uop_is_sfb : _slots_22_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_51
         ? _slots_24_io_out_uop_br_mask
         : _GEN_50 ? _slots_23_io_out_uop_br_mask : _slots_22_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_51
         ? _slots_24_io_out_uop_br_tag
         : _GEN_50 ? _slots_23_io_out_uop_br_tag : _slots_22_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_51
         ? _slots_24_io_out_uop_ftq_idx
         : _GEN_50 ? _slots_23_io_out_uop_ftq_idx : _slots_22_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_51
         ? _slots_24_io_out_uop_edge_inst
         : _GEN_50 ? _slots_23_io_out_uop_edge_inst : _slots_22_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_51
         ? _slots_24_io_out_uop_pc_lob
         : _GEN_50 ? _slots_23_io_out_uop_pc_lob : _slots_22_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_51
         ? _slots_24_io_out_uop_taken
         : _GEN_50 ? _slots_23_io_out_uop_taken : _slots_22_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_51
         ? _slots_24_io_out_uop_imm_packed
         : _GEN_50 ? _slots_23_io_out_uop_imm_packed : _slots_22_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_51
         ? _slots_24_io_out_uop_csr_addr
         : _GEN_50 ? _slots_23_io_out_uop_csr_addr : _slots_22_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_51
         ? _slots_24_io_out_uop_rob_idx
         : _GEN_50 ? _slots_23_io_out_uop_rob_idx : _slots_22_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_51
         ? _slots_24_io_out_uop_ldq_idx
         : _GEN_50 ? _slots_23_io_out_uop_ldq_idx : _slots_22_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_51
         ? _slots_24_io_out_uop_stq_idx
         : _GEN_50 ? _slots_23_io_out_uop_stq_idx : _slots_22_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_51
         ? _slots_24_io_out_uop_rxq_idx
         : _GEN_50 ? _slots_23_io_out_uop_rxq_idx : _slots_22_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_51
         ? _slots_24_io_out_uop_pdst
         : _GEN_50 ? _slots_23_io_out_uop_pdst : _slots_22_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_51
         ? _slots_24_io_out_uop_prs1
         : _GEN_50 ? _slots_23_io_out_uop_prs1 : _slots_22_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_51
         ? _slots_24_io_out_uop_prs2
         : _GEN_50 ? _slots_23_io_out_uop_prs2 : _slots_22_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_51
         ? _slots_24_io_out_uop_prs3
         : _GEN_50 ? _slots_23_io_out_uop_prs3 : _slots_22_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_51
         ? _slots_24_io_out_uop_ppred
         : _GEN_50 ? _slots_23_io_out_uop_ppred : _slots_22_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_51
         ? _slots_24_io_out_uop_prs1_busy
         : _GEN_50 ? _slots_23_io_out_uop_prs1_busy : _slots_22_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_51
         ? _slots_24_io_out_uop_prs2_busy
         : _GEN_50 ? _slots_23_io_out_uop_prs2_busy : _slots_22_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_51
         ? _slots_24_io_out_uop_prs3_busy
         : _GEN_50 ? _slots_23_io_out_uop_prs3_busy : _slots_22_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_51
         ? _slots_24_io_out_uop_ppred_busy
         : _GEN_50 ? _slots_23_io_out_uop_ppred_busy : _slots_22_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_51
         ? _slots_24_io_out_uop_stale_pdst
         : _GEN_50 ? _slots_23_io_out_uop_stale_pdst : _slots_22_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_51
         ? _slots_24_io_out_uop_exception
         : _GEN_50 ? _slots_23_io_out_uop_exception : _slots_22_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_51
         ? _slots_24_io_out_uop_exc_cause
         : _GEN_50 ? _slots_23_io_out_uop_exc_cause : _slots_22_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_51
         ? _slots_24_io_out_uop_bypassable
         : _GEN_50 ? _slots_23_io_out_uop_bypassable : _slots_22_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_51
         ? _slots_24_io_out_uop_mem_cmd
         : _GEN_50 ? _slots_23_io_out_uop_mem_cmd : _slots_22_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_51
         ? _slots_24_io_out_uop_mem_size
         : _GEN_50 ? _slots_23_io_out_uop_mem_size : _slots_22_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_51
         ? _slots_24_io_out_uop_mem_signed
         : _GEN_50 ? _slots_23_io_out_uop_mem_signed : _slots_22_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_51
         ? _slots_24_io_out_uop_is_fence
         : _GEN_50 ? _slots_23_io_out_uop_is_fence : _slots_22_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_51
         ? _slots_24_io_out_uop_is_fencei
         : _GEN_50 ? _slots_23_io_out_uop_is_fencei : _slots_22_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_51
         ? _slots_24_io_out_uop_is_amo
         : _GEN_50 ? _slots_23_io_out_uop_is_amo : _slots_22_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_51
         ? _slots_24_io_out_uop_uses_ldq
         : _GEN_50 ? _slots_23_io_out_uop_uses_ldq : _slots_22_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_51
         ? _slots_24_io_out_uop_uses_stq
         : _GEN_50 ? _slots_23_io_out_uop_uses_stq : _slots_22_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_51
         ? _slots_24_io_out_uop_is_sys_pc2epc
         : _GEN_50
             ? _slots_23_io_out_uop_is_sys_pc2epc
             : _slots_22_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_51
         ? _slots_24_io_out_uop_is_unique
         : _GEN_50 ? _slots_23_io_out_uop_is_unique : _slots_22_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_51
         ? _slots_24_io_out_uop_flush_on_commit
         : _GEN_50
             ? _slots_23_io_out_uop_flush_on_commit
             : _slots_22_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_51
         ? _slots_24_io_out_uop_ldst_is_rs1
         : _GEN_50 ? _slots_23_io_out_uop_ldst_is_rs1 : _slots_22_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_51
         ? _slots_24_io_out_uop_ldst
         : _GEN_50 ? _slots_23_io_out_uop_ldst : _slots_22_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_51
         ? _slots_24_io_out_uop_lrs1
         : _GEN_50 ? _slots_23_io_out_uop_lrs1 : _slots_22_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_51
         ? _slots_24_io_out_uop_lrs2
         : _GEN_50 ? _slots_23_io_out_uop_lrs2 : _slots_22_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_51
         ? _slots_24_io_out_uop_lrs3
         : _GEN_50 ? _slots_23_io_out_uop_lrs3 : _slots_22_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_51
         ? _slots_24_io_out_uop_ldst_val
         : _GEN_50 ? _slots_23_io_out_uop_ldst_val : _slots_22_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_51
         ? _slots_24_io_out_uop_dst_rtype
         : _GEN_50 ? _slots_23_io_out_uop_dst_rtype : _slots_22_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_51
         ? _slots_24_io_out_uop_lrs1_rtype
         : _GEN_50 ? _slots_23_io_out_uop_lrs1_rtype : _slots_22_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_51
         ? _slots_24_io_out_uop_lrs2_rtype
         : _GEN_50 ? _slots_23_io_out_uop_lrs2_rtype : _slots_22_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_51
         ? _slots_24_io_out_uop_frs3_en
         : _GEN_50 ? _slots_23_io_out_uop_frs3_en : _slots_22_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_51
         ? _slots_24_io_out_uop_fp_val
         : _GEN_50 ? _slots_23_io_out_uop_fp_val : _slots_22_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_51
         ? _slots_24_io_out_uop_fp_single
         : _GEN_50 ? _slots_23_io_out_uop_fp_single : _slots_22_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_51
         ? _slots_24_io_out_uop_xcpt_pf_if
         : _GEN_50 ? _slots_23_io_out_uop_xcpt_pf_if : _slots_22_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_51
         ? _slots_24_io_out_uop_xcpt_ae_if
         : _GEN_50 ? _slots_23_io_out_uop_xcpt_ae_if : _slots_22_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_51
         ? _slots_24_io_out_uop_xcpt_ma_if
         : _GEN_50 ? _slots_23_io_out_uop_xcpt_ma_if : _slots_22_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_51
         ? _slots_24_io_out_uop_bp_debug_if
         : _GEN_50 ? _slots_23_io_out_uop_bp_debug_if : _slots_22_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_51
         ? _slots_24_io_out_uop_bp_xcpt_if
         : _GEN_50 ? _slots_23_io_out_uop_bp_xcpt_if : _slots_22_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_51
         ? _slots_24_io_out_uop_debug_fsrc
         : _GEN_50 ? _slots_23_io_out_uop_debug_fsrc : _slots_22_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_51
         ? _slots_24_io_out_uop_debug_tsrc
         : _GEN_50 ? _slots_23_io_out_uop_debug_tsrc : _slots_22_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_21_io_valid),
    .io_will_be_valid               (_slots_21_io_will_be_valid),
    .io_request                     (_slots_21_io_request),
    .io_out_uop_uopc                (_slots_21_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_21_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_21_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_21_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_21_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_21_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_21_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_21_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_21_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_21_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_21_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_21_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_21_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_21_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_21_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_21_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_21_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_21_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_21_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_21_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_21_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_21_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_21_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_21_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_21_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_21_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_21_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_21_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_21_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_21_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_21_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_21_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_21_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_21_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_21_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_21_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_21_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_21_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_21_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_21_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_21_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_21_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_21_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_21_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_21_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_21_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_21_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_21_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_21_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_21_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_21_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_21_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_21_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_21_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_21_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_21_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_21_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_21_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_21_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_21_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_21_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_21_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_21_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_21_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_21_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_21_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_21_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_21_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_21_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_21_io_uop_uopc),
    .io_uop_inst                    (_slots_21_io_uop_inst),
    .io_uop_debug_inst              (_slots_21_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_21_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_21_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_21_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_21_io_uop_fu_code),
    .io_uop_iw_state                (_slots_21_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_21_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_21_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_21_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_21_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_21_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_21_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_21_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_21_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_21_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_21_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_21_io_uop_pc_lob),
    .io_uop_taken                   (_slots_21_io_uop_taken),
    .io_uop_imm_packed              (_slots_21_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_21_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_21_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_21_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_21_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_21_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_21_io_uop_pdst),
    .io_uop_prs1                    (_slots_21_io_uop_prs1),
    .io_uop_prs2                    (_slots_21_io_uop_prs2),
    .io_uop_prs3                    (_slots_21_io_uop_prs3),
    .io_uop_ppred                   (_slots_21_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_21_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_21_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_21_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_21_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_21_io_uop_stale_pdst),
    .io_uop_exception               (_slots_21_io_uop_exception),
    .io_uop_exc_cause               (_slots_21_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_21_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_21_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_21_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_21_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_21_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_21_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_21_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_21_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_21_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_21_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_21_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_21_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_21_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_21_io_uop_ldst),
    .io_uop_lrs1                    (_slots_21_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_21_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_21_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_21_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_21_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_21_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_21_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_21_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_21_io_uop_fp_val),
    .io_uop_fp_single               (_slots_21_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_21_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_21_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_21_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_21_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_21_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_21_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_21_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_22 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_22_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_21),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_22_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_53
         ? _slots_25_io_out_uop_uopc
         : _GEN_52 ? _slots_24_io_out_uop_uopc : _slots_23_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_53
         ? _slots_25_io_out_uop_inst
         : _GEN_52 ? _slots_24_io_out_uop_inst : _slots_23_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_53
         ? _slots_25_io_out_uop_debug_inst
         : _GEN_52 ? _slots_24_io_out_uop_debug_inst : _slots_23_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_53
         ? _slots_25_io_out_uop_is_rvc
         : _GEN_52 ? _slots_24_io_out_uop_is_rvc : _slots_23_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_53
         ? _slots_25_io_out_uop_debug_pc
         : _GEN_52 ? _slots_24_io_out_uop_debug_pc : _slots_23_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_53
         ? _slots_25_io_out_uop_iq_type
         : _GEN_52 ? _slots_24_io_out_uop_iq_type : _slots_23_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_53
         ? _slots_25_io_out_uop_fu_code
         : _GEN_52 ? _slots_24_io_out_uop_fu_code : _slots_23_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_53
         ? _slots_25_io_out_uop_iw_state
         : _GEN_52 ? _slots_24_io_out_uop_iw_state : _slots_23_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_53
         ? _slots_25_io_out_uop_iw_p1_poisoned
         : _GEN_52
             ? _slots_24_io_out_uop_iw_p1_poisoned
             : _slots_23_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_53
         ? _slots_25_io_out_uop_iw_p2_poisoned
         : _GEN_52
             ? _slots_24_io_out_uop_iw_p2_poisoned
             : _slots_23_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_53
         ? _slots_25_io_out_uop_is_br
         : _GEN_52 ? _slots_24_io_out_uop_is_br : _slots_23_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_53
         ? _slots_25_io_out_uop_is_jalr
         : _GEN_52 ? _slots_24_io_out_uop_is_jalr : _slots_23_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_53
         ? _slots_25_io_out_uop_is_jal
         : _GEN_52 ? _slots_24_io_out_uop_is_jal : _slots_23_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_53
         ? _slots_25_io_out_uop_is_sfb
         : _GEN_52 ? _slots_24_io_out_uop_is_sfb : _slots_23_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_53
         ? _slots_25_io_out_uop_br_mask
         : _GEN_52 ? _slots_24_io_out_uop_br_mask : _slots_23_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_53
         ? _slots_25_io_out_uop_br_tag
         : _GEN_52 ? _slots_24_io_out_uop_br_tag : _slots_23_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_53
         ? _slots_25_io_out_uop_ftq_idx
         : _GEN_52 ? _slots_24_io_out_uop_ftq_idx : _slots_23_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_53
         ? _slots_25_io_out_uop_edge_inst
         : _GEN_52 ? _slots_24_io_out_uop_edge_inst : _slots_23_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_53
         ? _slots_25_io_out_uop_pc_lob
         : _GEN_52 ? _slots_24_io_out_uop_pc_lob : _slots_23_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_53
         ? _slots_25_io_out_uop_taken
         : _GEN_52 ? _slots_24_io_out_uop_taken : _slots_23_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_53
         ? _slots_25_io_out_uop_imm_packed
         : _GEN_52 ? _slots_24_io_out_uop_imm_packed : _slots_23_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_53
         ? _slots_25_io_out_uop_csr_addr
         : _GEN_52 ? _slots_24_io_out_uop_csr_addr : _slots_23_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_53
         ? _slots_25_io_out_uop_rob_idx
         : _GEN_52 ? _slots_24_io_out_uop_rob_idx : _slots_23_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_53
         ? _slots_25_io_out_uop_ldq_idx
         : _GEN_52 ? _slots_24_io_out_uop_ldq_idx : _slots_23_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_53
         ? _slots_25_io_out_uop_stq_idx
         : _GEN_52 ? _slots_24_io_out_uop_stq_idx : _slots_23_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_53
         ? _slots_25_io_out_uop_rxq_idx
         : _GEN_52 ? _slots_24_io_out_uop_rxq_idx : _slots_23_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_53
         ? _slots_25_io_out_uop_pdst
         : _GEN_52 ? _slots_24_io_out_uop_pdst : _slots_23_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_53
         ? _slots_25_io_out_uop_prs1
         : _GEN_52 ? _slots_24_io_out_uop_prs1 : _slots_23_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_53
         ? _slots_25_io_out_uop_prs2
         : _GEN_52 ? _slots_24_io_out_uop_prs2 : _slots_23_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_53
         ? _slots_25_io_out_uop_prs3
         : _GEN_52 ? _slots_24_io_out_uop_prs3 : _slots_23_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_53
         ? _slots_25_io_out_uop_ppred
         : _GEN_52 ? _slots_24_io_out_uop_ppred : _slots_23_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_53
         ? _slots_25_io_out_uop_prs1_busy
         : _GEN_52 ? _slots_24_io_out_uop_prs1_busy : _slots_23_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_53
         ? _slots_25_io_out_uop_prs2_busy
         : _GEN_52 ? _slots_24_io_out_uop_prs2_busy : _slots_23_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_53
         ? _slots_25_io_out_uop_prs3_busy
         : _GEN_52 ? _slots_24_io_out_uop_prs3_busy : _slots_23_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_53
         ? _slots_25_io_out_uop_ppred_busy
         : _GEN_52 ? _slots_24_io_out_uop_ppred_busy : _slots_23_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_53
         ? _slots_25_io_out_uop_stale_pdst
         : _GEN_52 ? _slots_24_io_out_uop_stale_pdst : _slots_23_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_53
         ? _slots_25_io_out_uop_exception
         : _GEN_52 ? _slots_24_io_out_uop_exception : _slots_23_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_53
         ? _slots_25_io_out_uop_exc_cause
         : _GEN_52 ? _slots_24_io_out_uop_exc_cause : _slots_23_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_53
         ? _slots_25_io_out_uop_bypassable
         : _GEN_52 ? _slots_24_io_out_uop_bypassable : _slots_23_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_53
         ? _slots_25_io_out_uop_mem_cmd
         : _GEN_52 ? _slots_24_io_out_uop_mem_cmd : _slots_23_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_53
         ? _slots_25_io_out_uop_mem_size
         : _GEN_52 ? _slots_24_io_out_uop_mem_size : _slots_23_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_53
         ? _slots_25_io_out_uop_mem_signed
         : _GEN_52 ? _slots_24_io_out_uop_mem_signed : _slots_23_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_53
         ? _slots_25_io_out_uop_is_fence
         : _GEN_52 ? _slots_24_io_out_uop_is_fence : _slots_23_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_53
         ? _slots_25_io_out_uop_is_fencei
         : _GEN_52 ? _slots_24_io_out_uop_is_fencei : _slots_23_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_53
         ? _slots_25_io_out_uop_is_amo
         : _GEN_52 ? _slots_24_io_out_uop_is_amo : _slots_23_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_53
         ? _slots_25_io_out_uop_uses_ldq
         : _GEN_52 ? _slots_24_io_out_uop_uses_ldq : _slots_23_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_53
         ? _slots_25_io_out_uop_uses_stq
         : _GEN_52 ? _slots_24_io_out_uop_uses_stq : _slots_23_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_53
         ? _slots_25_io_out_uop_is_sys_pc2epc
         : _GEN_52
             ? _slots_24_io_out_uop_is_sys_pc2epc
             : _slots_23_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_53
         ? _slots_25_io_out_uop_is_unique
         : _GEN_52 ? _slots_24_io_out_uop_is_unique : _slots_23_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_53
         ? _slots_25_io_out_uop_flush_on_commit
         : _GEN_52
             ? _slots_24_io_out_uop_flush_on_commit
             : _slots_23_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_53
         ? _slots_25_io_out_uop_ldst_is_rs1
         : _GEN_52 ? _slots_24_io_out_uop_ldst_is_rs1 : _slots_23_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_53
         ? _slots_25_io_out_uop_ldst
         : _GEN_52 ? _slots_24_io_out_uop_ldst : _slots_23_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_53
         ? _slots_25_io_out_uop_lrs1
         : _GEN_52 ? _slots_24_io_out_uop_lrs1 : _slots_23_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_53
         ? _slots_25_io_out_uop_lrs2
         : _GEN_52 ? _slots_24_io_out_uop_lrs2 : _slots_23_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_53
         ? _slots_25_io_out_uop_lrs3
         : _GEN_52 ? _slots_24_io_out_uop_lrs3 : _slots_23_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_53
         ? _slots_25_io_out_uop_ldst_val
         : _GEN_52 ? _slots_24_io_out_uop_ldst_val : _slots_23_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_53
         ? _slots_25_io_out_uop_dst_rtype
         : _GEN_52 ? _slots_24_io_out_uop_dst_rtype : _slots_23_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_53
         ? _slots_25_io_out_uop_lrs1_rtype
         : _GEN_52 ? _slots_24_io_out_uop_lrs1_rtype : _slots_23_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_53
         ? _slots_25_io_out_uop_lrs2_rtype
         : _GEN_52 ? _slots_24_io_out_uop_lrs2_rtype : _slots_23_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_53
         ? _slots_25_io_out_uop_frs3_en
         : _GEN_52 ? _slots_24_io_out_uop_frs3_en : _slots_23_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_53
         ? _slots_25_io_out_uop_fp_val
         : _GEN_52 ? _slots_24_io_out_uop_fp_val : _slots_23_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_53
         ? _slots_25_io_out_uop_fp_single
         : _GEN_52 ? _slots_24_io_out_uop_fp_single : _slots_23_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_53
         ? _slots_25_io_out_uop_xcpt_pf_if
         : _GEN_52 ? _slots_24_io_out_uop_xcpt_pf_if : _slots_23_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_53
         ? _slots_25_io_out_uop_xcpt_ae_if
         : _GEN_52 ? _slots_24_io_out_uop_xcpt_ae_if : _slots_23_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_53
         ? _slots_25_io_out_uop_xcpt_ma_if
         : _GEN_52 ? _slots_24_io_out_uop_xcpt_ma_if : _slots_23_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_53
         ? _slots_25_io_out_uop_bp_debug_if
         : _GEN_52 ? _slots_24_io_out_uop_bp_debug_if : _slots_23_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_53
         ? _slots_25_io_out_uop_bp_xcpt_if
         : _GEN_52 ? _slots_24_io_out_uop_bp_xcpt_if : _slots_23_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_53
         ? _slots_25_io_out_uop_debug_fsrc
         : _GEN_52 ? _slots_24_io_out_uop_debug_fsrc : _slots_23_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_53
         ? _slots_25_io_out_uop_debug_tsrc
         : _GEN_52 ? _slots_24_io_out_uop_debug_tsrc : _slots_23_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_22_io_valid),
    .io_will_be_valid               (_slots_22_io_will_be_valid),
    .io_request                     (_slots_22_io_request),
    .io_out_uop_uopc                (_slots_22_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_22_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_22_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_22_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_22_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_22_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_22_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_22_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_22_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_22_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_22_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_22_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_22_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_22_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_22_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_22_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_22_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_22_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_22_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_22_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_22_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_22_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_22_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_22_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_22_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_22_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_22_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_22_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_22_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_22_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_22_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_22_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_22_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_22_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_22_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_22_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_22_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_22_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_22_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_22_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_22_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_22_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_22_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_22_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_22_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_22_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_22_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_22_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_22_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_22_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_22_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_22_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_22_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_22_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_22_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_22_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_22_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_22_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_22_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_22_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_22_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_22_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_22_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_22_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_22_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_22_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_22_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_22_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_22_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_22_io_uop_uopc),
    .io_uop_inst                    (_slots_22_io_uop_inst),
    .io_uop_debug_inst              (_slots_22_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_22_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_22_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_22_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_22_io_uop_fu_code),
    .io_uop_iw_state                (_slots_22_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_22_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_22_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_22_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_22_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_22_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_22_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_22_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_22_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_22_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_22_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_22_io_uop_pc_lob),
    .io_uop_taken                   (_slots_22_io_uop_taken),
    .io_uop_imm_packed              (_slots_22_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_22_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_22_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_22_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_22_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_22_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_22_io_uop_pdst),
    .io_uop_prs1                    (_slots_22_io_uop_prs1),
    .io_uop_prs2                    (_slots_22_io_uop_prs2),
    .io_uop_prs3                    (_slots_22_io_uop_prs3),
    .io_uop_ppred                   (_slots_22_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_22_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_22_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_22_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_22_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_22_io_uop_stale_pdst),
    .io_uop_exception               (_slots_22_io_uop_exception),
    .io_uop_exc_cause               (_slots_22_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_22_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_22_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_22_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_22_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_22_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_22_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_22_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_22_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_22_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_22_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_22_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_22_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_22_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_22_io_uop_ldst),
    .io_uop_lrs1                    (_slots_22_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_22_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_22_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_22_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_22_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_22_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_22_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_22_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_22_io_uop_fp_val),
    .io_uop_fp_single               (_slots_22_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_22_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_22_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_22_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_22_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_22_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_22_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_22_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_23 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_23_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_22),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_23_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_55
         ? _slots_26_io_out_uop_uopc
         : _GEN_54 ? _slots_25_io_out_uop_uopc : _slots_24_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_55
         ? _slots_26_io_out_uop_inst
         : _GEN_54 ? _slots_25_io_out_uop_inst : _slots_24_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_55
         ? _slots_26_io_out_uop_debug_inst
         : _GEN_54 ? _slots_25_io_out_uop_debug_inst : _slots_24_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_55
         ? _slots_26_io_out_uop_is_rvc
         : _GEN_54 ? _slots_25_io_out_uop_is_rvc : _slots_24_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_55
         ? _slots_26_io_out_uop_debug_pc
         : _GEN_54 ? _slots_25_io_out_uop_debug_pc : _slots_24_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_55
         ? _slots_26_io_out_uop_iq_type
         : _GEN_54 ? _slots_25_io_out_uop_iq_type : _slots_24_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_55
         ? _slots_26_io_out_uop_fu_code
         : _GEN_54 ? _slots_25_io_out_uop_fu_code : _slots_24_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_55
         ? _slots_26_io_out_uop_iw_state
         : _GEN_54 ? _slots_25_io_out_uop_iw_state : _slots_24_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_55
         ? _slots_26_io_out_uop_iw_p1_poisoned
         : _GEN_54
             ? _slots_25_io_out_uop_iw_p1_poisoned
             : _slots_24_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_55
         ? _slots_26_io_out_uop_iw_p2_poisoned
         : _GEN_54
             ? _slots_25_io_out_uop_iw_p2_poisoned
             : _slots_24_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_55
         ? _slots_26_io_out_uop_is_br
         : _GEN_54 ? _slots_25_io_out_uop_is_br : _slots_24_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_55
         ? _slots_26_io_out_uop_is_jalr
         : _GEN_54 ? _slots_25_io_out_uop_is_jalr : _slots_24_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_55
         ? _slots_26_io_out_uop_is_jal
         : _GEN_54 ? _slots_25_io_out_uop_is_jal : _slots_24_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_55
         ? _slots_26_io_out_uop_is_sfb
         : _GEN_54 ? _slots_25_io_out_uop_is_sfb : _slots_24_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_55
         ? _slots_26_io_out_uop_br_mask
         : _GEN_54 ? _slots_25_io_out_uop_br_mask : _slots_24_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_55
         ? _slots_26_io_out_uop_br_tag
         : _GEN_54 ? _slots_25_io_out_uop_br_tag : _slots_24_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_55
         ? _slots_26_io_out_uop_ftq_idx
         : _GEN_54 ? _slots_25_io_out_uop_ftq_idx : _slots_24_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_55
         ? _slots_26_io_out_uop_edge_inst
         : _GEN_54 ? _slots_25_io_out_uop_edge_inst : _slots_24_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_55
         ? _slots_26_io_out_uop_pc_lob
         : _GEN_54 ? _slots_25_io_out_uop_pc_lob : _slots_24_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_55
         ? _slots_26_io_out_uop_taken
         : _GEN_54 ? _slots_25_io_out_uop_taken : _slots_24_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_55
         ? _slots_26_io_out_uop_imm_packed
         : _GEN_54 ? _slots_25_io_out_uop_imm_packed : _slots_24_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_55
         ? _slots_26_io_out_uop_csr_addr
         : _GEN_54 ? _slots_25_io_out_uop_csr_addr : _slots_24_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_55
         ? _slots_26_io_out_uop_rob_idx
         : _GEN_54 ? _slots_25_io_out_uop_rob_idx : _slots_24_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_55
         ? _slots_26_io_out_uop_ldq_idx
         : _GEN_54 ? _slots_25_io_out_uop_ldq_idx : _slots_24_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_55
         ? _slots_26_io_out_uop_stq_idx
         : _GEN_54 ? _slots_25_io_out_uop_stq_idx : _slots_24_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_55
         ? _slots_26_io_out_uop_rxq_idx
         : _GEN_54 ? _slots_25_io_out_uop_rxq_idx : _slots_24_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_55
         ? _slots_26_io_out_uop_pdst
         : _GEN_54 ? _slots_25_io_out_uop_pdst : _slots_24_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_55
         ? _slots_26_io_out_uop_prs1
         : _GEN_54 ? _slots_25_io_out_uop_prs1 : _slots_24_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_55
         ? _slots_26_io_out_uop_prs2
         : _GEN_54 ? _slots_25_io_out_uop_prs2 : _slots_24_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_55
         ? _slots_26_io_out_uop_prs3
         : _GEN_54 ? _slots_25_io_out_uop_prs3 : _slots_24_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_55
         ? _slots_26_io_out_uop_ppred
         : _GEN_54 ? _slots_25_io_out_uop_ppred : _slots_24_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_55
         ? _slots_26_io_out_uop_prs1_busy
         : _GEN_54 ? _slots_25_io_out_uop_prs1_busy : _slots_24_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_55
         ? _slots_26_io_out_uop_prs2_busy
         : _GEN_54 ? _slots_25_io_out_uop_prs2_busy : _slots_24_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_55
         ? _slots_26_io_out_uop_prs3_busy
         : _GEN_54 ? _slots_25_io_out_uop_prs3_busy : _slots_24_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_55
         ? _slots_26_io_out_uop_ppred_busy
         : _GEN_54 ? _slots_25_io_out_uop_ppred_busy : _slots_24_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_55
         ? _slots_26_io_out_uop_stale_pdst
         : _GEN_54 ? _slots_25_io_out_uop_stale_pdst : _slots_24_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_55
         ? _slots_26_io_out_uop_exception
         : _GEN_54 ? _slots_25_io_out_uop_exception : _slots_24_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_55
         ? _slots_26_io_out_uop_exc_cause
         : _GEN_54 ? _slots_25_io_out_uop_exc_cause : _slots_24_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_55
         ? _slots_26_io_out_uop_bypassable
         : _GEN_54 ? _slots_25_io_out_uop_bypassable : _slots_24_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_55
         ? _slots_26_io_out_uop_mem_cmd
         : _GEN_54 ? _slots_25_io_out_uop_mem_cmd : _slots_24_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_55
         ? _slots_26_io_out_uop_mem_size
         : _GEN_54 ? _slots_25_io_out_uop_mem_size : _slots_24_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_55
         ? _slots_26_io_out_uop_mem_signed
         : _GEN_54 ? _slots_25_io_out_uop_mem_signed : _slots_24_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_55
         ? _slots_26_io_out_uop_is_fence
         : _GEN_54 ? _slots_25_io_out_uop_is_fence : _slots_24_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_55
         ? _slots_26_io_out_uop_is_fencei
         : _GEN_54 ? _slots_25_io_out_uop_is_fencei : _slots_24_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_55
         ? _slots_26_io_out_uop_is_amo
         : _GEN_54 ? _slots_25_io_out_uop_is_amo : _slots_24_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_55
         ? _slots_26_io_out_uop_uses_ldq
         : _GEN_54 ? _slots_25_io_out_uop_uses_ldq : _slots_24_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_55
         ? _slots_26_io_out_uop_uses_stq
         : _GEN_54 ? _slots_25_io_out_uop_uses_stq : _slots_24_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_55
         ? _slots_26_io_out_uop_is_sys_pc2epc
         : _GEN_54
             ? _slots_25_io_out_uop_is_sys_pc2epc
             : _slots_24_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_55
         ? _slots_26_io_out_uop_is_unique
         : _GEN_54 ? _slots_25_io_out_uop_is_unique : _slots_24_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_55
         ? _slots_26_io_out_uop_flush_on_commit
         : _GEN_54
             ? _slots_25_io_out_uop_flush_on_commit
             : _slots_24_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_55
         ? _slots_26_io_out_uop_ldst_is_rs1
         : _GEN_54 ? _slots_25_io_out_uop_ldst_is_rs1 : _slots_24_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_55
         ? _slots_26_io_out_uop_ldst
         : _GEN_54 ? _slots_25_io_out_uop_ldst : _slots_24_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_55
         ? _slots_26_io_out_uop_lrs1
         : _GEN_54 ? _slots_25_io_out_uop_lrs1 : _slots_24_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_55
         ? _slots_26_io_out_uop_lrs2
         : _GEN_54 ? _slots_25_io_out_uop_lrs2 : _slots_24_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_55
         ? _slots_26_io_out_uop_lrs3
         : _GEN_54 ? _slots_25_io_out_uop_lrs3 : _slots_24_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_55
         ? _slots_26_io_out_uop_ldst_val
         : _GEN_54 ? _slots_25_io_out_uop_ldst_val : _slots_24_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_55
         ? _slots_26_io_out_uop_dst_rtype
         : _GEN_54 ? _slots_25_io_out_uop_dst_rtype : _slots_24_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_55
         ? _slots_26_io_out_uop_lrs1_rtype
         : _GEN_54 ? _slots_25_io_out_uop_lrs1_rtype : _slots_24_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_55
         ? _slots_26_io_out_uop_lrs2_rtype
         : _GEN_54 ? _slots_25_io_out_uop_lrs2_rtype : _slots_24_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_55
         ? _slots_26_io_out_uop_frs3_en
         : _GEN_54 ? _slots_25_io_out_uop_frs3_en : _slots_24_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_55
         ? _slots_26_io_out_uop_fp_val
         : _GEN_54 ? _slots_25_io_out_uop_fp_val : _slots_24_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_55
         ? _slots_26_io_out_uop_fp_single
         : _GEN_54 ? _slots_25_io_out_uop_fp_single : _slots_24_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_55
         ? _slots_26_io_out_uop_xcpt_pf_if
         : _GEN_54 ? _slots_25_io_out_uop_xcpt_pf_if : _slots_24_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_55
         ? _slots_26_io_out_uop_xcpt_ae_if
         : _GEN_54 ? _slots_25_io_out_uop_xcpt_ae_if : _slots_24_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_55
         ? _slots_26_io_out_uop_xcpt_ma_if
         : _GEN_54 ? _slots_25_io_out_uop_xcpt_ma_if : _slots_24_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_55
         ? _slots_26_io_out_uop_bp_debug_if
         : _GEN_54 ? _slots_25_io_out_uop_bp_debug_if : _slots_24_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_55
         ? _slots_26_io_out_uop_bp_xcpt_if
         : _GEN_54 ? _slots_25_io_out_uop_bp_xcpt_if : _slots_24_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_55
         ? _slots_26_io_out_uop_debug_fsrc
         : _GEN_54 ? _slots_25_io_out_uop_debug_fsrc : _slots_24_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_55
         ? _slots_26_io_out_uop_debug_tsrc
         : _GEN_54 ? _slots_25_io_out_uop_debug_tsrc : _slots_24_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_23_io_valid),
    .io_will_be_valid               (_slots_23_io_will_be_valid),
    .io_request                     (_slots_23_io_request),
    .io_out_uop_uopc                (_slots_23_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_23_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_23_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_23_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_23_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_23_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_23_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_23_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_23_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_23_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_23_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_23_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_23_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_23_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_23_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_23_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_23_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_23_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_23_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_23_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_23_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_23_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_23_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_23_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_23_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_23_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_23_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_23_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_23_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_23_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_23_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_23_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_23_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_23_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_23_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_23_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_23_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_23_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_23_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_23_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_23_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_23_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_23_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_23_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_23_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_23_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_23_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_23_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_23_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_23_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_23_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_23_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_23_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_23_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_23_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_23_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_23_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_23_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_23_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_23_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_23_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_23_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_23_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_23_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_23_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_23_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_23_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_23_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_23_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_23_io_uop_uopc),
    .io_uop_inst                    (_slots_23_io_uop_inst),
    .io_uop_debug_inst              (_slots_23_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_23_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_23_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_23_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_23_io_uop_fu_code),
    .io_uop_iw_state                (_slots_23_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_23_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_23_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_23_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_23_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_23_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_23_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_23_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_23_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_23_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_23_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_23_io_uop_pc_lob),
    .io_uop_taken                   (_slots_23_io_uop_taken),
    .io_uop_imm_packed              (_slots_23_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_23_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_23_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_23_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_23_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_23_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_23_io_uop_pdst),
    .io_uop_prs1                    (_slots_23_io_uop_prs1),
    .io_uop_prs2                    (_slots_23_io_uop_prs2),
    .io_uop_prs3                    (_slots_23_io_uop_prs3),
    .io_uop_ppred                   (_slots_23_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_23_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_23_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_23_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_23_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_23_io_uop_stale_pdst),
    .io_uop_exception               (_slots_23_io_uop_exception),
    .io_uop_exc_cause               (_slots_23_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_23_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_23_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_23_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_23_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_23_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_23_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_23_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_23_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_23_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_23_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_23_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_23_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_23_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_23_io_uop_ldst),
    .io_uop_lrs1                    (_slots_23_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_23_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_23_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_23_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_23_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_23_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_23_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_23_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_23_io_uop_fp_val),
    .io_uop_fp_single               (_slots_23_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_23_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_23_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_23_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_23_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_23_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_23_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_23_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_24 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_24_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_23),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_24_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_57
         ? _slots_27_io_out_uop_uopc
         : _GEN_56 ? _slots_26_io_out_uop_uopc : _slots_25_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_57
         ? _slots_27_io_out_uop_inst
         : _GEN_56 ? _slots_26_io_out_uop_inst : _slots_25_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_57
         ? _slots_27_io_out_uop_debug_inst
         : _GEN_56 ? _slots_26_io_out_uop_debug_inst : _slots_25_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_57
         ? _slots_27_io_out_uop_is_rvc
         : _GEN_56 ? _slots_26_io_out_uop_is_rvc : _slots_25_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_57
         ? _slots_27_io_out_uop_debug_pc
         : _GEN_56 ? _slots_26_io_out_uop_debug_pc : _slots_25_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_57
         ? _slots_27_io_out_uop_iq_type
         : _GEN_56 ? _slots_26_io_out_uop_iq_type : _slots_25_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_57
         ? _slots_27_io_out_uop_fu_code
         : _GEN_56 ? _slots_26_io_out_uop_fu_code : _slots_25_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_57
         ? _slots_27_io_out_uop_iw_state
         : _GEN_56 ? _slots_26_io_out_uop_iw_state : _slots_25_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_57
         ? _slots_27_io_out_uop_iw_p1_poisoned
         : _GEN_56
             ? _slots_26_io_out_uop_iw_p1_poisoned
             : _slots_25_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_57
         ? _slots_27_io_out_uop_iw_p2_poisoned
         : _GEN_56
             ? _slots_26_io_out_uop_iw_p2_poisoned
             : _slots_25_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_57
         ? _slots_27_io_out_uop_is_br
         : _GEN_56 ? _slots_26_io_out_uop_is_br : _slots_25_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_57
         ? _slots_27_io_out_uop_is_jalr
         : _GEN_56 ? _slots_26_io_out_uop_is_jalr : _slots_25_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_57
         ? _slots_27_io_out_uop_is_jal
         : _GEN_56 ? _slots_26_io_out_uop_is_jal : _slots_25_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_57
         ? _slots_27_io_out_uop_is_sfb
         : _GEN_56 ? _slots_26_io_out_uop_is_sfb : _slots_25_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_57
         ? _slots_27_io_out_uop_br_mask
         : _GEN_56 ? _slots_26_io_out_uop_br_mask : _slots_25_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_57
         ? _slots_27_io_out_uop_br_tag
         : _GEN_56 ? _slots_26_io_out_uop_br_tag : _slots_25_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_57
         ? _slots_27_io_out_uop_ftq_idx
         : _GEN_56 ? _slots_26_io_out_uop_ftq_idx : _slots_25_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_57
         ? _slots_27_io_out_uop_edge_inst
         : _GEN_56 ? _slots_26_io_out_uop_edge_inst : _slots_25_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_57
         ? _slots_27_io_out_uop_pc_lob
         : _GEN_56 ? _slots_26_io_out_uop_pc_lob : _slots_25_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_57
         ? _slots_27_io_out_uop_taken
         : _GEN_56 ? _slots_26_io_out_uop_taken : _slots_25_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_57
         ? _slots_27_io_out_uop_imm_packed
         : _GEN_56 ? _slots_26_io_out_uop_imm_packed : _slots_25_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_57
         ? _slots_27_io_out_uop_csr_addr
         : _GEN_56 ? _slots_26_io_out_uop_csr_addr : _slots_25_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_57
         ? _slots_27_io_out_uop_rob_idx
         : _GEN_56 ? _slots_26_io_out_uop_rob_idx : _slots_25_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_57
         ? _slots_27_io_out_uop_ldq_idx
         : _GEN_56 ? _slots_26_io_out_uop_ldq_idx : _slots_25_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_57
         ? _slots_27_io_out_uop_stq_idx
         : _GEN_56 ? _slots_26_io_out_uop_stq_idx : _slots_25_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_57
         ? _slots_27_io_out_uop_rxq_idx
         : _GEN_56 ? _slots_26_io_out_uop_rxq_idx : _slots_25_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_57
         ? _slots_27_io_out_uop_pdst
         : _GEN_56 ? _slots_26_io_out_uop_pdst : _slots_25_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_57
         ? _slots_27_io_out_uop_prs1
         : _GEN_56 ? _slots_26_io_out_uop_prs1 : _slots_25_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_57
         ? _slots_27_io_out_uop_prs2
         : _GEN_56 ? _slots_26_io_out_uop_prs2 : _slots_25_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_57
         ? _slots_27_io_out_uop_prs3
         : _GEN_56 ? _slots_26_io_out_uop_prs3 : _slots_25_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_57
         ? _slots_27_io_out_uop_ppred
         : _GEN_56 ? _slots_26_io_out_uop_ppred : _slots_25_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_57
         ? _slots_27_io_out_uop_prs1_busy
         : _GEN_56 ? _slots_26_io_out_uop_prs1_busy : _slots_25_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_57
         ? _slots_27_io_out_uop_prs2_busy
         : _GEN_56 ? _slots_26_io_out_uop_prs2_busy : _slots_25_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_57
         ? _slots_27_io_out_uop_prs3_busy
         : _GEN_56 ? _slots_26_io_out_uop_prs3_busy : _slots_25_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_57
         ? _slots_27_io_out_uop_ppred_busy
         : _GEN_56 ? _slots_26_io_out_uop_ppred_busy : _slots_25_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_57
         ? _slots_27_io_out_uop_stale_pdst
         : _GEN_56 ? _slots_26_io_out_uop_stale_pdst : _slots_25_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_57
         ? _slots_27_io_out_uop_exception
         : _GEN_56 ? _slots_26_io_out_uop_exception : _slots_25_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_57
         ? _slots_27_io_out_uop_exc_cause
         : _GEN_56 ? _slots_26_io_out_uop_exc_cause : _slots_25_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_57
         ? _slots_27_io_out_uop_bypassable
         : _GEN_56 ? _slots_26_io_out_uop_bypassable : _slots_25_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_57
         ? _slots_27_io_out_uop_mem_cmd
         : _GEN_56 ? _slots_26_io_out_uop_mem_cmd : _slots_25_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_57
         ? _slots_27_io_out_uop_mem_size
         : _GEN_56 ? _slots_26_io_out_uop_mem_size : _slots_25_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_57
         ? _slots_27_io_out_uop_mem_signed
         : _GEN_56 ? _slots_26_io_out_uop_mem_signed : _slots_25_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_57
         ? _slots_27_io_out_uop_is_fence
         : _GEN_56 ? _slots_26_io_out_uop_is_fence : _slots_25_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_57
         ? _slots_27_io_out_uop_is_fencei
         : _GEN_56 ? _slots_26_io_out_uop_is_fencei : _slots_25_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_57
         ? _slots_27_io_out_uop_is_amo
         : _GEN_56 ? _slots_26_io_out_uop_is_amo : _slots_25_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_57
         ? _slots_27_io_out_uop_uses_ldq
         : _GEN_56 ? _slots_26_io_out_uop_uses_ldq : _slots_25_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_57
         ? _slots_27_io_out_uop_uses_stq
         : _GEN_56 ? _slots_26_io_out_uop_uses_stq : _slots_25_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_57
         ? _slots_27_io_out_uop_is_sys_pc2epc
         : _GEN_56
             ? _slots_26_io_out_uop_is_sys_pc2epc
             : _slots_25_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_57
         ? _slots_27_io_out_uop_is_unique
         : _GEN_56 ? _slots_26_io_out_uop_is_unique : _slots_25_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_57
         ? _slots_27_io_out_uop_flush_on_commit
         : _GEN_56
             ? _slots_26_io_out_uop_flush_on_commit
             : _slots_25_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_57
         ? _slots_27_io_out_uop_ldst_is_rs1
         : _GEN_56 ? _slots_26_io_out_uop_ldst_is_rs1 : _slots_25_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_57
         ? _slots_27_io_out_uop_ldst
         : _GEN_56 ? _slots_26_io_out_uop_ldst : _slots_25_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_57
         ? _slots_27_io_out_uop_lrs1
         : _GEN_56 ? _slots_26_io_out_uop_lrs1 : _slots_25_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_57
         ? _slots_27_io_out_uop_lrs2
         : _GEN_56 ? _slots_26_io_out_uop_lrs2 : _slots_25_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_57
         ? _slots_27_io_out_uop_lrs3
         : _GEN_56 ? _slots_26_io_out_uop_lrs3 : _slots_25_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_57
         ? _slots_27_io_out_uop_ldst_val
         : _GEN_56 ? _slots_26_io_out_uop_ldst_val : _slots_25_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_57
         ? _slots_27_io_out_uop_dst_rtype
         : _GEN_56 ? _slots_26_io_out_uop_dst_rtype : _slots_25_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_57
         ? _slots_27_io_out_uop_lrs1_rtype
         : _GEN_56 ? _slots_26_io_out_uop_lrs1_rtype : _slots_25_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_57
         ? _slots_27_io_out_uop_lrs2_rtype
         : _GEN_56 ? _slots_26_io_out_uop_lrs2_rtype : _slots_25_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_57
         ? _slots_27_io_out_uop_frs3_en
         : _GEN_56 ? _slots_26_io_out_uop_frs3_en : _slots_25_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_57
         ? _slots_27_io_out_uop_fp_val
         : _GEN_56 ? _slots_26_io_out_uop_fp_val : _slots_25_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_57
         ? _slots_27_io_out_uop_fp_single
         : _GEN_56 ? _slots_26_io_out_uop_fp_single : _slots_25_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_57
         ? _slots_27_io_out_uop_xcpt_pf_if
         : _GEN_56 ? _slots_26_io_out_uop_xcpt_pf_if : _slots_25_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_57
         ? _slots_27_io_out_uop_xcpt_ae_if
         : _GEN_56 ? _slots_26_io_out_uop_xcpt_ae_if : _slots_25_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_57
         ? _slots_27_io_out_uop_xcpt_ma_if
         : _GEN_56 ? _slots_26_io_out_uop_xcpt_ma_if : _slots_25_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_57
         ? _slots_27_io_out_uop_bp_debug_if
         : _GEN_56 ? _slots_26_io_out_uop_bp_debug_if : _slots_25_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_57
         ? _slots_27_io_out_uop_bp_xcpt_if
         : _GEN_56 ? _slots_26_io_out_uop_bp_xcpt_if : _slots_25_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_57
         ? _slots_27_io_out_uop_debug_fsrc
         : _GEN_56 ? _slots_26_io_out_uop_debug_fsrc : _slots_25_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_57
         ? _slots_27_io_out_uop_debug_tsrc
         : _GEN_56 ? _slots_26_io_out_uop_debug_tsrc : _slots_25_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_24_io_valid),
    .io_will_be_valid               (_slots_24_io_will_be_valid),
    .io_request                     (_slots_24_io_request),
    .io_out_uop_uopc                (_slots_24_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_24_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_24_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_24_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_24_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_24_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_24_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_24_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_24_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_24_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_24_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_24_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_24_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_24_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_24_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_24_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_24_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_24_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_24_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_24_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_24_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_24_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_24_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_24_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_24_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_24_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_24_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_24_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_24_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_24_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_24_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_24_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_24_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_24_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_24_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_24_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_24_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_24_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_24_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_24_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_24_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_24_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_24_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_24_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_24_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_24_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_24_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_24_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_24_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_24_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_24_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_24_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_24_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_24_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_24_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_24_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_24_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_24_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_24_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_24_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_24_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_24_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_24_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_24_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_24_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_24_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_24_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_24_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_24_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_24_io_uop_uopc),
    .io_uop_inst                    (_slots_24_io_uop_inst),
    .io_uop_debug_inst              (_slots_24_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_24_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_24_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_24_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_24_io_uop_fu_code),
    .io_uop_iw_state                (_slots_24_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_24_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_24_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_24_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_24_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_24_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_24_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_24_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_24_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_24_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_24_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_24_io_uop_pc_lob),
    .io_uop_taken                   (_slots_24_io_uop_taken),
    .io_uop_imm_packed              (_slots_24_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_24_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_24_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_24_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_24_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_24_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_24_io_uop_pdst),
    .io_uop_prs1                    (_slots_24_io_uop_prs1),
    .io_uop_prs2                    (_slots_24_io_uop_prs2),
    .io_uop_prs3                    (_slots_24_io_uop_prs3),
    .io_uop_ppred                   (_slots_24_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_24_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_24_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_24_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_24_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_24_io_uop_stale_pdst),
    .io_uop_exception               (_slots_24_io_uop_exception),
    .io_uop_exc_cause               (_slots_24_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_24_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_24_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_24_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_24_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_24_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_24_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_24_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_24_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_24_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_24_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_24_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_24_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_24_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_24_io_uop_ldst),
    .io_uop_lrs1                    (_slots_24_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_24_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_24_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_24_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_24_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_24_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_24_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_24_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_24_io_uop_fp_val),
    .io_uop_fp_single               (_slots_24_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_24_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_24_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_24_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_24_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_24_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_24_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_24_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_25 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_25_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_24),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_25_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_59
         ? _slots_28_io_out_uop_uopc
         : _GEN_58 ? _slots_27_io_out_uop_uopc : _slots_26_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_59
         ? _slots_28_io_out_uop_inst
         : _GEN_58 ? _slots_27_io_out_uop_inst : _slots_26_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_59
         ? _slots_28_io_out_uop_debug_inst
         : _GEN_58 ? _slots_27_io_out_uop_debug_inst : _slots_26_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_59
         ? _slots_28_io_out_uop_is_rvc
         : _GEN_58 ? _slots_27_io_out_uop_is_rvc : _slots_26_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_59
         ? _slots_28_io_out_uop_debug_pc
         : _GEN_58 ? _slots_27_io_out_uop_debug_pc : _slots_26_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_59
         ? _slots_28_io_out_uop_iq_type
         : _GEN_58 ? _slots_27_io_out_uop_iq_type : _slots_26_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_59
         ? _slots_28_io_out_uop_fu_code
         : _GEN_58 ? _slots_27_io_out_uop_fu_code : _slots_26_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_59
         ? _slots_28_io_out_uop_iw_state
         : _GEN_58 ? _slots_27_io_out_uop_iw_state : _slots_26_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_59
         ? _slots_28_io_out_uop_iw_p1_poisoned
         : _GEN_58
             ? _slots_27_io_out_uop_iw_p1_poisoned
             : _slots_26_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_59
         ? _slots_28_io_out_uop_iw_p2_poisoned
         : _GEN_58
             ? _slots_27_io_out_uop_iw_p2_poisoned
             : _slots_26_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_59
         ? _slots_28_io_out_uop_is_br
         : _GEN_58 ? _slots_27_io_out_uop_is_br : _slots_26_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_59
         ? _slots_28_io_out_uop_is_jalr
         : _GEN_58 ? _slots_27_io_out_uop_is_jalr : _slots_26_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_59
         ? _slots_28_io_out_uop_is_jal
         : _GEN_58 ? _slots_27_io_out_uop_is_jal : _slots_26_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_59
         ? _slots_28_io_out_uop_is_sfb
         : _GEN_58 ? _slots_27_io_out_uop_is_sfb : _slots_26_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_59
         ? _slots_28_io_out_uop_br_mask
         : _GEN_58 ? _slots_27_io_out_uop_br_mask : _slots_26_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_59
         ? _slots_28_io_out_uop_br_tag
         : _GEN_58 ? _slots_27_io_out_uop_br_tag : _slots_26_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_59
         ? _slots_28_io_out_uop_ftq_idx
         : _GEN_58 ? _slots_27_io_out_uop_ftq_idx : _slots_26_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_59
         ? _slots_28_io_out_uop_edge_inst
         : _GEN_58 ? _slots_27_io_out_uop_edge_inst : _slots_26_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_59
         ? _slots_28_io_out_uop_pc_lob
         : _GEN_58 ? _slots_27_io_out_uop_pc_lob : _slots_26_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_59
         ? _slots_28_io_out_uop_taken
         : _GEN_58 ? _slots_27_io_out_uop_taken : _slots_26_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_59
         ? _slots_28_io_out_uop_imm_packed
         : _GEN_58 ? _slots_27_io_out_uop_imm_packed : _slots_26_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_59
         ? _slots_28_io_out_uop_csr_addr
         : _GEN_58 ? _slots_27_io_out_uop_csr_addr : _slots_26_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_59
         ? _slots_28_io_out_uop_rob_idx
         : _GEN_58 ? _slots_27_io_out_uop_rob_idx : _slots_26_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_59
         ? _slots_28_io_out_uop_ldq_idx
         : _GEN_58 ? _slots_27_io_out_uop_ldq_idx : _slots_26_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_59
         ? _slots_28_io_out_uop_stq_idx
         : _GEN_58 ? _slots_27_io_out_uop_stq_idx : _slots_26_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_59
         ? _slots_28_io_out_uop_rxq_idx
         : _GEN_58 ? _slots_27_io_out_uop_rxq_idx : _slots_26_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_59
         ? _slots_28_io_out_uop_pdst
         : _GEN_58 ? _slots_27_io_out_uop_pdst : _slots_26_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_59
         ? _slots_28_io_out_uop_prs1
         : _GEN_58 ? _slots_27_io_out_uop_prs1 : _slots_26_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_59
         ? _slots_28_io_out_uop_prs2
         : _GEN_58 ? _slots_27_io_out_uop_prs2 : _slots_26_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_59
         ? _slots_28_io_out_uop_prs3
         : _GEN_58 ? _slots_27_io_out_uop_prs3 : _slots_26_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_59
         ? _slots_28_io_out_uop_ppred
         : _GEN_58 ? _slots_27_io_out_uop_ppred : _slots_26_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_59
         ? _slots_28_io_out_uop_prs1_busy
         : _GEN_58 ? _slots_27_io_out_uop_prs1_busy : _slots_26_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_59
         ? _slots_28_io_out_uop_prs2_busy
         : _GEN_58 ? _slots_27_io_out_uop_prs2_busy : _slots_26_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_59
         ? _slots_28_io_out_uop_prs3_busy
         : _GEN_58 ? _slots_27_io_out_uop_prs3_busy : _slots_26_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_59
         ? _slots_28_io_out_uop_ppred_busy
         : _GEN_58 ? _slots_27_io_out_uop_ppred_busy : _slots_26_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_59
         ? _slots_28_io_out_uop_stale_pdst
         : _GEN_58 ? _slots_27_io_out_uop_stale_pdst : _slots_26_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_59
         ? _slots_28_io_out_uop_exception
         : _GEN_58 ? _slots_27_io_out_uop_exception : _slots_26_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_59
         ? _slots_28_io_out_uop_exc_cause
         : _GEN_58 ? _slots_27_io_out_uop_exc_cause : _slots_26_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_59
         ? _slots_28_io_out_uop_bypassable
         : _GEN_58 ? _slots_27_io_out_uop_bypassable : _slots_26_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_59
         ? _slots_28_io_out_uop_mem_cmd
         : _GEN_58 ? _slots_27_io_out_uop_mem_cmd : _slots_26_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_59
         ? _slots_28_io_out_uop_mem_size
         : _GEN_58 ? _slots_27_io_out_uop_mem_size : _slots_26_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_59
         ? _slots_28_io_out_uop_mem_signed
         : _GEN_58 ? _slots_27_io_out_uop_mem_signed : _slots_26_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_59
         ? _slots_28_io_out_uop_is_fence
         : _GEN_58 ? _slots_27_io_out_uop_is_fence : _slots_26_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_59
         ? _slots_28_io_out_uop_is_fencei
         : _GEN_58 ? _slots_27_io_out_uop_is_fencei : _slots_26_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_59
         ? _slots_28_io_out_uop_is_amo
         : _GEN_58 ? _slots_27_io_out_uop_is_amo : _slots_26_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_59
         ? _slots_28_io_out_uop_uses_ldq
         : _GEN_58 ? _slots_27_io_out_uop_uses_ldq : _slots_26_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_59
         ? _slots_28_io_out_uop_uses_stq
         : _GEN_58 ? _slots_27_io_out_uop_uses_stq : _slots_26_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_59
         ? _slots_28_io_out_uop_is_sys_pc2epc
         : _GEN_58
             ? _slots_27_io_out_uop_is_sys_pc2epc
             : _slots_26_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_59
         ? _slots_28_io_out_uop_is_unique
         : _GEN_58 ? _slots_27_io_out_uop_is_unique : _slots_26_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_59
         ? _slots_28_io_out_uop_flush_on_commit
         : _GEN_58
             ? _slots_27_io_out_uop_flush_on_commit
             : _slots_26_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_59
         ? _slots_28_io_out_uop_ldst_is_rs1
         : _GEN_58 ? _slots_27_io_out_uop_ldst_is_rs1 : _slots_26_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_59
         ? _slots_28_io_out_uop_ldst
         : _GEN_58 ? _slots_27_io_out_uop_ldst : _slots_26_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_59
         ? _slots_28_io_out_uop_lrs1
         : _GEN_58 ? _slots_27_io_out_uop_lrs1 : _slots_26_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_59
         ? _slots_28_io_out_uop_lrs2
         : _GEN_58 ? _slots_27_io_out_uop_lrs2 : _slots_26_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_59
         ? _slots_28_io_out_uop_lrs3
         : _GEN_58 ? _slots_27_io_out_uop_lrs3 : _slots_26_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_59
         ? _slots_28_io_out_uop_ldst_val
         : _GEN_58 ? _slots_27_io_out_uop_ldst_val : _slots_26_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_59
         ? _slots_28_io_out_uop_dst_rtype
         : _GEN_58 ? _slots_27_io_out_uop_dst_rtype : _slots_26_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_59
         ? _slots_28_io_out_uop_lrs1_rtype
         : _GEN_58 ? _slots_27_io_out_uop_lrs1_rtype : _slots_26_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_59
         ? _slots_28_io_out_uop_lrs2_rtype
         : _GEN_58 ? _slots_27_io_out_uop_lrs2_rtype : _slots_26_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_59
         ? _slots_28_io_out_uop_frs3_en
         : _GEN_58 ? _slots_27_io_out_uop_frs3_en : _slots_26_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_59
         ? _slots_28_io_out_uop_fp_val
         : _GEN_58 ? _slots_27_io_out_uop_fp_val : _slots_26_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_59
         ? _slots_28_io_out_uop_fp_single
         : _GEN_58 ? _slots_27_io_out_uop_fp_single : _slots_26_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_59
         ? _slots_28_io_out_uop_xcpt_pf_if
         : _GEN_58 ? _slots_27_io_out_uop_xcpt_pf_if : _slots_26_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_59
         ? _slots_28_io_out_uop_xcpt_ae_if
         : _GEN_58 ? _slots_27_io_out_uop_xcpt_ae_if : _slots_26_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_59
         ? _slots_28_io_out_uop_xcpt_ma_if
         : _GEN_58 ? _slots_27_io_out_uop_xcpt_ma_if : _slots_26_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_59
         ? _slots_28_io_out_uop_bp_debug_if
         : _GEN_58 ? _slots_27_io_out_uop_bp_debug_if : _slots_26_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_59
         ? _slots_28_io_out_uop_bp_xcpt_if
         : _GEN_58 ? _slots_27_io_out_uop_bp_xcpt_if : _slots_26_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_59
         ? _slots_28_io_out_uop_debug_fsrc
         : _GEN_58 ? _slots_27_io_out_uop_debug_fsrc : _slots_26_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_59
         ? _slots_28_io_out_uop_debug_tsrc
         : _GEN_58 ? _slots_27_io_out_uop_debug_tsrc : _slots_26_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_25_io_valid),
    .io_will_be_valid               (_slots_25_io_will_be_valid),
    .io_request                     (_slots_25_io_request),
    .io_out_uop_uopc                (_slots_25_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_25_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_25_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_25_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_25_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_25_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_25_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_25_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_25_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_25_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_25_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_25_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_25_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_25_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_25_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_25_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_25_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_25_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_25_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_25_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_25_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_25_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_25_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_25_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_25_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_25_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_25_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_25_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_25_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_25_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_25_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_25_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_25_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_25_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_25_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_25_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_25_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_25_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_25_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_25_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_25_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_25_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_25_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_25_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_25_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_25_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_25_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_25_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_25_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_25_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_25_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_25_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_25_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_25_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_25_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_25_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_25_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_25_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_25_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_25_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_25_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_25_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_25_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_25_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_25_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_25_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_25_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_25_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_25_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_25_io_uop_uopc),
    .io_uop_inst                    (_slots_25_io_uop_inst),
    .io_uop_debug_inst              (_slots_25_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_25_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_25_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_25_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_25_io_uop_fu_code),
    .io_uop_iw_state                (_slots_25_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_25_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_25_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_25_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_25_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_25_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_25_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_25_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_25_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_25_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_25_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_25_io_uop_pc_lob),
    .io_uop_taken                   (_slots_25_io_uop_taken),
    .io_uop_imm_packed              (_slots_25_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_25_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_25_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_25_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_25_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_25_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_25_io_uop_pdst),
    .io_uop_prs1                    (_slots_25_io_uop_prs1),
    .io_uop_prs2                    (_slots_25_io_uop_prs2),
    .io_uop_prs3                    (_slots_25_io_uop_prs3),
    .io_uop_ppred                   (_slots_25_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_25_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_25_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_25_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_25_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_25_io_uop_stale_pdst),
    .io_uop_exception               (_slots_25_io_uop_exception),
    .io_uop_exc_cause               (_slots_25_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_25_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_25_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_25_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_25_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_25_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_25_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_25_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_25_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_25_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_25_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_25_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_25_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_25_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_25_io_uop_ldst),
    .io_uop_lrs1                    (_slots_25_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_25_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_25_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_25_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_25_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_25_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_25_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_25_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_25_io_uop_fp_val),
    .io_uop_fp_single               (_slots_25_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_25_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_25_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_25_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_25_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_25_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_25_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_25_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_26 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_26_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_25),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_26_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_61
         ? _slots_29_io_out_uop_uopc
         : _GEN_60 ? _slots_28_io_out_uop_uopc : _slots_27_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_61
         ? _slots_29_io_out_uop_inst
         : _GEN_60 ? _slots_28_io_out_uop_inst : _slots_27_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_61
         ? _slots_29_io_out_uop_debug_inst
         : _GEN_60 ? _slots_28_io_out_uop_debug_inst : _slots_27_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_61
         ? _slots_29_io_out_uop_is_rvc
         : _GEN_60 ? _slots_28_io_out_uop_is_rvc : _slots_27_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_61
         ? _slots_29_io_out_uop_debug_pc
         : _GEN_60 ? _slots_28_io_out_uop_debug_pc : _slots_27_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_61
         ? _slots_29_io_out_uop_iq_type
         : _GEN_60 ? _slots_28_io_out_uop_iq_type : _slots_27_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_61
         ? _slots_29_io_out_uop_fu_code
         : _GEN_60 ? _slots_28_io_out_uop_fu_code : _slots_27_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_61
         ? _slots_29_io_out_uop_iw_state
         : _GEN_60 ? _slots_28_io_out_uop_iw_state : _slots_27_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_61
         ? _slots_29_io_out_uop_iw_p1_poisoned
         : _GEN_60
             ? _slots_28_io_out_uop_iw_p1_poisoned
             : _slots_27_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_61
         ? _slots_29_io_out_uop_iw_p2_poisoned
         : _GEN_60
             ? _slots_28_io_out_uop_iw_p2_poisoned
             : _slots_27_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_61
         ? _slots_29_io_out_uop_is_br
         : _GEN_60 ? _slots_28_io_out_uop_is_br : _slots_27_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_61
         ? _slots_29_io_out_uop_is_jalr
         : _GEN_60 ? _slots_28_io_out_uop_is_jalr : _slots_27_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_61
         ? _slots_29_io_out_uop_is_jal
         : _GEN_60 ? _slots_28_io_out_uop_is_jal : _slots_27_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_61
         ? _slots_29_io_out_uop_is_sfb
         : _GEN_60 ? _slots_28_io_out_uop_is_sfb : _slots_27_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_61
         ? _slots_29_io_out_uop_br_mask
         : _GEN_60 ? _slots_28_io_out_uop_br_mask : _slots_27_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_61
         ? _slots_29_io_out_uop_br_tag
         : _GEN_60 ? _slots_28_io_out_uop_br_tag : _slots_27_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_61
         ? _slots_29_io_out_uop_ftq_idx
         : _GEN_60 ? _slots_28_io_out_uop_ftq_idx : _slots_27_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_61
         ? _slots_29_io_out_uop_edge_inst
         : _GEN_60 ? _slots_28_io_out_uop_edge_inst : _slots_27_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_61
         ? _slots_29_io_out_uop_pc_lob
         : _GEN_60 ? _slots_28_io_out_uop_pc_lob : _slots_27_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_61
         ? _slots_29_io_out_uop_taken
         : _GEN_60 ? _slots_28_io_out_uop_taken : _slots_27_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_61
         ? _slots_29_io_out_uop_imm_packed
         : _GEN_60 ? _slots_28_io_out_uop_imm_packed : _slots_27_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_61
         ? _slots_29_io_out_uop_csr_addr
         : _GEN_60 ? _slots_28_io_out_uop_csr_addr : _slots_27_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_61
         ? _slots_29_io_out_uop_rob_idx
         : _GEN_60 ? _slots_28_io_out_uop_rob_idx : _slots_27_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_61
         ? _slots_29_io_out_uop_ldq_idx
         : _GEN_60 ? _slots_28_io_out_uop_ldq_idx : _slots_27_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_61
         ? _slots_29_io_out_uop_stq_idx
         : _GEN_60 ? _slots_28_io_out_uop_stq_idx : _slots_27_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_61
         ? _slots_29_io_out_uop_rxq_idx
         : _GEN_60 ? _slots_28_io_out_uop_rxq_idx : _slots_27_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_61
         ? _slots_29_io_out_uop_pdst
         : _GEN_60 ? _slots_28_io_out_uop_pdst : _slots_27_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_61
         ? _slots_29_io_out_uop_prs1
         : _GEN_60 ? _slots_28_io_out_uop_prs1 : _slots_27_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_61
         ? _slots_29_io_out_uop_prs2
         : _GEN_60 ? _slots_28_io_out_uop_prs2 : _slots_27_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_61
         ? _slots_29_io_out_uop_prs3
         : _GEN_60 ? _slots_28_io_out_uop_prs3 : _slots_27_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_61
         ? _slots_29_io_out_uop_ppred
         : _GEN_60 ? _slots_28_io_out_uop_ppred : _slots_27_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_61
         ? _slots_29_io_out_uop_prs1_busy
         : _GEN_60 ? _slots_28_io_out_uop_prs1_busy : _slots_27_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_61
         ? _slots_29_io_out_uop_prs2_busy
         : _GEN_60 ? _slots_28_io_out_uop_prs2_busy : _slots_27_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_61
         ? _slots_29_io_out_uop_prs3_busy
         : _GEN_60 ? _slots_28_io_out_uop_prs3_busy : _slots_27_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_61
         ? _slots_29_io_out_uop_ppred_busy
         : _GEN_60 ? _slots_28_io_out_uop_ppred_busy : _slots_27_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_61
         ? _slots_29_io_out_uop_stale_pdst
         : _GEN_60 ? _slots_28_io_out_uop_stale_pdst : _slots_27_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_61
         ? _slots_29_io_out_uop_exception
         : _GEN_60 ? _slots_28_io_out_uop_exception : _slots_27_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_61
         ? _slots_29_io_out_uop_exc_cause
         : _GEN_60 ? _slots_28_io_out_uop_exc_cause : _slots_27_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_61
         ? _slots_29_io_out_uop_bypassable
         : _GEN_60 ? _slots_28_io_out_uop_bypassable : _slots_27_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_61
         ? _slots_29_io_out_uop_mem_cmd
         : _GEN_60 ? _slots_28_io_out_uop_mem_cmd : _slots_27_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_61
         ? _slots_29_io_out_uop_mem_size
         : _GEN_60 ? _slots_28_io_out_uop_mem_size : _slots_27_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_61
         ? _slots_29_io_out_uop_mem_signed
         : _GEN_60 ? _slots_28_io_out_uop_mem_signed : _slots_27_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_61
         ? _slots_29_io_out_uop_is_fence
         : _GEN_60 ? _slots_28_io_out_uop_is_fence : _slots_27_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_61
         ? _slots_29_io_out_uop_is_fencei
         : _GEN_60 ? _slots_28_io_out_uop_is_fencei : _slots_27_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_61
         ? _slots_29_io_out_uop_is_amo
         : _GEN_60 ? _slots_28_io_out_uop_is_amo : _slots_27_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_61
         ? _slots_29_io_out_uop_uses_ldq
         : _GEN_60 ? _slots_28_io_out_uop_uses_ldq : _slots_27_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_61
         ? _slots_29_io_out_uop_uses_stq
         : _GEN_60 ? _slots_28_io_out_uop_uses_stq : _slots_27_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_61
         ? _slots_29_io_out_uop_is_sys_pc2epc
         : _GEN_60
             ? _slots_28_io_out_uop_is_sys_pc2epc
             : _slots_27_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_61
         ? _slots_29_io_out_uop_is_unique
         : _GEN_60 ? _slots_28_io_out_uop_is_unique : _slots_27_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_61
         ? _slots_29_io_out_uop_flush_on_commit
         : _GEN_60
             ? _slots_28_io_out_uop_flush_on_commit
             : _slots_27_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_61
         ? _slots_29_io_out_uop_ldst_is_rs1
         : _GEN_60 ? _slots_28_io_out_uop_ldst_is_rs1 : _slots_27_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_61
         ? _slots_29_io_out_uop_ldst
         : _GEN_60 ? _slots_28_io_out_uop_ldst : _slots_27_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_61
         ? _slots_29_io_out_uop_lrs1
         : _GEN_60 ? _slots_28_io_out_uop_lrs1 : _slots_27_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_61
         ? _slots_29_io_out_uop_lrs2
         : _GEN_60 ? _slots_28_io_out_uop_lrs2 : _slots_27_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_61
         ? _slots_29_io_out_uop_lrs3
         : _GEN_60 ? _slots_28_io_out_uop_lrs3 : _slots_27_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_61
         ? _slots_29_io_out_uop_ldst_val
         : _GEN_60 ? _slots_28_io_out_uop_ldst_val : _slots_27_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_61
         ? _slots_29_io_out_uop_dst_rtype
         : _GEN_60 ? _slots_28_io_out_uop_dst_rtype : _slots_27_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_61
         ? _slots_29_io_out_uop_lrs1_rtype
         : _GEN_60 ? _slots_28_io_out_uop_lrs1_rtype : _slots_27_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_61
         ? _slots_29_io_out_uop_lrs2_rtype
         : _GEN_60 ? _slots_28_io_out_uop_lrs2_rtype : _slots_27_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_61
         ? _slots_29_io_out_uop_frs3_en
         : _GEN_60 ? _slots_28_io_out_uop_frs3_en : _slots_27_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_61
         ? _slots_29_io_out_uop_fp_val
         : _GEN_60 ? _slots_28_io_out_uop_fp_val : _slots_27_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_61
         ? _slots_29_io_out_uop_fp_single
         : _GEN_60 ? _slots_28_io_out_uop_fp_single : _slots_27_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_61
         ? _slots_29_io_out_uop_xcpt_pf_if
         : _GEN_60 ? _slots_28_io_out_uop_xcpt_pf_if : _slots_27_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_61
         ? _slots_29_io_out_uop_xcpt_ae_if
         : _GEN_60 ? _slots_28_io_out_uop_xcpt_ae_if : _slots_27_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_61
         ? _slots_29_io_out_uop_xcpt_ma_if
         : _GEN_60 ? _slots_28_io_out_uop_xcpt_ma_if : _slots_27_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_61
         ? _slots_29_io_out_uop_bp_debug_if
         : _GEN_60 ? _slots_28_io_out_uop_bp_debug_if : _slots_27_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_61
         ? _slots_29_io_out_uop_bp_xcpt_if
         : _GEN_60 ? _slots_28_io_out_uop_bp_xcpt_if : _slots_27_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_61
         ? _slots_29_io_out_uop_debug_fsrc
         : _GEN_60 ? _slots_28_io_out_uop_debug_fsrc : _slots_27_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_61
         ? _slots_29_io_out_uop_debug_tsrc
         : _GEN_60 ? _slots_28_io_out_uop_debug_tsrc : _slots_27_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_26_io_valid),
    .io_will_be_valid               (_slots_26_io_will_be_valid),
    .io_request                     (_slots_26_io_request),
    .io_out_uop_uopc                (_slots_26_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_26_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_26_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_26_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_26_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_26_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_26_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_26_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_26_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_26_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_26_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_26_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_26_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_26_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_26_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_26_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_26_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_26_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_26_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_26_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_26_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_26_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_26_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_26_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_26_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_26_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_26_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_26_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_26_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_26_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_26_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_26_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_26_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_26_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_26_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_26_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_26_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_26_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_26_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_26_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_26_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_26_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_26_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_26_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_26_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_26_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_26_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_26_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_26_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_26_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_26_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_26_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_26_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_26_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_26_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_26_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_26_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_26_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_26_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_26_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_26_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_26_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_26_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_26_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_26_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_26_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_26_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_26_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_26_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_26_io_uop_uopc),
    .io_uop_inst                    (_slots_26_io_uop_inst),
    .io_uop_debug_inst              (_slots_26_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_26_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_26_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_26_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_26_io_uop_fu_code),
    .io_uop_iw_state                (_slots_26_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_26_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_26_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_26_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_26_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_26_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_26_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_26_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_26_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_26_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_26_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_26_io_uop_pc_lob),
    .io_uop_taken                   (_slots_26_io_uop_taken),
    .io_uop_imm_packed              (_slots_26_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_26_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_26_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_26_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_26_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_26_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_26_io_uop_pdst),
    .io_uop_prs1                    (_slots_26_io_uop_prs1),
    .io_uop_prs2                    (_slots_26_io_uop_prs2),
    .io_uop_prs3                    (_slots_26_io_uop_prs3),
    .io_uop_ppred                   (_slots_26_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_26_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_26_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_26_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_26_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_26_io_uop_stale_pdst),
    .io_uop_exception               (_slots_26_io_uop_exception),
    .io_uop_exc_cause               (_slots_26_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_26_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_26_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_26_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_26_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_26_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_26_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_26_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_26_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_26_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_26_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_26_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_26_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_26_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_26_io_uop_ldst),
    .io_uop_lrs1                    (_slots_26_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_26_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_26_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_26_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_26_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_26_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_26_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_26_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_26_io_uop_fp_val),
    .io_uop_fp_single               (_slots_26_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_26_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_26_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_26_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_26_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_26_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_26_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_26_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_27 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_27_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_26),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_27_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_63
         ? _slots_30_io_out_uop_uopc
         : _GEN_62 ? _slots_29_io_out_uop_uopc : _slots_28_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_63
         ? _slots_30_io_out_uop_inst
         : _GEN_62 ? _slots_29_io_out_uop_inst : _slots_28_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_63
         ? _slots_30_io_out_uop_debug_inst
         : _GEN_62 ? _slots_29_io_out_uop_debug_inst : _slots_28_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_63
         ? _slots_30_io_out_uop_is_rvc
         : _GEN_62 ? _slots_29_io_out_uop_is_rvc : _slots_28_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_63
         ? _slots_30_io_out_uop_debug_pc
         : _GEN_62 ? _slots_29_io_out_uop_debug_pc : _slots_28_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_63
         ? _slots_30_io_out_uop_iq_type
         : _GEN_62 ? _slots_29_io_out_uop_iq_type : _slots_28_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_63
         ? _slots_30_io_out_uop_fu_code
         : _GEN_62 ? _slots_29_io_out_uop_fu_code : _slots_28_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_63
         ? _slots_30_io_out_uop_iw_state
         : _GEN_62 ? _slots_29_io_out_uop_iw_state : _slots_28_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_63
         ? _slots_30_io_out_uop_iw_p1_poisoned
         : _GEN_62
             ? _slots_29_io_out_uop_iw_p1_poisoned
             : _slots_28_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_63
         ? _slots_30_io_out_uop_iw_p2_poisoned
         : _GEN_62
             ? _slots_29_io_out_uop_iw_p2_poisoned
             : _slots_28_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_63
         ? _slots_30_io_out_uop_is_br
         : _GEN_62 ? _slots_29_io_out_uop_is_br : _slots_28_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_63
         ? _slots_30_io_out_uop_is_jalr
         : _GEN_62 ? _slots_29_io_out_uop_is_jalr : _slots_28_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_63
         ? _slots_30_io_out_uop_is_jal
         : _GEN_62 ? _slots_29_io_out_uop_is_jal : _slots_28_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_63
         ? _slots_30_io_out_uop_is_sfb
         : _GEN_62 ? _slots_29_io_out_uop_is_sfb : _slots_28_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_63
         ? _slots_30_io_out_uop_br_mask
         : _GEN_62 ? _slots_29_io_out_uop_br_mask : _slots_28_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_63
         ? _slots_30_io_out_uop_br_tag
         : _GEN_62 ? _slots_29_io_out_uop_br_tag : _slots_28_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_63
         ? _slots_30_io_out_uop_ftq_idx
         : _GEN_62 ? _slots_29_io_out_uop_ftq_idx : _slots_28_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_63
         ? _slots_30_io_out_uop_edge_inst
         : _GEN_62 ? _slots_29_io_out_uop_edge_inst : _slots_28_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_63
         ? _slots_30_io_out_uop_pc_lob
         : _GEN_62 ? _slots_29_io_out_uop_pc_lob : _slots_28_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_63
         ? _slots_30_io_out_uop_taken
         : _GEN_62 ? _slots_29_io_out_uop_taken : _slots_28_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_63
         ? _slots_30_io_out_uop_imm_packed
         : _GEN_62 ? _slots_29_io_out_uop_imm_packed : _slots_28_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_63
         ? _slots_30_io_out_uop_csr_addr
         : _GEN_62 ? _slots_29_io_out_uop_csr_addr : _slots_28_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_63
         ? _slots_30_io_out_uop_rob_idx
         : _GEN_62 ? _slots_29_io_out_uop_rob_idx : _slots_28_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_63
         ? _slots_30_io_out_uop_ldq_idx
         : _GEN_62 ? _slots_29_io_out_uop_ldq_idx : _slots_28_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_63
         ? _slots_30_io_out_uop_stq_idx
         : _GEN_62 ? _slots_29_io_out_uop_stq_idx : _slots_28_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_63
         ? _slots_30_io_out_uop_rxq_idx
         : _GEN_62 ? _slots_29_io_out_uop_rxq_idx : _slots_28_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_63
         ? _slots_30_io_out_uop_pdst
         : _GEN_62 ? _slots_29_io_out_uop_pdst : _slots_28_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_63
         ? _slots_30_io_out_uop_prs1
         : _GEN_62 ? _slots_29_io_out_uop_prs1 : _slots_28_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_63
         ? _slots_30_io_out_uop_prs2
         : _GEN_62 ? _slots_29_io_out_uop_prs2 : _slots_28_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_63
         ? _slots_30_io_out_uop_prs3
         : _GEN_62 ? _slots_29_io_out_uop_prs3 : _slots_28_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_63
         ? _slots_30_io_out_uop_ppred
         : _GEN_62 ? _slots_29_io_out_uop_ppred : _slots_28_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_63
         ? _slots_30_io_out_uop_prs1_busy
         : _GEN_62 ? _slots_29_io_out_uop_prs1_busy : _slots_28_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_63
         ? _slots_30_io_out_uop_prs2_busy
         : _GEN_62 ? _slots_29_io_out_uop_prs2_busy : _slots_28_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_63
         ? _slots_30_io_out_uop_prs3_busy
         : _GEN_62 ? _slots_29_io_out_uop_prs3_busy : _slots_28_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_63
         ? _slots_30_io_out_uop_ppred_busy
         : _GEN_62 ? _slots_29_io_out_uop_ppred_busy : _slots_28_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_63
         ? _slots_30_io_out_uop_stale_pdst
         : _GEN_62 ? _slots_29_io_out_uop_stale_pdst : _slots_28_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_63
         ? _slots_30_io_out_uop_exception
         : _GEN_62 ? _slots_29_io_out_uop_exception : _slots_28_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_63
         ? _slots_30_io_out_uop_exc_cause
         : _GEN_62 ? _slots_29_io_out_uop_exc_cause : _slots_28_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_63
         ? _slots_30_io_out_uop_bypassable
         : _GEN_62 ? _slots_29_io_out_uop_bypassable : _slots_28_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_63
         ? _slots_30_io_out_uop_mem_cmd
         : _GEN_62 ? _slots_29_io_out_uop_mem_cmd : _slots_28_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_63
         ? _slots_30_io_out_uop_mem_size
         : _GEN_62 ? _slots_29_io_out_uop_mem_size : _slots_28_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_63
         ? _slots_30_io_out_uop_mem_signed
         : _GEN_62 ? _slots_29_io_out_uop_mem_signed : _slots_28_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_63
         ? _slots_30_io_out_uop_is_fence
         : _GEN_62 ? _slots_29_io_out_uop_is_fence : _slots_28_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_63
         ? _slots_30_io_out_uop_is_fencei
         : _GEN_62 ? _slots_29_io_out_uop_is_fencei : _slots_28_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_63
         ? _slots_30_io_out_uop_is_amo
         : _GEN_62 ? _slots_29_io_out_uop_is_amo : _slots_28_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_63
         ? _slots_30_io_out_uop_uses_ldq
         : _GEN_62 ? _slots_29_io_out_uop_uses_ldq : _slots_28_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_63
         ? _slots_30_io_out_uop_uses_stq
         : _GEN_62 ? _slots_29_io_out_uop_uses_stq : _slots_28_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_63
         ? _slots_30_io_out_uop_is_sys_pc2epc
         : _GEN_62
             ? _slots_29_io_out_uop_is_sys_pc2epc
             : _slots_28_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_63
         ? _slots_30_io_out_uop_is_unique
         : _GEN_62 ? _slots_29_io_out_uop_is_unique : _slots_28_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_63
         ? _slots_30_io_out_uop_flush_on_commit
         : _GEN_62
             ? _slots_29_io_out_uop_flush_on_commit
             : _slots_28_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_63
         ? _slots_30_io_out_uop_ldst_is_rs1
         : _GEN_62 ? _slots_29_io_out_uop_ldst_is_rs1 : _slots_28_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_63
         ? _slots_30_io_out_uop_ldst
         : _GEN_62 ? _slots_29_io_out_uop_ldst : _slots_28_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_63
         ? _slots_30_io_out_uop_lrs1
         : _GEN_62 ? _slots_29_io_out_uop_lrs1 : _slots_28_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_63
         ? _slots_30_io_out_uop_lrs2
         : _GEN_62 ? _slots_29_io_out_uop_lrs2 : _slots_28_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_63
         ? _slots_30_io_out_uop_lrs3
         : _GEN_62 ? _slots_29_io_out_uop_lrs3 : _slots_28_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_63
         ? _slots_30_io_out_uop_ldst_val
         : _GEN_62 ? _slots_29_io_out_uop_ldst_val : _slots_28_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_63
         ? _slots_30_io_out_uop_dst_rtype
         : _GEN_62 ? _slots_29_io_out_uop_dst_rtype : _slots_28_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_63
         ? _slots_30_io_out_uop_lrs1_rtype
         : _GEN_62 ? _slots_29_io_out_uop_lrs1_rtype : _slots_28_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_63
         ? _slots_30_io_out_uop_lrs2_rtype
         : _GEN_62 ? _slots_29_io_out_uop_lrs2_rtype : _slots_28_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_63
         ? _slots_30_io_out_uop_frs3_en
         : _GEN_62 ? _slots_29_io_out_uop_frs3_en : _slots_28_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_63
         ? _slots_30_io_out_uop_fp_val
         : _GEN_62 ? _slots_29_io_out_uop_fp_val : _slots_28_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_63
         ? _slots_30_io_out_uop_fp_single
         : _GEN_62 ? _slots_29_io_out_uop_fp_single : _slots_28_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_63
         ? _slots_30_io_out_uop_xcpt_pf_if
         : _GEN_62 ? _slots_29_io_out_uop_xcpt_pf_if : _slots_28_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_63
         ? _slots_30_io_out_uop_xcpt_ae_if
         : _GEN_62 ? _slots_29_io_out_uop_xcpt_ae_if : _slots_28_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_63
         ? _slots_30_io_out_uop_xcpt_ma_if
         : _GEN_62 ? _slots_29_io_out_uop_xcpt_ma_if : _slots_28_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_63
         ? _slots_30_io_out_uop_bp_debug_if
         : _GEN_62 ? _slots_29_io_out_uop_bp_debug_if : _slots_28_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_63
         ? _slots_30_io_out_uop_bp_xcpt_if
         : _GEN_62 ? _slots_29_io_out_uop_bp_xcpt_if : _slots_28_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_63
         ? _slots_30_io_out_uop_debug_fsrc
         : _GEN_62 ? _slots_29_io_out_uop_debug_fsrc : _slots_28_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_63
         ? _slots_30_io_out_uop_debug_tsrc
         : _GEN_62 ? _slots_29_io_out_uop_debug_tsrc : _slots_28_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_27_io_valid),
    .io_will_be_valid               (_slots_27_io_will_be_valid),
    .io_request                     (_slots_27_io_request),
    .io_out_uop_uopc                (_slots_27_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_27_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_27_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_27_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_27_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_27_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_27_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_27_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_27_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_27_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_27_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_27_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_27_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_27_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_27_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_27_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_27_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_27_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_27_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_27_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_27_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_27_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_27_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_27_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_27_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_27_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_27_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_27_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_27_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_27_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_27_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_27_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_27_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_27_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_27_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_27_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_27_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_27_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_27_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_27_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_27_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_27_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_27_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_27_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_27_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_27_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_27_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_27_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_27_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_27_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_27_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_27_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_27_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_27_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_27_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_27_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_27_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_27_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_27_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_27_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_27_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_27_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_27_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_27_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_27_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_27_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_27_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_27_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_27_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_27_io_uop_uopc),
    .io_uop_inst                    (_slots_27_io_uop_inst),
    .io_uop_debug_inst              (_slots_27_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_27_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_27_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_27_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_27_io_uop_fu_code),
    .io_uop_iw_state                (_slots_27_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_27_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_27_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_27_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_27_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_27_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_27_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_27_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_27_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_27_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_27_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_27_io_uop_pc_lob),
    .io_uop_taken                   (_slots_27_io_uop_taken),
    .io_uop_imm_packed              (_slots_27_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_27_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_27_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_27_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_27_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_27_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_27_io_uop_pdst),
    .io_uop_prs1                    (_slots_27_io_uop_prs1),
    .io_uop_prs2                    (_slots_27_io_uop_prs2),
    .io_uop_prs3                    (_slots_27_io_uop_prs3),
    .io_uop_ppred                   (_slots_27_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_27_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_27_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_27_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_27_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_27_io_uop_stale_pdst),
    .io_uop_exception               (_slots_27_io_uop_exception),
    .io_uop_exc_cause               (_slots_27_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_27_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_27_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_27_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_27_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_27_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_27_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_27_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_27_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_27_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_27_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_27_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_27_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_27_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_27_io_uop_ldst),
    .io_uop_lrs1                    (_slots_27_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_27_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_27_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_27_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_27_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_27_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_27_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_27_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_27_io_uop_fp_val),
    .io_uop_fp_single               (_slots_27_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_27_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_27_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_27_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_27_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_27_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_27_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_27_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_28 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_28_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_27),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_28_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_65
         ? _slots_31_io_out_uop_uopc
         : _GEN_64 ? _slots_30_io_out_uop_uopc : _slots_29_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_65
         ? _slots_31_io_out_uop_inst
         : _GEN_64 ? _slots_30_io_out_uop_inst : _slots_29_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_65
         ? _slots_31_io_out_uop_debug_inst
         : _GEN_64 ? _slots_30_io_out_uop_debug_inst : _slots_29_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_65
         ? _slots_31_io_out_uop_is_rvc
         : _GEN_64 ? _slots_30_io_out_uop_is_rvc : _slots_29_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_65
         ? _slots_31_io_out_uop_debug_pc
         : _GEN_64 ? _slots_30_io_out_uop_debug_pc : _slots_29_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_65
         ? _slots_31_io_out_uop_iq_type
         : _GEN_64 ? _slots_30_io_out_uop_iq_type : _slots_29_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_65
         ? _slots_31_io_out_uop_fu_code
         : _GEN_64 ? _slots_30_io_out_uop_fu_code : _slots_29_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_65
         ? _slots_31_io_out_uop_iw_state
         : _GEN_64 ? _slots_30_io_out_uop_iw_state : _slots_29_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p1_poisoned
      (_GEN_65
         ? _slots_31_io_out_uop_iw_p1_poisoned
         : _GEN_64
             ? _slots_30_io_out_uop_iw_p1_poisoned
             : _slots_29_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (_GEN_65
         ? _slots_31_io_out_uop_iw_p2_poisoned
         : _GEN_64
             ? _slots_30_io_out_uop_iw_p2_poisoned
             : _slots_29_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_65
         ? _slots_31_io_out_uop_is_br
         : _GEN_64 ? _slots_30_io_out_uop_is_br : _slots_29_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_65
         ? _slots_31_io_out_uop_is_jalr
         : _GEN_64 ? _slots_30_io_out_uop_is_jalr : _slots_29_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_65
         ? _slots_31_io_out_uop_is_jal
         : _GEN_64 ? _slots_30_io_out_uop_is_jal : _slots_29_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_65
         ? _slots_31_io_out_uop_is_sfb
         : _GEN_64 ? _slots_30_io_out_uop_is_sfb : _slots_29_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_65
         ? _slots_31_io_out_uop_br_mask
         : _GEN_64 ? _slots_30_io_out_uop_br_mask : _slots_29_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_65
         ? _slots_31_io_out_uop_br_tag
         : _GEN_64 ? _slots_30_io_out_uop_br_tag : _slots_29_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_65
         ? _slots_31_io_out_uop_ftq_idx
         : _GEN_64 ? _slots_30_io_out_uop_ftq_idx : _slots_29_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_65
         ? _slots_31_io_out_uop_edge_inst
         : _GEN_64 ? _slots_30_io_out_uop_edge_inst : _slots_29_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_65
         ? _slots_31_io_out_uop_pc_lob
         : _GEN_64 ? _slots_30_io_out_uop_pc_lob : _slots_29_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_65
         ? _slots_31_io_out_uop_taken
         : _GEN_64 ? _slots_30_io_out_uop_taken : _slots_29_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_65
         ? _slots_31_io_out_uop_imm_packed
         : _GEN_64 ? _slots_30_io_out_uop_imm_packed : _slots_29_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_65
         ? _slots_31_io_out_uop_csr_addr
         : _GEN_64 ? _slots_30_io_out_uop_csr_addr : _slots_29_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_65
         ? _slots_31_io_out_uop_rob_idx
         : _GEN_64 ? _slots_30_io_out_uop_rob_idx : _slots_29_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_65
         ? _slots_31_io_out_uop_ldq_idx
         : _GEN_64 ? _slots_30_io_out_uop_ldq_idx : _slots_29_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_65
         ? _slots_31_io_out_uop_stq_idx
         : _GEN_64 ? _slots_30_io_out_uop_stq_idx : _slots_29_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_65
         ? _slots_31_io_out_uop_rxq_idx
         : _GEN_64 ? _slots_30_io_out_uop_rxq_idx : _slots_29_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_65
         ? _slots_31_io_out_uop_pdst
         : _GEN_64 ? _slots_30_io_out_uop_pdst : _slots_29_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_65
         ? _slots_31_io_out_uop_prs1
         : _GEN_64 ? _slots_30_io_out_uop_prs1 : _slots_29_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_65
         ? _slots_31_io_out_uop_prs2
         : _GEN_64 ? _slots_30_io_out_uop_prs2 : _slots_29_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_65
         ? _slots_31_io_out_uop_prs3
         : _GEN_64 ? _slots_30_io_out_uop_prs3 : _slots_29_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_65
         ? _slots_31_io_out_uop_ppred
         : _GEN_64 ? _slots_30_io_out_uop_ppred : _slots_29_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1_busy
      (_GEN_65
         ? _slots_31_io_out_uop_prs1_busy
         : _GEN_64 ? _slots_30_io_out_uop_prs1_busy : _slots_29_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_65
         ? _slots_31_io_out_uop_prs2_busy
         : _GEN_64 ? _slots_30_io_out_uop_prs2_busy : _slots_29_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3_busy
      (_GEN_65
         ? _slots_31_io_out_uop_prs3_busy
         : _GEN_64 ? _slots_30_io_out_uop_prs3_busy : _slots_29_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (_GEN_65
         ? _slots_31_io_out_uop_ppred_busy
         : _GEN_64 ? _slots_30_io_out_uop_ppred_busy : _slots_29_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_65
         ? _slots_31_io_out_uop_stale_pdst
         : _GEN_64 ? _slots_30_io_out_uop_stale_pdst : _slots_29_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_65
         ? _slots_31_io_out_uop_exception
         : _GEN_64 ? _slots_30_io_out_uop_exception : _slots_29_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_65
         ? _slots_31_io_out_uop_exc_cause
         : _GEN_64 ? _slots_30_io_out_uop_exc_cause : _slots_29_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_65
         ? _slots_31_io_out_uop_bypassable
         : _GEN_64 ? _slots_30_io_out_uop_bypassable : _slots_29_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_65
         ? _slots_31_io_out_uop_mem_cmd
         : _GEN_64 ? _slots_30_io_out_uop_mem_cmd : _slots_29_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_65
         ? _slots_31_io_out_uop_mem_size
         : _GEN_64 ? _slots_30_io_out_uop_mem_size : _slots_29_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_65
         ? _slots_31_io_out_uop_mem_signed
         : _GEN_64 ? _slots_30_io_out_uop_mem_signed : _slots_29_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_65
         ? _slots_31_io_out_uop_is_fence
         : _GEN_64 ? _slots_30_io_out_uop_is_fence : _slots_29_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_65
         ? _slots_31_io_out_uop_is_fencei
         : _GEN_64 ? _slots_30_io_out_uop_is_fencei : _slots_29_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_65
         ? _slots_31_io_out_uop_is_amo
         : _GEN_64 ? _slots_30_io_out_uop_is_amo : _slots_29_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_65
         ? _slots_31_io_out_uop_uses_ldq
         : _GEN_64 ? _slots_30_io_out_uop_uses_ldq : _slots_29_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_65
         ? _slots_31_io_out_uop_uses_stq
         : _GEN_64 ? _slots_30_io_out_uop_uses_stq : _slots_29_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_65
         ? _slots_31_io_out_uop_is_sys_pc2epc
         : _GEN_64
             ? _slots_30_io_out_uop_is_sys_pc2epc
             : _slots_29_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_65
         ? _slots_31_io_out_uop_is_unique
         : _GEN_64 ? _slots_30_io_out_uop_is_unique : _slots_29_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_65
         ? _slots_31_io_out_uop_flush_on_commit
         : _GEN_64
             ? _slots_30_io_out_uop_flush_on_commit
             : _slots_29_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_65
         ? _slots_31_io_out_uop_ldst_is_rs1
         : _GEN_64 ? _slots_30_io_out_uop_ldst_is_rs1 : _slots_29_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_65
         ? _slots_31_io_out_uop_ldst
         : _GEN_64 ? _slots_30_io_out_uop_ldst : _slots_29_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_65
         ? _slots_31_io_out_uop_lrs1
         : _GEN_64 ? _slots_30_io_out_uop_lrs1 : _slots_29_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_65
         ? _slots_31_io_out_uop_lrs2
         : _GEN_64 ? _slots_30_io_out_uop_lrs2 : _slots_29_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_65
         ? _slots_31_io_out_uop_lrs3
         : _GEN_64 ? _slots_30_io_out_uop_lrs3 : _slots_29_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_65
         ? _slots_31_io_out_uop_ldst_val
         : _GEN_64 ? _slots_30_io_out_uop_ldst_val : _slots_29_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_65
         ? _slots_31_io_out_uop_dst_rtype
         : _GEN_64 ? _slots_30_io_out_uop_dst_rtype : _slots_29_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_65
         ? _slots_31_io_out_uop_lrs1_rtype
         : _GEN_64 ? _slots_30_io_out_uop_lrs1_rtype : _slots_29_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_65
         ? _slots_31_io_out_uop_lrs2_rtype
         : _GEN_64 ? _slots_30_io_out_uop_lrs2_rtype : _slots_29_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_frs3_en
      (_GEN_65
         ? _slots_31_io_out_uop_frs3_en
         : _GEN_64 ? _slots_30_io_out_uop_frs3_en : _slots_29_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_65
         ? _slots_31_io_out_uop_fp_val
         : _GEN_64 ? _slots_30_io_out_uop_fp_val : _slots_29_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_65
         ? _slots_31_io_out_uop_fp_single
         : _GEN_64 ? _slots_30_io_out_uop_fp_single : _slots_29_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_65
         ? _slots_31_io_out_uop_xcpt_pf_if
         : _GEN_64 ? _slots_30_io_out_uop_xcpt_pf_if : _slots_29_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_65
         ? _slots_31_io_out_uop_xcpt_ae_if
         : _GEN_64 ? _slots_30_io_out_uop_xcpt_ae_if : _slots_29_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_65
         ? _slots_31_io_out_uop_xcpt_ma_if
         : _GEN_64 ? _slots_30_io_out_uop_xcpt_ma_if : _slots_29_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_65
         ? _slots_31_io_out_uop_bp_debug_if
         : _GEN_64 ? _slots_30_io_out_uop_bp_debug_if : _slots_29_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_65
         ? _slots_31_io_out_uop_bp_xcpt_if
         : _GEN_64 ? _slots_30_io_out_uop_bp_xcpt_if : _slots_29_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_65
         ? _slots_31_io_out_uop_debug_fsrc
         : _GEN_64 ? _slots_30_io_out_uop_debug_fsrc : _slots_29_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_65
         ? _slots_31_io_out_uop_debug_tsrc
         : _GEN_64 ? _slots_30_io_out_uop_debug_tsrc : _slots_29_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_28_io_valid),
    .io_will_be_valid               (_slots_28_io_will_be_valid),
    .io_request                     (_slots_28_io_request),
    .io_out_uop_uopc                (_slots_28_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_28_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_28_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_28_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_28_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_28_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_28_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_28_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_28_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_28_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_28_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_28_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_28_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_28_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_28_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_28_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_28_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_28_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_28_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_28_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_28_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_28_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_28_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_28_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_28_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_28_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_28_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_28_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_28_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_28_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_28_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_28_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_28_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_28_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_28_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_28_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_28_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_28_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_28_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_28_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_28_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_28_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_28_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_28_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_28_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_28_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_28_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_28_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_28_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_28_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_28_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_28_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_28_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_28_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_28_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_28_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_28_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_28_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_28_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_28_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_28_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_28_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_28_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_28_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_28_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_28_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_28_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_28_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_28_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_28_io_uop_uopc),
    .io_uop_inst                    (_slots_28_io_uop_inst),
    .io_uop_debug_inst              (_slots_28_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_28_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_28_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_28_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_28_io_uop_fu_code),
    .io_uop_iw_state                (_slots_28_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_28_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_28_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_28_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_28_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_28_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_28_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_28_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_28_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_28_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_28_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_28_io_uop_pc_lob),
    .io_uop_taken                   (_slots_28_io_uop_taken),
    .io_uop_imm_packed              (_slots_28_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_28_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_28_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_28_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_28_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_28_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_28_io_uop_pdst),
    .io_uop_prs1                    (_slots_28_io_uop_prs1),
    .io_uop_prs2                    (_slots_28_io_uop_prs2),
    .io_uop_prs3                    (_slots_28_io_uop_prs3),
    .io_uop_ppred                   (_slots_28_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_28_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_28_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_28_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_28_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_28_io_uop_stale_pdst),
    .io_uop_exception               (_slots_28_io_uop_exception),
    .io_uop_exc_cause               (_slots_28_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_28_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_28_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_28_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_28_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_28_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_28_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_28_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_28_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_28_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_28_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_28_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_28_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_28_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_28_io_uop_ldst),
    .io_uop_lrs1                    (_slots_28_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_28_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_28_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_28_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_28_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_28_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_28_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_28_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_28_io_uop_fp_val),
    .io_uop_fp_single               (_slots_28_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_28_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_28_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_28_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_28_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_28_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_28_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_28_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_29 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_29_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_28),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_29_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_67
         ? io_dis_uops_0_bits_uopc
         : _GEN_66 ? _slots_31_io_out_uop_uopc : _slots_30_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_67
         ? io_dis_uops_0_bits_inst
         : _GEN_66 ? _slots_31_io_out_uop_inst : _slots_30_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_67
         ? io_dis_uops_0_bits_debug_inst
         : _GEN_66 ? _slots_31_io_out_uop_debug_inst : _slots_30_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_67
         ? io_dis_uops_0_bits_is_rvc
         : _GEN_66 ? _slots_31_io_out_uop_is_rvc : _slots_30_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_67
         ? io_dis_uops_0_bits_debug_pc
         : _GEN_66 ? _slots_31_io_out_uop_debug_pc : _slots_30_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_67
         ? io_dis_uops_0_bits_iq_type
         : _GEN_66 ? _slots_31_io_out_uop_iq_type : _slots_30_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_67
         ? io_dis_uops_0_bits_fu_code
         : _GEN_66 ? _slots_31_io_out_uop_fu_code : _slots_30_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_67
         ? uops_32_iw_state
         : _GEN_66 ? _slots_31_io_out_uop_iw_state : _slots_30_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:123:26, :128:54, :129:30, :153:73
    .io_in_uop_bits_iw_p1_poisoned
      (~_GEN_67
       & (_GEN_66
            ? _slots_31_io_out_uop_iw_p1_poisoned
            : _slots_30_io_out_uop_iw_p1_poisoned)),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned
      (~_GEN_67
       & (_GEN_66
            ? _slots_31_io_out_uop_iw_p2_poisoned
            : _slots_30_io_out_uop_iw_p2_poisoned)),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_67
         ? io_dis_uops_0_bits_is_br
         : _GEN_66 ? _slots_31_io_out_uop_is_br : _slots_30_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_67
         ? io_dis_uops_0_bits_is_jalr
         : _GEN_66 ? _slots_31_io_out_uop_is_jalr : _slots_30_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_67
         ? io_dis_uops_0_bits_is_jal
         : _GEN_66 ? _slots_31_io_out_uop_is_jal : _slots_30_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_67
         ? io_dis_uops_0_bits_is_sfb
         : _GEN_66 ? _slots_31_io_out_uop_is_sfb : _slots_30_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_67
         ? io_dis_uops_0_bits_br_mask
         : _GEN_66 ? _slots_31_io_out_uop_br_mask : _slots_30_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_67
         ? io_dis_uops_0_bits_br_tag
         : _GEN_66 ? _slots_31_io_out_uop_br_tag : _slots_30_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_67
         ? io_dis_uops_0_bits_ftq_idx
         : _GEN_66 ? _slots_31_io_out_uop_ftq_idx : _slots_30_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_67
         ? io_dis_uops_0_bits_edge_inst
         : _GEN_66 ? _slots_31_io_out_uop_edge_inst : _slots_30_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_67
         ? io_dis_uops_0_bits_pc_lob
         : _GEN_66 ? _slots_31_io_out_uop_pc_lob : _slots_30_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_67
         ? io_dis_uops_0_bits_taken
         : _GEN_66 ? _slots_31_io_out_uop_taken : _slots_30_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_67
         ? io_dis_uops_0_bits_imm_packed
         : _GEN_66 ? _slots_31_io_out_uop_imm_packed : _slots_30_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_67
         ? io_dis_uops_0_bits_csr_addr
         : _GEN_66 ? _slots_31_io_out_uop_csr_addr : _slots_30_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_67
         ? io_dis_uops_0_bits_rob_idx
         : _GEN_66 ? _slots_31_io_out_uop_rob_idx : _slots_30_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_67
         ? io_dis_uops_0_bits_ldq_idx
         : _GEN_66 ? _slots_31_io_out_uop_ldq_idx : _slots_30_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_67
         ? io_dis_uops_0_bits_stq_idx
         : _GEN_66 ? _slots_31_io_out_uop_stq_idx : _slots_30_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_67
         ? io_dis_uops_0_bits_rxq_idx
         : _GEN_66 ? _slots_31_io_out_uop_rxq_idx : _slots_30_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_67
         ? io_dis_uops_0_bits_pdst
         : _GEN_66 ? _slots_31_io_out_uop_pdst : _slots_30_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_67
         ? io_dis_uops_0_bits_prs1
         : _GEN_66 ? _slots_31_io_out_uop_prs1 : _slots_30_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_67
         ? io_dis_uops_0_bits_prs2
         : _GEN_66 ? _slots_31_io_out_uop_prs2 : _slots_30_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_67
         ? io_dis_uops_0_bits_prs3
         : _GEN_66 ? _slots_31_io_out_uop_prs3 : _slots_30_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred
      (_GEN_67
         ? 5'h0
         : _GEN_66 ? _slots_31_io_out_uop_ppred : _slots_30_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73, :154:28
    .io_in_uop_bits_prs1_busy
      (_GEN_67
         ? io_dis_uops_0_bits_prs1_busy
         : _GEN_66 ? _slots_31_io_out_uop_prs1_busy : _slots_30_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_67
         ? uops_32_prs2_busy
         : _GEN_66 ? _slots_31_io_out_uop_prs2_busy : _slots_30_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:120:17, :128:54, :131:102, :153:73
    .io_in_uop_bits_prs3_busy
      (~_GEN_67
       & (_GEN_66 ? _slots_31_io_out_uop_prs3_busy : _slots_30_io_out_uop_prs3_busy)),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy
      (~_GEN_67
       & (_GEN_66 ? _slots_31_io_out_uop_ppred_busy : _slots_30_io_out_uop_ppred_busy)),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_67
         ? io_dis_uops_0_bits_stale_pdst
         : _GEN_66 ? _slots_31_io_out_uop_stale_pdst : _slots_30_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_67
         ? io_dis_uops_0_bits_exception
         : _GEN_66 ? _slots_31_io_out_uop_exception : _slots_30_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_67
         ? io_dis_uops_0_bits_exc_cause
         : _GEN_66 ? _slots_31_io_out_uop_exc_cause : _slots_30_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_67
         ? io_dis_uops_0_bits_bypassable
         : _GEN_66 ? _slots_31_io_out_uop_bypassable : _slots_30_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_67
         ? io_dis_uops_0_bits_mem_cmd
         : _GEN_66 ? _slots_31_io_out_uop_mem_cmd : _slots_30_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_67
         ? io_dis_uops_0_bits_mem_size
         : _GEN_66 ? _slots_31_io_out_uop_mem_size : _slots_30_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_67
         ? io_dis_uops_0_bits_mem_signed
         : _GEN_66 ? _slots_31_io_out_uop_mem_signed : _slots_30_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_67
         ? io_dis_uops_0_bits_is_fence
         : _GEN_66 ? _slots_31_io_out_uop_is_fence : _slots_30_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_67
         ? io_dis_uops_0_bits_is_fencei
         : _GEN_66 ? _slots_31_io_out_uop_is_fencei : _slots_30_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_67
         ? io_dis_uops_0_bits_is_amo
         : _GEN_66 ? _slots_31_io_out_uop_is_amo : _slots_30_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_67
         ? io_dis_uops_0_bits_uses_ldq
         : _GEN_66 ? _slots_31_io_out_uop_uses_ldq : _slots_30_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_67
         ? io_dis_uops_0_bits_uses_stq
         : _GEN_66 ? _slots_31_io_out_uop_uses_stq : _slots_30_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_67
         ? io_dis_uops_0_bits_is_sys_pc2epc
         : _GEN_66
             ? _slots_31_io_out_uop_is_sys_pc2epc
             : _slots_30_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_67
         ? io_dis_uops_0_bits_is_unique
         : _GEN_66 ? _slots_31_io_out_uop_is_unique : _slots_30_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_67
         ? io_dis_uops_0_bits_flush_on_commit
         : _GEN_66
             ? _slots_31_io_out_uop_flush_on_commit
             : _slots_30_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_67
         ? io_dis_uops_0_bits_ldst_is_rs1
         : _GEN_66 ? _slots_31_io_out_uop_ldst_is_rs1 : _slots_30_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_67
         ? io_dis_uops_0_bits_ldst
         : _GEN_66 ? _slots_31_io_out_uop_ldst : _slots_30_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_67
         ? io_dis_uops_0_bits_lrs1
         : _GEN_66 ? _slots_31_io_out_uop_lrs1 : _slots_30_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_67
         ? io_dis_uops_0_bits_lrs2
         : _GEN_66 ? _slots_31_io_out_uop_lrs2 : _slots_30_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_67
         ? io_dis_uops_0_bits_lrs3
         : _GEN_66 ? _slots_31_io_out_uop_lrs3 : _slots_30_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_67
         ? io_dis_uops_0_bits_ldst_val
         : _GEN_66 ? _slots_31_io_out_uop_ldst_val : _slots_30_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_67
         ? io_dis_uops_0_bits_dst_rtype
         : _GEN_66 ? _slots_31_io_out_uop_dst_rtype : _slots_30_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_67
         ? io_dis_uops_0_bits_lrs1_rtype
         : _GEN_66 ? _slots_31_io_out_uop_lrs1_rtype : _slots_30_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_67
         ? uops_32_lrs2_rtype
         : _GEN_66 ? _slots_31_io_out_uop_lrs2_rtype : _slots_30_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:120:17, :128:54, :131:102, :153:73
    .io_in_uop_bits_frs3_en
      (_GEN_67
         ? io_dis_uops_0_bits_frs3_en
         : _GEN_66 ? _slots_31_io_out_uop_frs3_en : _slots_30_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_67
         ? io_dis_uops_0_bits_fp_val
         : _GEN_66 ? _slots_31_io_out_uop_fp_val : _slots_30_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_67
         ? io_dis_uops_0_bits_fp_single
         : _GEN_66 ? _slots_31_io_out_uop_fp_single : _slots_30_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_67
         ? io_dis_uops_0_bits_xcpt_pf_if
         : _GEN_66 ? _slots_31_io_out_uop_xcpt_pf_if : _slots_30_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_67
         ? io_dis_uops_0_bits_xcpt_ae_if
         : _GEN_66 ? _slots_31_io_out_uop_xcpt_ae_if : _slots_30_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_67
         ? io_dis_uops_0_bits_xcpt_ma_if
         : _GEN_66 ? _slots_31_io_out_uop_xcpt_ma_if : _slots_30_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_67
         ? io_dis_uops_0_bits_bp_debug_if
         : _GEN_66 ? _slots_31_io_out_uop_bp_debug_if : _slots_30_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_67
         ? io_dis_uops_0_bits_bp_xcpt_if
         : _GEN_66 ? _slots_31_io_out_uop_bp_xcpt_if : _slots_30_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_67
         ? io_dis_uops_0_bits_debug_fsrc
         : _GEN_66 ? _slots_31_io_out_uop_debug_fsrc : _slots_30_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_67
         ? io_dis_uops_0_bits_debug_tsrc
         : _GEN_66 ? _slots_31_io_out_uop_debug_tsrc : _slots_30_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_29_io_valid),
    .io_will_be_valid               (_slots_29_io_will_be_valid),
    .io_request                     (_slots_29_io_request),
    .io_out_uop_uopc                (_slots_29_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_29_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_29_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_29_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_29_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_29_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_29_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_29_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_29_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_29_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_29_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_29_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_29_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_29_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_29_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_29_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_29_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_29_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_29_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_29_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_29_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_29_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_29_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_29_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_29_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_29_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_29_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_29_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_29_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_29_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_29_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_29_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_29_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_29_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_29_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_29_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_29_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_29_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_29_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_29_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_29_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_29_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_29_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_29_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_29_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_29_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_29_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_29_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_29_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_29_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_29_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_29_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_29_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_29_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_29_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_29_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_29_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_29_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_29_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_29_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_29_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_29_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_29_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_29_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_29_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_29_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_29_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_29_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_29_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_29_io_uop_uopc),
    .io_uop_inst                    (_slots_29_io_uop_inst),
    .io_uop_debug_inst              (_slots_29_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_29_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_29_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_29_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_29_io_uop_fu_code),
    .io_uop_iw_state                (_slots_29_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_29_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_29_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_29_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_29_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_29_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_29_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_29_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_29_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_29_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_29_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_29_io_uop_pc_lob),
    .io_uop_taken                   (_slots_29_io_uop_taken),
    .io_uop_imm_packed              (_slots_29_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_29_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_29_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_29_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_29_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_29_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_29_io_uop_pdst),
    .io_uop_prs1                    (_slots_29_io_uop_prs1),
    .io_uop_prs2                    (_slots_29_io_uop_prs2),
    .io_uop_prs3                    (_slots_29_io_uop_prs3),
    .io_uop_ppred                   (_slots_29_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_29_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_29_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_29_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_29_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_29_io_uop_stale_pdst),
    .io_uop_exception               (_slots_29_io_uop_exception),
    .io_uop_exc_cause               (_slots_29_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_29_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_29_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_29_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_29_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_29_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_29_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_29_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_29_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_29_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_29_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_29_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_29_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_29_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_29_io_uop_ldst),
    .io_uop_lrs1                    (_slots_29_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_29_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_29_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_29_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_29_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_29_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_29_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_29_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_29_io_uop_fp_val),
    .io_uop_fp_single               (_slots_29_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_29_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_29_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_29_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_29_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_29_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_29_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_29_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_30 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_30_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_29),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_30_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_69
         ? io_dis_uops_1_bits_uopc
         : _GEN_68 ? io_dis_uops_0_bits_uopc : _slots_31_io_out_uop_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_inst
      (_GEN_69
         ? io_dis_uops_1_bits_inst
         : _GEN_68 ? io_dis_uops_0_bits_inst : _slots_31_io_out_uop_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_inst
      (_GEN_69
         ? io_dis_uops_1_bits_debug_inst
         : _GEN_68 ? io_dis_uops_0_bits_debug_inst : _slots_31_io_out_uop_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_rvc
      (_GEN_69
         ? io_dis_uops_1_bits_is_rvc
         : _GEN_68 ? io_dis_uops_0_bits_is_rvc : _slots_31_io_out_uop_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_pc
      (_GEN_69
         ? io_dis_uops_1_bits_debug_pc
         : _GEN_68 ? io_dis_uops_0_bits_debug_pc : _slots_31_io_out_uop_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iq_type
      (_GEN_69
         ? io_dis_uops_1_bits_iq_type
         : _GEN_68 ? io_dis_uops_0_bits_iq_type : _slots_31_io_out_uop_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fu_code
      (_GEN_69
         ? io_dis_uops_1_bits_fu_code
         : _GEN_68 ? io_dis_uops_0_bits_fu_code : _slots_31_io_out_uop_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_state
      (_GEN_69
         ? (_GEN_3 ? 2'h2 : 2'h1)
         : _GEN_68 ? uops_32_iw_state : _slots_31_io_out_uop_iw_state),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:123:26, :127:96, :128:54, :129:30, :153:73
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_70 & _slots_31_io_out_uop_iw_p1_poisoned),	// issue-unit-age-ordered.scala:71:48, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_70 & _slots_31_io_out_uop_iw_p2_poisoned),	// issue-unit-age-ordered.scala:71:48, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_br
      (_GEN_69
         ? io_dis_uops_1_bits_is_br
         : _GEN_68 ? io_dis_uops_0_bits_is_br : _slots_31_io_out_uop_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jalr
      (_GEN_69
         ? io_dis_uops_1_bits_is_jalr
         : _GEN_68 ? io_dis_uops_0_bits_is_jalr : _slots_31_io_out_uop_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_jal
      (_GEN_69
         ? io_dis_uops_1_bits_is_jal
         : _GEN_68 ? io_dis_uops_0_bits_is_jal : _slots_31_io_out_uop_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sfb
      (_GEN_69
         ? io_dis_uops_1_bits_is_sfb
         : _GEN_68 ? io_dis_uops_0_bits_is_sfb : _slots_31_io_out_uop_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_mask
      (_GEN_69
         ? io_dis_uops_1_bits_br_mask
         : _GEN_68 ? io_dis_uops_0_bits_br_mask : _slots_31_io_out_uop_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_br_tag
      (_GEN_69
         ? io_dis_uops_1_bits_br_tag
         : _GEN_68 ? io_dis_uops_0_bits_br_tag : _slots_31_io_out_uop_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ftq_idx
      (_GEN_69
         ? io_dis_uops_1_bits_ftq_idx
         : _GEN_68 ? io_dis_uops_0_bits_ftq_idx : _slots_31_io_out_uop_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_edge_inst
      (_GEN_69
         ? io_dis_uops_1_bits_edge_inst
         : _GEN_68 ? io_dis_uops_0_bits_edge_inst : _slots_31_io_out_uop_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pc_lob
      (_GEN_69
         ? io_dis_uops_1_bits_pc_lob
         : _GEN_68 ? io_dis_uops_0_bits_pc_lob : _slots_31_io_out_uop_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_taken
      (_GEN_69
         ? io_dis_uops_1_bits_taken
         : _GEN_68 ? io_dis_uops_0_bits_taken : _slots_31_io_out_uop_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_imm_packed
      (_GEN_69
         ? io_dis_uops_1_bits_imm_packed
         : _GEN_68 ? io_dis_uops_0_bits_imm_packed : _slots_31_io_out_uop_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_csr_addr
      (_GEN_69
         ? io_dis_uops_1_bits_csr_addr
         : _GEN_68 ? io_dis_uops_0_bits_csr_addr : _slots_31_io_out_uop_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rob_idx
      (_GEN_69
         ? io_dis_uops_1_bits_rob_idx
         : _GEN_68 ? io_dis_uops_0_bits_rob_idx : _slots_31_io_out_uop_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldq_idx
      (_GEN_69
         ? io_dis_uops_1_bits_ldq_idx
         : _GEN_68 ? io_dis_uops_0_bits_ldq_idx : _slots_31_io_out_uop_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stq_idx
      (_GEN_69
         ? io_dis_uops_1_bits_stq_idx
         : _GEN_68 ? io_dis_uops_0_bits_stq_idx : _slots_31_io_out_uop_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_rxq_idx
      (_GEN_69
         ? io_dis_uops_1_bits_rxq_idx
         : _GEN_68 ? io_dis_uops_0_bits_rxq_idx : _slots_31_io_out_uop_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_pdst
      (_GEN_69
         ? io_dis_uops_1_bits_pdst
         : _GEN_68 ? io_dis_uops_0_bits_pdst : _slots_31_io_out_uop_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs1
      (_GEN_69
         ? io_dis_uops_1_bits_prs1
         : _GEN_68 ? io_dis_uops_0_bits_prs1 : _slots_31_io_out_uop_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2
      (_GEN_69
         ? io_dis_uops_1_bits_prs2
         : _GEN_68 ? io_dis_uops_0_bits_prs2 : _slots_31_io_out_uop_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs3
      (_GEN_69
         ? io_dis_uops_1_bits_prs3
         : _GEN_68 ? io_dis_uops_0_bits_prs3 : _slots_31_io_out_uop_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred           (_GEN_70 ? 5'h0 : _slots_31_io_out_uop_ppred),	// issue-unit-age-ordered.scala:71:48, :73:37, issue-unit.scala:153:73, :154:28
    .io_in_uop_bits_prs1_busy
      (_GEN_69
         ? io_dis_uops_1_bits_prs1_busy
         : _GEN_68 ? io_dis_uops_0_bits_prs1_busy : _slots_31_io_out_uop_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_prs2_busy
      (_GEN_69
         ? uops_33_prs2_busy
         : _GEN_68 ? uops_32_prs2_busy : _slots_31_io_out_uop_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:120:17, :128:54, :131:102, :153:73
    .io_in_uop_bits_prs3_busy       (~_GEN_70 & _slots_31_io_out_uop_prs3_busy),	// issue-unit-age-ordered.scala:71:48, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ppred_busy      (~_GEN_70 & _slots_31_io_out_uop_ppred_busy),	// issue-unit-age-ordered.scala:71:48, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_stale_pdst
      (_GEN_69
         ? io_dis_uops_1_bits_stale_pdst
         : _GEN_68 ? io_dis_uops_0_bits_stale_pdst : _slots_31_io_out_uop_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exception
      (_GEN_69
         ? io_dis_uops_1_bits_exception
         : _GEN_68 ? io_dis_uops_0_bits_exception : _slots_31_io_out_uop_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_exc_cause
      (_GEN_69
         ? io_dis_uops_1_bits_exc_cause
         : _GEN_68 ? io_dis_uops_0_bits_exc_cause : _slots_31_io_out_uop_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bypassable
      (_GEN_69
         ? io_dis_uops_1_bits_bypassable
         : _GEN_68 ? io_dis_uops_0_bits_bypassable : _slots_31_io_out_uop_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_cmd
      (_GEN_69
         ? io_dis_uops_1_bits_mem_cmd
         : _GEN_68 ? io_dis_uops_0_bits_mem_cmd : _slots_31_io_out_uop_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_size
      (_GEN_69
         ? io_dis_uops_1_bits_mem_size
         : _GEN_68 ? io_dis_uops_0_bits_mem_size : _slots_31_io_out_uop_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_mem_signed
      (_GEN_69
         ? io_dis_uops_1_bits_mem_signed
         : _GEN_68 ? io_dis_uops_0_bits_mem_signed : _slots_31_io_out_uop_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fence
      (_GEN_69
         ? io_dis_uops_1_bits_is_fence
         : _GEN_68 ? io_dis_uops_0_bits_is_fence : _slots_31_io_out_uop_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_fencei
      (_GEN_69
         ? io_dis_uops_1_bits_is_fencei
         : _GEN_68 ? io_dis_uops_0_bits_is_fencei : _slots_31_io_out_uop_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_amo
      (_GEN_69
         ? io_dis_uops_1_bits_is_amo
         : _GEN_68 ? io_dis_uops_0_bits_is_amo : _slots_31_io_out_uop_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_ldq
      (_GEN_69
         ? io_dis_uops_1_bits_uses_ldq
         : _GEN_68 ? io_dis_uops_0_bits_uses_ldq : _slots_31_io_out_uop_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_uses_stq
      (_GEN_69
         ? io_dis_uops_1_bits_uses_stq
         : _GEN_68 ? io_dis_uops_0_bits_uses_stq : _slots_31_io_out_uop_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_69
         ? io_dis_uops_1_bits_is_sys_pc2epc
         : _GEN_68
             ? io_dis_uops_0_bits_is_sys_pc2epc
             : _slots_31_io_out_uop_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_is_unique
      (_GEN_69
         ? io_dis_uops_1_bits_is_unique
         : _GEN_68 ? io_dis_uops_0_bits_is_unique : _slots_31_io_out_uop_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_flush_on_commit
      (_GEN_69
         ? io_dis_uops_1_bits_flush_on_commit
         : _GEN_68
             ? io_dis_uops_0_bits_flush_on_commit
             : _slots_31_io_out_uop_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_69
         ? io_dis_uops_1_bits_ldst_is_rs1
         : _GEN_68 ? io_dis_uops_0_bits_ldst_is_rs1 : _slots_31_io_out_uop_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst
      (_GEN_69
         ? io_dis_uops_1_bits_ldst
         : _GEN_68 ? io_dis_uops_0_bits_ldst : _slots_31_io_out_uop_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1
      (_GEN_69
         ? io_dis_uops_1_bits_lrs1
         : _GEN_68 ? io_dis_uops_0_bits_lrs1 : _slots_31_io_out_uop_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2
      (_GEN_69
         ? io_dis_uops_1_bits_lrs2
         : _GEN_68 ? io_dis_uops_0_bits_lrs2 : _slots_31_io_out_uop_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs3
      (_GEN_69
         ? io_dis_uops_1_bits_lrs3
         : _GEN_68 ? io_dis_uops_0_bits_lrs3 : _slots_31_io_out_uop_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_ldst_val
      (_GEN_69
         ? io_dis_uops_1_bits_ldst_val
         : _GEN_68 ? io_dis_uops_0_bits_ldst_val : _slots_31_io_out_uop_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_dst_rtype
      (_GEN_69
         ? io_dis_uops_1_bits_dst_rtype
         : _GEN_68 ? io_dis_uops_0_bits_dst_rtype : _slots_31_io_out_uop_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs1_rtype
      (_GEN_69
         ? io_dis_uops_1_bits_lrs1_rtype
         : _GEN_68 ? io_dis_uops_0_bits_lrs1_rtype : _slots_31_io_out_uop_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_lrs2_rtype
      (_GEN_69
         ? uops_33_lrs2_rtype
         : _GEN_68 ? uops_32_lrs2_rtype : _slots_31_io_out_uop_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:120:17, :128:54, :131:102, :153:73
    .io_in_uop_bits_frs3_en
      (_GEN_69
         ? io_dis_uops_1_bits_frs3_en
         : _GEN_68 ? io_dis_uops_0_bits_frs3_en : _slots_31_io_out_uop_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_val
      (_GEN_69
         ? io_dis_uops_1_bits_fp_val
         : _GEN_68 ? io_dis_uops_0_bits_fp_val : _slots_31_io_out_uop_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_fp_single
      (_GEN_69
         ? io_dis_uops_1_bits_fp_single
         : _GEN_68 ? io_dis_uops_0_bits_fp_single : _slots_31_io_out_uop_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_69
         ? io_dis_uops_1_bits_xcpt_pf_if
         : _GEN_68 ? io_dis_uops_0_bits_xcpt_pf_if : _slots_31_io_out_uop_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_69
         ? io_dis_uops_1_bits_xcpt_ae_if
         : _GEN_68 ? io_dis_uops_0_bits_xcpt_ae_if : _slots_31_io_out_uop_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_69
         ? io_dis_uops_1_bits_xcpt_ma_if
         : _GEN_68 ? io_dis_uops_0_bits_xcpt_ma_if : _slots_31_io_out_uop_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_debug_if
      (_GEN_69
         ? io_dis_uops_1_bits_bp_debug_if
         : _GEN_68 ? io_dis_uops_0_bits_bp_debug_if : _slots_31_io_out_uop_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_69
         ? io_dis_uops_1_bits_bp_xcpt_if
         : _GEN_68 ? io_dis_uops_0_bits_bp_xcpt_if : _slots_31_io_out_uop_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_fsrc
      (_GEN_69
         ? io_dis_uops_1_bits_debug_fsrc
         : _GEN_68 ? io_dis_uops_0_bits_debug_fsrc : _slots_31_io_out_uop_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_in_uop_bits_debug_tsrc
      (_GEN_69
         ? io_dis_uops_1_bits_debug_tsrc
         : _GEN_68 ? io_dis_uops_0_bits_debug_tsrc : _slots_31_io_out_uop_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:153:73
    .io_valid                       (_slots_30_io_valid),
    .io_will_be_valid               (_slots_30_io_will_be_valid),
    .io_request                     (_slots_30_io_request),
    .io_out_uop_uopc                (_slots_30_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_30_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_30_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_30_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_30_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_30_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_30_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_30_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_30_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_30_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_30_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_30_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_30_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_30_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_30_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_30_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_30_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_30_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_30_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_30_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_30_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_30_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_30_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_30_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_30_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_30_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_30_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_30_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_30_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_30_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_30_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_30_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_30_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_30_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_30_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_30_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_30_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_30_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_30_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_30_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_30_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_30_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_30_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_30_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_30_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_30_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_30_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_30_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_30_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_30_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_30_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_30_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_30_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_30_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_30_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_30_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_30_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_30_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_30_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_30_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_30_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_30_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_30_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_30_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_30_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_30_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_30_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_30_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_30_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_30_io_uop_uopc),
    .io_uop_inst                    (_slots_30_io_uop_inst),
    .io_uop_debug_inst              (_slots_30_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_30_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_30_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_30_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_30_io_uop_fu_code),
    .io_uop_iw_state                (_slots_30_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_30_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_30_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_30_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_30_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_30_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_30_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_30_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_30_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_30_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_30_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_30_io_uop_pc_lob),
    .io_uop_taken                   (_slots_30_io_uop_taken),
    .io_uop_imm_packed              (_slots_30_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_30_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_30_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_30_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_30_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_30_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_30_io_uop_pdst),
    .io_uop_prs1                    (_slots_30_io_uop_prs1),
    .io_uop_prs2                    (_slots_30_io_uop_prs2),
    .io_uop_prs3                    (_slots_30_io_uop_prs3),
    .io_uop_ppred                   (_slots_30_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_30_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_30_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_30_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_30_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_30_io_uop_stale_pdst),
    .io_uop_exception               (_slots_30_io_uop_exception),
    .io_uop_exc_cause               (_slots_30_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_30_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_30_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_30_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_30_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_30_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_30_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_30_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_30_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_30_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_30_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_30_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_30_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_30_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_30_io_uop_ldst),
    .io_uop_lrs1                    (_slots_30_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_30_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_30_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_30_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_30_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_30_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_30_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_30_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_30_io_uop_fp_val),
    .io_uop_fp_single               (_slots_30_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_30_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_30_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_30_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_30_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_30_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_30_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_30_io_uop_debug_tsrc)
  );
  IssueSlot_120 slots_31 (	// issue-unit.scala:153:73
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_31_grant),	// issue-unit-age-ordered.scala:118:76, :119:30
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_30),	// issue-unit-age-ordered.scala:45:37, :46:13, :47:44, :76:49
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid                (issue_slots_31_in_uop_valid),	// issue-unit-age-ordered.scala:71:48, :72:37
    .io_in_uop_bits_uopc
      (_GEN_72
         ? io_dis_uops_2_bits_uopc
         : _GEN_71 ? io_dis_uops_1_bits_uopc : io_dis_uops_0_bits_uopc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_inst
      (_GEN_72
         ? io_dis_uops_2_bits_inst
         : _GEN_71 ? io_dis_uops_1_bits_inst : io_dis_uops_0_bits_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_debug_inst
      (_GEN_72
         ? io_dis_uops_2_bits_debug_inst
         : _GEN_71 ? io_dis_uops_1_bits_debug_inst : io_dis_uops_0_bits_debug_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_rvc
      (_GEN_72
         ? io_dis_uops_2_bits_is_rvc
         : _GEN_71 ? io_dis_uops_1_bits_is_rvc : io_dis_uops_0_bits_is_rvc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_debug_pc
      (_GEN_72
         ? io_dis_uops_2_bits_debug_pc
         : _GEN_71 ? io_dis_uops_1_bits_debug_pc : io_dis_uops_0_bits_debug_pc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_iq_type
      (_GEN_72
         ? io_dis_uops_2_bits_iq_type
         : _GEN_71 ? io_dis_uops_1_bits_iq_type : io_dis_uops_0_bits_iq_type),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_fu_code
      (_GEN_72
         ? io_dis_uops_2_bits_fu_code
         : _GEN_71 ? io_dis_uops_1_bits_fu_code : io_dis_uops_0_bits_fu_code),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_iw_state
      ((_GEN_72 ? _GEN_6 : _GEN_71 ? _GEN_3 : _GEN_0) ? 2'h2 : 2'h1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:123:26, :127:96, :128:54, :129:30
    .io_in_uop_bits_iw_p1_poisoned  (1'h0),
    .io_in_uop_bits_iw_p2_poisoned  (1'h0),
    .io_in_uop_bits_is_br
      (_GEN_72
         ? io_dis_uops_2_bits_is_br
         : _GEN_71 ? io_dis_uops_1_bits_is_br : io_dis_uops_0_bits_is_br),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_jalr
      (_GEN_72
         ? io_dis_uops_2_bits_is_jalr
         : _GEN_71 ? io_dis_uops_1_bits_is_jalr : io_dis_uops_0_bits_is_jalr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_jal
      (_GEN_72
         ? io_dis_uops_2_bits_is_jal
         : _GEN_71 ? io_dis_uops_1_bits_is_jal : io_dis_uops_0_bits_is_jal),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_sfb
      (_GEN_72
         ? io_dis_uops_2_bits_is_sfb
         : _GEN_71 ? io_dis_uops_1_bits_is_sfb : io_dis_uops_0_bits_is_sfb),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_br_mask
      (_GEN_72
         ? io_dis_uops_2_bits_br_mask
         : _GEN_71 ? io_dis_uops_1_bits_br_mask : io_dis_uops_0_bits_br_mask),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_br_tag
      (_GEN_72
         ? io_dis_uops_2_bits_br_tag
         : _GEN_71 ? io_dis_uops_1_bits_br_tag : io_dis_uops_0_bits_br_tag),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_ftq_idx
      (_GEN_72
         ? io_dis_uops_2_bits_ftq_idx
         : _GEN_71 ? io_dis_uops_1_bits_ftq_idx : io_dis_uops_0_bits_ftq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_edge_inst
      (_GEN_72
         ? io_dis_uops_2_bits_edge_inst
         : _GEN_71 ? io_dis_uops_1_bits_edge_inst : io_dis_uops_0_bits_edge_inst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_pc_lob
      (_GEN_72
         ? io_dis_uops_2_bits_pc_lob
         : _GEN_71 ? io_dis_uops_1_bits_pc_lob : io_dis_uops_0_bits_pc_lob),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_taken
      (_GEN_72
         ? io_dis_uops_2_bits_taken
         : _GEN_71 ? io_dis_uops_1_bits_taken : io_dis_uops_0_bits_taken),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_imm_packed
      (_GEN_72
         ? io_dis_uops_2_bits_imm_packed
         : _GEN_71 ? io_dis_uops_1_bits_imm_packed : io_dis_uops_0_bits_imm_packed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_csr_addr
      (_GEN_72
         ? io_dis_uops_2_bits_csr_addr
         : _GEN_71 ? io_dis_uops_1_bits_csr_addr : io_dis_uops_0_bits_csr_addr),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_rob_idx
      (_GEN_72
         ? io_dis_uops_2_bits_rob_idx
         : _GEN_71 ? io_dis_uops_1_bits_rob_idx : io_dis_uops_0_bits_rob_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_ldq_idx
      (_GEN_72
         ? io_dis_uops_2_bits_ldq_idx
         : _GEN_71 ? io_dis_uops_1_bits_ldq_idx : io_dis_uops_0_bits_ldq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_stq_idx
      (_GEN_72
         ? io_dis_uops_2_bits_stq_idx
         : _GEN_71 ? io_dis_uops_1_bits_stq_idx : io_dis_uops_0_bits_stq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_rxq_idx
      (_GEN_72
         ? io_dis_uops_2_bits_rxq_idx
         : _GEN_71 ? io_dis_uops_1_bits_rxq_idx : io_dis_uops_0_bits_rxq_idx),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_pdst
      (_GEN_72
         ? io_dis_uops_2_bits_pdst
         : _GEN_71 ? io_dis_uops_1_bits_pdst : io_dis_uops_0_bits_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_prs1
      (_GEN_72
         ? io_dis_uops_2_bits_prs1
         : _GEN_71 ? io_dis_uops_1_bits_prs1 : io_dis_uops_0_bits_prs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_prs2
      (_GEN_72
         ? io_dis_uops_2_bits_prs2
         : _GEN_71 ? io_dis_uops_1_bits_prs2 : io_dis_uops_0_bits_prs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_prs3
      (_GEN_72
         ? io_dis_uops_2_bits_prs3
         : _GEN_71 ? io_dis_uops_1_bits_prs3 : io_dis_uops_0_bits_prs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_ppred           (5'h0),	// issue-unit.scala:153:73, :154:28
    .io_in_uop_bits_prs1_busy
      (_GEN_72
         ? io_dis_uops_2_bits_prs1_busy
         : _GEN_71 ? io_dis_uops_1_bits_prs1_busy : io_dis_uops_0_bits_prs1_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_prs2_busy
      (_GEN_72
         ? _GEN_7 & io_dis_uops_2_bits_prs2_busy
         : _GEN_71 ? uops_33_prs2_busy : uops_32_prs2_busy),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:120:17, :128:54, :131:102
    .io_in_uop_bits_prs3_busy       (1'h0),
    .io_in_uop_bits_ppred_busy      (1'h0),
    .io_in_uop_bits_stale_pdst
      (_GEN_72
         ? io_dis_uops_2_bits_stale_pdst
         : _GEN_71 ? io_dis_uops_1_bits_stale_pdst : io_dis_uops_0_bits_stale_pdst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_exception
      (_GEN_72
         ? io_dis_uops_2_bits_exception
         : _GEN_71 ? io_dis_uops_1_bits_exception : io_dis_uops_0_bits_exception),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_exc_cause
      (_GEN_72
         ? io_dis_uops_2_bits_exc_cause
         : _GEN_71 ? io_dis_uops_1_bits_exc_cause : io_dis_uops_0_bits_exc_cause),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_bypassable
      (_GEN_72
         ? io_dis_uops_2_bits_bypassable
         : _GEN_71 ? io_dis_uops_1_bits_bypassable : io_dis_uops_0_bits_bypassable),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_mem_cmd
      (_GEN_72
         ? io_dis_uops_2_bits_mem_cmd
         : _GEN_71 ? io_dis_uops_1_bits_mem_cmd : io_dis_uops_0_bits_mem_cmd),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_mem_size
      (_GEN_72
         ? io_dis_uops_2_bits_mem_size
         : _GEN_71 ? io_dis_uops_1_bits_mem_size : io_dis_uops_0_bits_mem_size),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_mem_signed
      (_GEN_72
         ? io_dis_uops_2_bits_mem_signed
         : _GEN_71 ? io_dis_uops_1_bits_mem_signed : io_dis_uops_0_bits_mem_signed),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_fence
      (_GEN_72
         ? io_dis_uops_2_bits_is_fence
         : _GEN_71 ? io_dis_uops_1_bits_is_fence : io_dis_uops_0_bits_is_fence),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_fencei
      (_GEN_72
         ? io_dis_uops_2_bits_is_fencei
         : _GEN_71 ? io_dis_uops_1_bits_is_fencei : io_dis_uops_0_bits_is_fencei),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_amo
      (_GEN_72
         ? io_dis_uops_2_bits_is_amo
         : _GEN_71 ? io_dis_uops_1_bits_is_amo : io_dis_uops_0_bits_is_amo),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_uses_ldq
      (_GEN_72
         ? io_dis_uops_2_bits_uses_ldq
         : _GEN_71 ? io_dis_uops_1_bits_uses_ldq : io_dis_uops_0_bits_uses_ldq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_uses_stq
      (_GEN_72
         ? io_dis_uops_2_bits_uses_stq
         : _GEN_71 ? io_dis_uops_1_bits_uses_stq : io_dis_uops_0_bits_uses_stq),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_sys_pc2epc
      (_GEN_72
         ? io_dis_uops_2_bits_is_sys_pc2epc
         : _GEN_71 ? io_dis_uops_1_bits_is_sys_pc2epc : io_dis_uops_0_bits_is_sys_pc2epc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_is_unique
      (_GEN_72
         ? io_dis_uops_2_bits_is_unique
         : _GEN_71 ? io_dis_uops_1_bits_is_unique : io_dis_uops_0_bits_is_unique),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_flush_on_commit
      (_GEN_72
         ? io_dis_uops_2_bits_flush_on_commit
         : _GEN_71
             ? io_dis_uops_1_bits_flush_on_commit
             : io_dis_uops_0_bits_flush_on_commit),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_ldst_is_rs1
      (_GEN_72
         ? io_dis_uops_2_bits_ldst_is_rs1
         : _GEN_71 ? io_dis_uops_1_bits_ldst_is_rs1 : io_dis_uops_0_bits_ldst_is_rs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_ldst
      (_GEN_72
         ? io_dis_uops_2_bits_ldst
         : _GEN_71 ? io_dis_uops_1_bits_ldst : io_dis_uops_0_bits_ldst),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_lrs1
      (_GEN_72
         ? io_dis_uops_2_bits_lrs1
         : _GEN_71 ? io_dis_uops_1_bits_lrs1 : io_dis_uops_0_bits_lrs1),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_lrs2
      (_GEN_72
         ? io_dis_uops_2_bits_lrs2
         : _GEN_71 ? io_dis_uops_1_bits_lrs2 : io_dis_uops_0_bits_lrs2),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_lrs3
      (_GEN_72
         ? io_dis_uops_2_bits_lrs3
         : _GEN_71 ? io_dis_uops_1_bits_lrs3 : io_dis_uops_0_bits_lrs3),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_ldst_val
      (_GEN_72
         ? io_dis_uops_2_bits_ldst_val
         : _GEN_71 ? io_dis_uops_1_bits_ldst_val : io_dis_uops_0_bits_ldst_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_dst_rtype
      (_GEN_72
         ? io_dis_uops_2_bits_dst_rtype
         : _GEN_71 ? io_dis_uops_1_bits_dst_rtype : io_dis_uops_0_bits_dst_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_lrs1_rtype
      (_GEN_72
         ? io_dis_uops_2_bits_lrs1_rtype
         : _GEN_71 ? io_dis_uops_1_bits_lrs1_rtype : io_dis_uops_0_bits_lrs1_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_lrs2_rtype
      (_GEN_72
         ? (_GEN_7 ? io_dis_uops_2_bits_lrs2_rtype : 2'h2)
         : _GEN_71 ? uops_33_lrs2_rtype : uops_32_lrs2_rtype),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37, issue-unit.scala:120:17, :128:54, :129:30, :131:102
    .io_in_uop_bits_frs3_en
      (_GEN_72
         ? io_dis_uops_2_bits_frs3_en
         : _GEN_71 ? io_dis_uops_1_bits_frs3_en : io_dis_uops_0_bits_frs3_en),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_fp_val
      (_GEN_72
         ? io_dis_uops_2_bits_fp_val
         : _GEN_71 ? io_dis_uops_1_bits_fp_val : io_dis_uops_0_bits_fp_val),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_fp_single
      (_GEN_72
         ? io_dis_uops_2_bits_fp_single
         : _GEN_71 ? io_dis_uops_1_bits_fp_single : io_dis_uops_0_bits_fp_single),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_xcpt_pf_if
      (_GEN_72
         ? io_dis_uops_2_bits_xcpt_pf_if
         : _GEN_71 ? io_dis_uops_1_bits_xcpt_pf_if : io_dis_uops_0_bits_xcpt_pf_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_xcpt_ae_if
      (_GEN_72
         ? io_dis_uops_2_bits_xcpt_ae_if
         : _GEN_71 ? io_dis_uops_1_bits_xcpt_ae_if : io_dis_uops_0_bits_xcpt_ae_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_xcpt_ma_if
      (_GEN_72
         ? io_dis_uops_2_bits_xcpt_ma_if
         : _GEN_71 ? io_dis_uops_1_bits_xcpt_ma_if : io_dis_uops_0_bits_xcpt_ma_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_bp_debug_if
      (_GEN_72
         ? io_dis_uops_2_bits_bp_debug_if
         : _GEN_71 ? io_dis_uops_1_bits_bp_debug_if : io_dis_uops_0_bits_bp_debug_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_bp_xcpt_if
      (_GEN_72
         ? io_dis_uops_2_bits_bp_xcpt_if
         : _GEN_71 ? io_dis_uops_1_bits_bp_xcpt_if : io_dis_uops_0_bits_bp_xcpt_if),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_debug_fsrc
      (_GEN_72
         ? io_dis_uops_2_bits_debug_fsrc
         : _GEN_71 ? io_dis_uops_1_bits_debug_fsrc : io_dis_uops_0_bits_debug_fsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_in_uop_bits_debug_tsrc
      (_GEN_72
         ? io_dis_uops_2_bits_debug_tsrc
         : _GEN_71 ? io_dis_uops_1_bits_debug_tsrc : io_dis_uops_0_bits_debug_tsrc),	// issue-unit-age-ordered.scala:71:{28,48}, :73:37
    .io_valid                       (_slots_31_io_valid),
    .io_will_be_valid               (_slots_31_io_will_be_valid),
    .io_request                     (_slots_31_io_request),
    .io_out_uop_uopc                (_slots_31_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_31_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_31_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_31_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_31_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_31_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_31_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_31_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_31_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_31_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_31_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_31_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_31_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_31_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_31_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_31_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_31_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_31_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_31_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_31_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_31_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_31_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_31_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_31_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_31_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_31_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_31_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_31_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_31_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_31_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_31_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_31_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_31_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_31_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_31_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_31_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_31_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_31_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_31_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_31_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_31_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_31_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_31_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_31_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_31_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_31_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_31_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_31_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_31_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_31_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_31_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_31_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_31_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_31_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_31_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_31_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_31_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_31_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_31_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_31_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_31_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_31_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_31_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_31_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_31_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_31_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_31_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_31_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_31_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_31_io_uop_uopc),
    .io_uop_inst                    (_slots_31_io_uop_inst),
    .io_uop_debug_inst              (_slots_31_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_31_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_31_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_31_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_31_io_uop_fu_code),
    .io_uop_iw_state                (_slots_31_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_31_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_31_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_31_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_31_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_31_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_31_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_31_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_31_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_31_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_31_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_31_io_uop_pc_lob),
    .io_uop_taken                   (_slots_31_io_uop_taken),
    .io_uop_imm_packed              (_slots_31_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_31_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_31_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_31_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_31_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_31_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_31_io_uop_pdst),
    .io_uop_prs1                    (_slots_31_io_uop_prs1),
    .io_uop_prs2                    (_slots_31_io_uop_prs2),
    .io_uop_prs3                    (_slots_31_io_uop_prs3),
    .io_uop_ppred                   (_slots_31_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_31_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_31_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_31_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_31_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_31_io_uop_stale_pdst),
    .io_uop_exception               (_slots_31_io_uop_exception),
    .io_uop_exc_cause               (_slots_31_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_31_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_31_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_31_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_31_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_31_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_31_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_31_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_31_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_31_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_31_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_31_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_31_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_31_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_31_io_uop_ldst),
    .io_uop_lrs1                    (_slots_31_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_31_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_31_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_31_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_31_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_31_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_31_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_31_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_31_io_uop_fp_val),
    .io_uop_fp_single               (_slots_31_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_31_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_31_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_31_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_31_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_31_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_31_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_31_io_uop_debug_tsrc)
  );
  assign io_dis_uops_0_ready = io_dis_uops_0_ready_REG;	// issue-unit-age-ordered.scala:87:36
  assign io_dis_uops_1_ready = io_dis_uops_1_ready_REG;	// issue-unit-age-ordered.scala:87:36
  assign io_dis_uops_2_ready = io_dis_uops_2_ready_REG;	// issue-unit-age-ordered.scala:87:36
  assign io_iss_valids_0 =
    _GEN_344 | _GEN_338 | _GEN_329 | _GEN_320 | _GEN_311 | _GEN_302 | _GEN_293 | _GEN_284
    | _GEN_275 | _GEN_266 | _GEN_257 | _GEN_248 | _GEN_239 | _GEN_230 | _GEN_221
    | _GEN_212 | _GEN_203 | _GEN_194 | _GEN_185 | _GEN_176 | _GEN_167 | _GEN_158
    | _GEN_149 | _GEN_140 | _GEN_131 | _GEN_122 | _GEN_113 | _GEN_104 | _GEN_95 | _GEN_86
    | _GEN_77 | _GEN_73;	// issue-unit-age-ordered.scala:118:{40,56,76}, :120:26
  assign io_iss_valids_1 =
    _GEN_345 | _GEN_340 | _GEN_332 | _GEN_323 | _GEN_314 | _GEN_305 | _GEN_296 | _GEN_287
    | _GEN_278 | _GEN_269 | _GEN_260 | _GEN_251 | _GEN_242 | _GEN_233 | _GEN_224
    | _GEN_215 | _GEN_206 | _GEN_197 | _GEN_188 | _GEN_179 | _GEN_170 | _GEN_161
    | _GEN_152 | _GEN_143 | _GEN_134 | _GEN_125 | _GEN_116 | _GEN_107 | _GEN_98 | _GEN_89
    | _GEN_80 | _GEN_74;	// issue-unit-age-ordered.scala:118:{40,56,76}, :120:26
  assign io_iss_valids_2 =
    _GEN_346 | _GEN_343 | _GEN_335 | _GEN_326 | _GEN_317 | _GEN_308 | _GEN_299 | _GEN_290
    | _GEN_281 | _GEN_272 | _GEN_263 | _GEN_254 | _GEN_245 | _GEN_236 | _GEN_227
    | _GEN_218 | _GEN_209 | _GEN_200 | _GEN_191 | _GEN_182 | _GEN_173 | _GEN_164
    | _GEN_155 | _GEN_146 | _GEN_137 | _GEN_128 | _GEN_119 | _GEN_110 | _GEN_101 | _GEN_92
    | _GEN_83 | _GEN_75;	// issue-unit-age-ordered.scala:118:{40,56,76}, :120:26
  assign io_iss_uops_0_uopc =
    _GEN_344
      ? _slots_31_io_uop_uopc
      : _GEN_338
          ? _slots_30_io_uop_uopc
          : _GEN_329
              ? _slots_29_io_uop_uopc
              : _GEN_320
                  ? _slots_28_io_uop_uopc
                  : _GEN_311
                      ? _slots_27_io_uop_uopc
                      : _GEN_302
                          ? _slots_26_io_uop_uopc
                          : _GEN_293
                              ? _slots_25_io_uop_uopc
                              : _GEN_284
                                  ? _slots_24_io_uop_uopc
                                  : _GEN_275
                                      ? _slots_23_io_uop_uopc
                                      : _GEN_266
                                          ? _slots_22_io_uop_uopc
                                          : _GEN_257
                                              ? _slots_21_io_uop_uopc
                                              : _GEN_248
                                                  ? _slots_20_io_uop_uopc
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_uopc
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_uopc
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_uopc
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_uopc
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_uopc
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_uopc
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_uopc
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_uopc
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_uopc
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_uopc
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_uopc
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_uopc
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_uopc
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_uopc
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_uopc
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_uopc
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_uopc
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_uopc
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_uopc
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_uopc
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_is_rvc =
    _GEN_344
      ? _slots_31_io_uop_is_rvc
      : _GEN_338
          ? _slots_30_io_uop_is_rvc
          : _GEN_329
              ? _slots_29_io_uop_is_rvc
              : _GEN_320
                  ? _slots_28_io_uop_is_rvc
                  : _GEN_311
                      ? _slots_27_io_uop_is_rvc
                      : _GEN_302
                          ? _slots_26_io_uop_is_rvc
                          : _GEN_293
                              ? _slots_25_io_uop_is_rvc
                              : _GEN_284
                                  ? _slots_24_io_uop_is_rvc
                                  : _GEN_275
                                      ? _slots_23_io_uop_is_rvc
                                      : _GEN_266
                                          ? _slots_22_io_uop_is_rvc
                                          : _GEN_257
                                              ? _slots_21_io_uop_is_rvc
                                              : _GEN_248
                                                  ? _slots_20_io_uop_is_rvc
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_is_rvc
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_is_rvc
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_is_rvc
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_is_rvc
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_is_rvc
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_is_rvc
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_is_rvc
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_is_rvc
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_is_rvc
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_is_rvc
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_is_rvc
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_is_rvc
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_is_rvc
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_is_rvc
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_is_rvc
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_is_rvc
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_is_rvc
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_is_rvc
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_is_rvc
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_is_rvc;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_fu_code =
    _GEN_344
      ? _slots_31_io_uop_fu_code
      : _GEN_338
          ? _slots_30_io_uop_fu_code
          : _GEN_329
              ? _slots_29_io_uop_fu_code
              : _GEN_320
                  ? _slots_28_io_uop_fu_code
                  : _GEN_311
                      ? _slots_27_io_uop_fu_code
                      : _GEN_302
                          ? _slots_26_io_uop_fu_code
                          : _GEN_293
                              ? _slots_25_io_uop_fu_code
                              : _GEN_284
                                  ? _slots_24_io_uop_fu_code
                                  : _GEN_275
                                      ? _slots_23_io_uop_fu_code
                                      : _GEN_266
                                          ? _slots_22_io_uop_fu_code
                                          : _GEN_257
                                              ? _slots_21_io_uop_fu_code
                                              : _GEN_248
                                                  ? _slots_20_io_uop_fu_code
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_fu_code
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_fu_code
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_fu_code
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_fu_code
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_fu_code
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_fu_code
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_fu_code
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_fu_code
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_fu_code
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_fu_code
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_fu_code
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_fu_code
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_fu_code
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_fu_code
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_fu_code
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_fu_code
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_fu_code
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_fu_code
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_fu_code
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_fu_code
                                                                                                                                  : 10'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_iw_p1_poisoned =
    _GEN_344
      ? _slots_31_io_uop_iw_p1_poisoned
      : _GEN_338
          ? _slots_30_io_uop_iw_p1_poisoned
          : _GEN_329
              ? _slots_29_io_uop_iw_p1_poisoned
              : _GEN_320
                  ? _slots_28_io_uop_iw_p1_poisoned
                  : _GEN_311
                      ? _slots_27_io_uop_iw_p1_poisoned
                      : _GEN_302
                          ? _slots_26_io_uop_iw_p1_poisoned
                          : _GEN_293
                              ? _slots_25_io_uop_iw_p1_poisoned
                              : _GEN_284
                                  ? _slots_24_io_uop_iw_p1_poisoned
                                  : _GEN_275
                                      ? _slots_23_io_uop_iw_p1_poisoned
                                      : _GEN_266
                                          ? _slots_22_io_uop_iw_p1_poisoned
                                          : _GEN_257
                                              ? _slots_21_io_uop_iw_p1_poisoned
                                              : _GEN_248
                                                  ? _slots_20_io_uop_iw_p1_poisoned
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_iw_p1_poisoned
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_iw_p1_poisoned
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_iw_p1_poisoned
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_iw_p1_poisoned
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_iw_p1_poisoned
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_iw_p1_poisoned
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_iw_p1_poisoned
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_iw_p1_poisoned
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_iw_p1_poisoned
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_iw_p1_poisoned
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_iw_p1_poisoned
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_iw_p1_poisoned
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_iw_p1_poisoned
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_iw_p1_poisoned
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_iw_p1_poisoned
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_iw_p1_poisoned
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_iw_p1_poisoned
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_iw_p1_poisoned
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_iw_p1_poisoned
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_iw_p1_poisoned;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_iw_p2_poisoned =
    _GEN_344
      ? _slots_31_io_uop_iw_p2_poisoned
      : _GEN_338
          ? _slots_30_io_uop_iw_p2_poisoned
          : _GEN_329
              ? _slots_29_io_uop_iw_p2_poisoned
              : _GEN_320
                  ? _slots_28_io_uop_iw_p2_poisoned
                  : _GEN_311
                      ? _slots_27_io_uop_iw_p2_poisoned
                      : _GEN_302
                          ? _slots_26_io_uop_iw_p2_poisoned
                          : _GEN_293
                              ? _slots_25_io_uop_iw_p2_poisoned
                              : _GEN_284
                                  ? _slots_24_io_uop_iw_p2_poisoned
                                  : _GEN_275
                                      ? _slots_23_io_uop_iw_p2_poisoned
                                      : _GEN_266
                                          ? _slots_22_io_uop_iw_p2_poisoned
                                          : _GEN_257
                                              ? _slots_21_io_uop_iw_p2_poisoned
                                              : _GEN_248
                                                  ? _slots_20_io_uop_iw_p2_poisoned
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_iw_p2_poisoned
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_iw_p2_poisoned
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_iw_p2_poisoned
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_iw_p2_poisoned
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_iw_p2_poisoned
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_iw_p2_poisoned
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_iw_p2_poisoned
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_iw_p2_poisoned
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_iw_p2_poisoned
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_iw_p2_poisoned
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_iw_p2_poisoned
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_iw_p2_poisoned
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_iw_p2_poisoned
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_iw_p2_poisoned
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_iw_p2_poisoned
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_iw_p2_poisoned
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_iw_p2_poisoned
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_iw_p2_poisoned
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_iw_p2_poisoned
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_iw_p2_poisoned;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_is_br =
    _GEN_344
      ? _slots_31_io_uop_is_br
      : _GEN_338
          ? _slots_30_io_uop_is_br
          : _GEN_329
              ? _slots_29_io_uop_is_br
              : _GEN_320
                  ? _slots_28_io_uop_is_br
                  : _GEN_311
                      ? _slots_27_io_uop_is_br
                      : _GEN_302
                          ? _slots_26_io_uop_is_br
                          : _GEN_293
                              ? _slots_25_io_uop_is_br
                              : _GEN_284
                                  ? _slots_24_io_uop_is_br
                                  : _GEN_275
                                      ? _slots_23_io_uop_is_br
                                      : _GEN_266
                                          ? _slots_22_io_uop_is_br
                                          : _GEN_257
                                              ? _slots_21_io_uop_is_br
                                              : _GEN_248
                                                  ? _slots_20_io_uop_is_br
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_is_br
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_is_br
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_is_br
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_is_br
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_is_br
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_is_br
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_is_br
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_is_br
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_is_br
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_is_br
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_is_br
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_is_br
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_is_br
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_is_br
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_is_br
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_is_br
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_is_br
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_is_br
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_is_br
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_is_br;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_is_jalr =
    _GEN_344
      ? _slots_31_io_uop_is_jalr
      : _GEN_338
          ? _slots_30_io_uop_is_jalr
          : _GEN_329
              ? _slots_29_io_uop_is_jalr
              : _GEN_320
                  ? _slots_28_io_uop_is_jalr
                  : _GEN_311
                      ? _slots_27_io_uop_is_jalr
                      : _GEN_302
                          ? _slots_26_io_uop_is_jalr
                          : _GEN_293
                              ? _slots_25_io_uop_is_jalr
                              : _GEN_284
                                  ? _slots_24_io_uop_is_jalr
                                  : _GEN_275
                                      ? _slots_23_io_uop_is_jalr
                                      : _GEN_266
                                          ? _slots_22_io_uop_is_jalr
                                          : _GEN_257
                                              ? _slots_21_io_uop_is_jalr
                                              : _GEN_248
                                                  ? _slots_20_io_uop_is_jalr
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_is_jalr
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_is_jalr
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_is_jalr
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_is_jalr
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_is_jalr
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_is_jalr
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_is_jalr
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_is_jalr
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_is_jalr
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_is_jalr
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_is_jalr
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_is_jalr
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_is_jalr
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_is_jalr
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_is_jalr
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_is_jalr
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_is_jalr
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_is_jalr
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_is_jalr
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_is_jalr;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_is_jal =
    _GEN_344
      ? _slots_31_io_uop_is_jal
      : _GEN_338
          ? _slots_30_io_uop_is_jal
          : _GEN_329
              ? _slots_29_io_uop_is_jal
              : _GEN_320
                  ? _slots_28_io_uop_is_jal
                  : _GEN_311
                      ? _slots_27_io_uop_is_jal
                      : _GEN_302
                          ? _slots_26_io_uop_is_jal
                          : _GEN_293
                              ? _slots_25_io_uop_is_jal
                              : _GEN_284
                                  ? _slots_24_io_uop_is_jal
                                  : _GEN_275
                                      ? _slots_23_io_uop_is_jal
                                      : _GEN_266
                                          ? _slots_22_io_uop_is_jal
                                          : _GEN_257
                                              ? _slots_21_io_uop_is_jal
                                              : _GEN_248
                                                  ? _slots_20_io_uop_is_jal
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_is_jal
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_is_jal
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_is_jal
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_is_jal
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_is_jal
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_is_jal
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_is_jal
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_is_jal
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_is_jal
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_is_jal
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_is_jal
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_is_jal
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_is_jal
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_is_jal
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_is_jal
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_is_jal
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_is_jal
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_is_jal
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_is_jal
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_is_jal;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_is_sfb =
    _GEN_344
      ? _slots_31_io_uop_is_sfb
      : _GEN_338
          ? _slots_30_io_uop_is_sfb
          : _GEN_329
              ? _slots_29_io_uop_is_sfb
              : _GEN_320
                  ? _slots_28_io_uop_is_sfb
                  : _GEN_311
                      ? _slots_27_io_uop_is_sfb
                      : _GEN_302
                          ? _slots_26_io_uop_is_sfb
                          : _GEN_293
                              ? _slots_25_io_uop_is_sfb
                              : _GEN_284
                                  ? _slots_24_io_uop_is_sfb
                                  : _GEN_275
                                      ? _slots_23_io_uop_is_sfb
                                      : _GEN_266
                                          ? _slots_22_io_uop_is_sfb
                                          : _GEN_257
                                              ? _slots_21_io_uop_is_sfb
                                              : _GEN_248
                                                  ? _slots_20_io_uop_is_sfb
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_is_sfb
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_is_sfb
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_is_sfb
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_is_sfb
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_is_sfb
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_is_sfb
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_is_sfb
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_is_sfb
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_is_sfb
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_is_sfb
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_is_sfb
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_is_sfb
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_is_sfb
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_is_sfb
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_is_sfb
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_is_sfb
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_is_sfb
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_is_sfb
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_is_sfb
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_is_sfb;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_br_mask =
    _GEN_344
      ? _slots_31_io_uop_br_mask
      : _GEN_338
          ? _slots_30_io_uop_br_mask
          : _GEN_329
              ? _slots_29_io_uop_br_mask
              : _GEN_320
                  ? _slots_28_io_uop_br_mask
                  : _GEN_311
                      ? _slots_27_io_uop_br_mask
                      : _GEN_302
                          ? _slots_26_io_uop_br_mask
                          : _GEN_293
                              ? _slots_25_io_uop_br_mask
                              : _GEN_284
                                  ? _slots_24_io_uop_br_mask
                                  : _GEN_275
                                      ? _slots_23_io_uop_br_mask
                                      : _GEN_266
                                          ? _slots_22_io_uop_br_mask
                                          : _GEN_257
                                              ? _slots_21_io_uop_br_mask
                                              : _GEN_248
                                                  ? _slots_20_io_uop_br_mask
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_br_mask
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_br_mask
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_br_mask
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_br_mask
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_br_mask
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_br_mask
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_br_mask
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_br_mask
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_br_mask
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_br_mask
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_br_mask
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_br_mask
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_br_mask
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_br_mask
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_br_mask
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_br_mask
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_br_mask
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_br_mask
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_br_mask
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_br_mask
                                                                                                                                  : 16'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_br_tag =
    _GEN_344
      ? _slots_31_io_uop_br_tag
      : _GEN_338
          ? _slots_30_io_uop_br_tag
          : _GEN_329
              ? _slots_29_io_uop_br_tag
              : _GEN_320
                  ? _slots_28_io_uop_br_tag
                  : _GEN_311
                      ? _slots_27_io_uop_br_tag
                      : _GEN_302
                          ? _slots_26_io_uop_br_tag
                          : _GEN_293
                              ? _slots_25_io_uop_br_tag
                              : _GEN_284
                                  ? _slots_24_io_uop_br_tag
                                  : _GEN_275
                                      ? _slots_23_io_uop_br_tag
                                      : _GEN_266
                                          ? _slots_22_io_uop_br_tag
                                          : _GEN_257
                                              ? _slots_21_io_uop_br_tag
                                              : _GEN_248
                                                  ? _slots_20_io_uop_br_tag
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_br_tag
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_br_tag
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_br_tag
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_br_tag
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_br_tag
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_br_tag
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_br_tag
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_br_tag
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_br_tag
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_br_tag
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_br_tag
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_br_tag
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_br_tag
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_br_tag
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_br_tag
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_br_tag
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_br_tag
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_br_tag
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_br_tag
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_br_tag
                                                                                                                                  : 4'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_ftq_idx =
    _GEN_344
      ? _slots_31_io_uop_ftq_idx
      : _GEN_338
          ? _slots_30_io_uop_ftq_idx
          : _GEN_329
              ? _slots_29_io_uop_ftq_idx
              : _GEN_320
                  ? _slots_28_io_uop_ftq_idx
                  : _GEN_311
                      ? _slots_27_io_uop_ftq_idx
                      : _GEN_302
                          ? _slots_26_io_uop_ftq_idx
                          : _GEN_293
                              ? _slots_25_io_uop_ftq_idx
                              : _GEN_284
                                  ? _slots_24_io_uop_ftq_idx
                                  : _GEN_275
                                      ? _slots_23_io_uop_ftq_idx
                                      : _GEN_266
                                          ? _slots_22_io_uop_ftq_idx
                                          : _GEN_257
                                              ? _slots_21_io_uop_ftq_idx
                                              : _GEN_248
                                                  ? _slots_20_io_uop_ftq_idx
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_ftq_idx
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_ftq_idx
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_ftq_idx
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_ftq_idx
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_ftq_idx
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_ftq_idx
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_ftq_idx
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_ftq_idx
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_ftq_idx
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_ftq_idx
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_ftq_idx
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_ftq_idx
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_ftq_idx
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_ftq_idx
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_ftq_idx
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_ftq_idx
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_ftq_idx
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_ftq_idx
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_ftq_idx
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_ftq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_0_edge_inst =
    _GEN_344
      ? _slots_31_io_uop_edge_inst
      : _GEN_338
          ? _slots_30_io_uop_edge_inst
          : _GEN_329
              ? _slots_29_io_uop_edge_inst
              : _GEN_320
                  ? _slots_28_io_uop_edge_inst
                  : _GEN_311
                      ? _slots_27_io_uop_edge_inst
                      : _GEN_302
                          ? _slots_26_io_uop_edge_inst
                          : _GEN_293
                              ? _slots_25_io_uop_edge_inst
                              : _GEN_284
                                  ? _slots_24_io_uop_edge_inst
                                  : _GEN_275
                                      ? _slots_23_io_uop_edge_inst
                                      : _GEN_266
                                          ? _slots_22_io_uop_edge_inst
                                          : _GEN_257
                                              ? _slots_21_io_uop_edge_inst
                                              : _GEN_248
                                                  ? _slots_20_io_uop_edge_inst
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_edge_inst
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_edge_inst
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_edge_inst
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_edge_inst
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_edge_inst
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_edge_inst
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_edge_inst
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_edge_inst
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_edge_inst
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_edge_inst
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_edge_inst
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_edge_inst
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_edge_inst
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_edge_inst
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_edge_inst
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_edge_inst
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_edge_inst
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_edge_inst
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_edge_inst
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_edge_inst;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_pc_lob =
    _GEN_344
      ? _slots_31_io_uop_pc_lob
      : _GEN_338
          ? _slots_30_io_uop_pc_lob
          : _GEN_329
              ? _slots_29_io_uop_pc_lob
              : _GEN_320
                  ? _slots_28_io_uop_pc_lob
                  : _GEN_311
                      ? _slots_27_io_uop_pc_lob
                      : _GEN_302
                          ? _slots_26_io_uop_pc_lob
                          : _GEN_293
                              ? _slots_25_io_uop_pc_lob
                              : _GEN_284
                                  ? _slots_24_io_uop_pc_lob
                                  : _GEN_275
                                      ? _slots_23_io_uop_pc_lob
                                      : _GEN_266
                                          ? _slots_22_io_uop_pc_lob
                                          : _GEN_257
                                              ? _slots_21_io_uop_pc_lob
                                              : _GEN_248
                                                  ? _slots_20_io_uop_pc_lob
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_pc_lob
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_pc_lob
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_pc_lob
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_pc_lob
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_pc_lob
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_pc_lob
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_pc_lob
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_pc_lob
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_pc_lob
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_pc_lob
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_pc_lob
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_pc_lob
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_pc_lob
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_pc_lob
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_pc_lob
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_pc_lob
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_pc_lob
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_pc_lob
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_pc_lob
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_pc_lob
                                                                                                                                  : 6'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_taken =
    _GEN_344
      ? _slots_31_io_uop_taken
      : _GEN_338
          ? _slots_30_io_uop_taken
          : _GEN_329
              ? _slots_29_io_uop_taken
              : _GEN_320
                  ? _slots_28_io_uop_taken
                  : _GEN_311
                      ? _slots_27_io_uop_taken
                      : _GEN_302
                          ? _slots_26_io_uop_taken
                          : _GEN_293
                              ? _slots_25_io_uop_taken
                              : _GEN_284
                                  ? _slots_24_io_uop_taken
                                  : _GEN_275
                                      ? _slots_23_io_uop_taken
                                      : _GEN_266
                                          ? _slots_22_io_uop_taken
                                          : _GEN_257
                                              ? _slots_21_io_uop_taken
                                              : _GEN_248
                                                  ? _slots_20_io_uop_taken
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_taken
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_taken
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_taken
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_taken
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_taken
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_taken
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_taken
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_taken
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_taken
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_taken
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_taken
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_taken
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_taken
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_taken
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_taken
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_taken
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_taken
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_taken
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_taken
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_taken;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_imm_packed =
    _GEN_344
      ? _slots_31_io_uop_imm_packed
      : _GEN_338
          ? _slots_30_io_uop_imm_packed
          : _GEN_329
              ? _slots_29_io_uop_imm_packed
              : _GEN_320
                  ? _slots_28_io_uop_imm_packed
                  : _GEN_311
                      ? _slots_27_io_uop_imm_packed
                      : _GEN_302
                          ? _slots_26_io_uop_imm_packed
                          : _GEN_293
                              ? _slots_25_io_uop_imm_packed
                              : _GEN_284
                                  ? _slots_24_io_uop_imm_packed
                                  : _GEN_275
                                      ? _slots_23_io_uop_imm_packed
                                      : _GEN_266
                                          ? _slots_22_io_uop_imm_packed
                                          : _GEN_257
                                              ? _slots_21_io_uop_imm_packed
                                              : _GEN_248
                                                  ? _slots_20_io_uop_imm_packed
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_imm_packed
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_imm_packed
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_imm_packed
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_imm_packed
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_imm_packed
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_imm_packed
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_imm_packed
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_imm_packed
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_imm_packed
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_imm_packed
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_imm_packed
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_imm_packed
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_imm_packed
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_imm_packed
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_imm_packed
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_imm_packed
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_imm_packed
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_imm_packed
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_imm_packed
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_imm_packed
                                                                                                                                  : 20'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_rob_idx =
    _GEN_344
      ? _slots_31_io_uop_rob_idx
      : _GEN_338
          ? _slots_30_io_uop_rob_idx
          : _GEN_329
              ? _slots_29_io_uop_rob_idx
              : _GEN_320
                  ? _slots_28_io_uop_rob_idx
                  : _GEN_311
                      ? _slots_27_io_uop_rob_idx
                      : _GEN_302
                          ? _slots_26_io_uop_rob_idx
                          : _GEN_293
                              ? _slots_25_io_uop_rob_idx
                              : _GEN_284
                                  ? _slots_24_io_uop_rob_idx
                                  : _GEN_275
                                      ? _slots_23_io_uop_rob_idx
                                      : _GEN_266
                                          ? _slots_22_io_uop_rob_idx
                                          : _GEN_257
                                              ? _slots_21_io_uop_rob_idx
                                              : _GEN_248
                                                  ? _slots_20_io_uop_rob_idx
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_rob_idx
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_rob_idx
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_rob_idx
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_rob_idx
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_rob_idx
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_rob_idx
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_rob_idx
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_rob_idx
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_rob_idx
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_rob_idx
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_rob_idx
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_rob_idx
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_rob_idx
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_rob_idx
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_rob_idx
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_rob_idx
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_rob_idx
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_rob_idx
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_rob_idx
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_rob_idx
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_ldq_idx =
    _GEN_344
      ? _slots_31_io_uop_ldq_idx
      : _GEN_338
          ? _slots_30_io_uop_ldq_idx
          : _GEN_329
              ? _slots_29_io_uop_ldq_idx
              : _GEN_320
                  ? _slots_28_io_uop_ldq_idx
                  : _GEN_311
                      ? _slots_27_io_uop_ldq_idx
                      : _GEN_302
                          ? _slots_26_io_uop_ldq_idx
                          : _GEN_293
                              ? _slots_25_io_uop_ldq_idx
                              : _GEN_284
                                  ? _slots_24_io_uop_ldq_idx
                                  : _GEN_275
                                      ? _slots_23_io_uop_ldq_idx
                                      : _GEN_266
                                          ? _slots_22_io_uop_ldq_idx
                                          : _GEN_257
                                              ? _slots_21_io_uop_ldq_idx
                                              : _GEN_248
                                                  ? _slots_20_io_uop_ldq_idx
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_ldq_idx
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_ldq_idx
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_ldq_idx
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_ldq_idx
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_ldq_idx
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_ldq_idx
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_ldq_idx
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_ldq_idx
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_ldq_idx
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_ldq_idx
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_ldq_idx
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_ldq_idx
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_ldq_idx
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_ldq_idx
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_ldq_idx
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_ldq_idx
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_ldq_idx
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_ldq_idx
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_ldq_idx
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_ldq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_0_stq_idx =
    _GEN_344
      ? _slots_31_io_uop_stq_idx
      : _GEN_338
          ? _slots_30_io_uop_stq_idx
          : _GEN_329
              ? _slots_29_io_uop_stq_idx
              : _GEN_320
                  ? _slots_28_io_uop_stq_idx
                  : _GEN_311
                      ? _slots_27_io_uop_stq_idx
                      : _GEN_302
                          ? _slots_26_io_uop_stq_idx
                          : _GEN_293
                              ? _slots_25_io_uop_stq_idx
                              : _GEN_284
                                  ? _slots_24_io_uop_stq_idx
                                  : _GEN_275
                                      ? _slots_23_io_uop_stq_idx
                                      : _GEN_266
                                          ? _slots_22_io_uop_stq_idx
                                          : _GEN_257
                                              ? _slots_21_io_uop_stq_idx
                                              : _GEN_248
                                                  ? _slots_20_io_uop_stq_idx
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_stq_idx
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_stq_idx
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_stq_idx
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_stq_idx
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_stq_idx
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_stq_idx
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_stq_idx
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_stq_idx
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_stq_idx
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_stq_idx
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_stq_idx
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_stq_idx
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_stq_idx
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_stq_idx
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_stq_idx
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_stq_idx
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_stq_idx
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_stq_idx
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_stq_idx
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_stq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_0_pdst =
    _GEN_344
      ? _slots_31_io_uop_pdst
      : _GEN_338
          ? _slots_30_io_uop_pdst
          : _GEN_329
              ? _slots_29_io_uop_pdst
              : _GEN_320
                  ? _slots_28_io_uop_pdst
                  : _GEN_311
                      ? _slots_27_io_uop_pdst
                      : _GEN_302
                          ? _slots_26_io_uop_pdst
                          : _GEN_293
                              ? _slots_25_io_uop_pdst
                              : _GEN_284
                                  ? _slots_24_io_uop_pdst
                                  : _GEN_275
                                      ? _slots_23_io_uop_pdst
                                      : _GEN_266
                                          ? _slots_22_io_uop_pdst
                                          : _GEN_257
                                              ? _slots_21_io_uop_pdst
                                              : _GEN_248
                                                  ? _slots_20_io_uop_pdst
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_pdst
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_pdst
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_pdst
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_pdst
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_pdst
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_pdst
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_pdst
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_pdst
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_pdst
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_pdst
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_pdst
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_pdst
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_pdst
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_pdst
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_pdst
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_pdst
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_pdst
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_pdst
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_pdst
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_pdst
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_prs1 =
    _GEN_344
      ? _slots_31_io_uop_prs1
      : _GEN_338
          ? _slots_30_io_uop_prs1
          : _GEN_329
              ? _slots_29_io_uop_prs1
              : _GEN_320
                  ? _slots_28_io_uop_prs1
                  : _GEN_311
                      ? _slots_27_io_uop_prs1
                      : _GEN_302
                          ? _slots_26_io_uop_prs1
                          : _GEN_293
                              ? _slots_25_io_uop_prs1
                              : _GEN_284
                                  ? _slots_24_io_uop_prs1
                                  : _GEN_275
                                      ? _slots_23_io_uop_prs1
                                      : _GEN_266
                                          ? _slots_22_io_uop_prs1
                                          : _GEN_257
                                              ? _slots_21_io_uop_prs1
                                              : _GEN_248
                                                  ? _slots_20_io_uop_prs1
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_prs1
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_prs1
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_prs1
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_prs1
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_prs1
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_prs1
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_prs1
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_prs1
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_prs1
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_prs1
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_prs1
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_prs1
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_prs1
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_prs1
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_prs1
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_prs1
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_prs1
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_prs1
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_prs1
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_prs1
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:98:25, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_prs2 =
    _GEN_344
      ? _slots_31_io_uop_prs2
      : _GEN_338
          ? _slots_30_io_uop_prs2
          : _GEN_329
              ? _slots_29_io_uop_prs2
              : _GEN_320
                  ? _slots_28_io_uop_prs2
                  : _GEN_311
                      ? _slots_27_io_uop_prs2
                      : _GEN_302
                          ? _slots_26_io_uop_prs2
                          : _GEN_293
                              ? _slots_25_io_uop_prs2
                              : _GEN_284
                                  ? _slots_24_io_uop_prs2
                                  : _GEN_275
                                      ? _slots_23_io_uop_prs2
                                      : _GEN_266
                                          ? _slots_22_io_uop_prs2
                                          : _GEN_257
                                              ? _slots_21_io_uop_prs2
                                              : _GEN_248
                                                  ? _slots_20_io_uop_prs2
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_prs2
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_prs2
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_prs2
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_prs2
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_prs2
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_prs2
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_prs2
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_prs2
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_prs2
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_prs2
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_prs2
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_prs2
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_prs2
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_prs2
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_prs2
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_prs2
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_prs2
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_prs2
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_prs2
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_prs2
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:99:25, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_bypassable =
    _GEN_344
      ? _slots_31_io_uop_bypassable
      : _GEN_338
          ? _slots_30_io_uop_bypassable
          : _GEN_329
              ? _slots_29_io_uop_bypassable
              : _GEN_320
                  ? _slots_28_io_uop_bypassable
                  : _GEN_311
                      ? _slots_27_io_uop_bypassable
                      : _GEN_302
                          ? _slots_26_io_uop_bypassable
                          : _GEN_293
                              ? _slots_25_io_uop_bypassable
                              : _GEN_284
                                  ? _slots_24_io_uop_bypassable
                                  : _GEN_275
                                      ? _slots_23_io_uop_bypassable
                                      : _GEN_266
                                          ? _slots_22_io_uop_bypassable
                                          : _GEN_257
                                              ? _slots_21_io_uop_bypassable
                                              : _GEN_248
                                                  ? _slots_20_io_uop_bypassable
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_bypassable
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_bypassable
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_bypassable
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_bypassable
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_bypassable
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_bypassable
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_bypassable
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_bypassable
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_bypassable
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_bypassable
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_bypassable
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_bypassable
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_bypassable
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_bypassable
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_bypassable
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_bypassable
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_bypassable
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_bypassable
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_bypassable
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_bypassable;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_mem_cmd =
    _GEN_344
      ? _slots_31_io_uop_mem_cmd
      : _GEN_338
          ? _slots_30_io_uop_mem_cmd
          : _GEN_329
              ? _slots_29_io_uop_mem_cmd
              : _GEN_320
                  ? _slots_28_io_uop_mem_cmd
                  : _GEN_311
                      ? _slots_27_io_uop_mem_cmd
                      : _GEN_302
                          ? _slots_26_io_uop_mem_cmd
                          : _GEN_293
                              ? _slots_25_io_uop_mem_cmd
                              : _GEN_284
                                  ? _slots_24_io_uop_mem_cmd
                                  : _GEN_275
                                      ? _slots_23_io_uop_mem_cmd
                                      : _GEN_266
                                          ? _slots_22_io_uop_mem_cmd
                                          : _GEN_257
                                              ? _slots_21_io_uop_mem_cmd
                                              : _GEN_248
                                                  ? _slots_20_io_uop_mem_cmd
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_mem_cmd
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_mem_cmd
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_mem_cmd
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_mem_cmd
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_mem_cmd
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_mem_cmd
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_mem_cmd
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_mem_cmd
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_mem_cmd
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_mem_cmd
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_mem_cmd
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_mem_cmd
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_mem_cmd
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_mem_cmd
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_mem_cmd
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_mem_cmd
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_mem_cmd
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_mem_cmd
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_mem_cmd
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_mem_cmd
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_0_is_amo =
    _GEN_344
      ? _slots_31_io_uop_is_amo
      : _GEN_338
          ? _slots_30_io_uop_is_amo
          : _GEN_329
              ? _slots_29_io_uop_is_amo
              : _GEN_320
                  ? _slots_28_io_uop_is_amo
                  : _GEN_311
                      ? _slots_27_io_uop_is_amo
                      : _GEN_302
                          ? _slots_26_io_uop_is_amo
                          : _GEN_293
                              ? _slots_25_io_uop_is_amo
                              : _GEN_284
                                  ? _slots_24_io_uop_is_amo
                                  : _GEN_275
                                      ? _slots_23_io_uop_is_amo
                                      : _GEN_266
                                          ? _slots_22_io_uop_is_amo
                                          : _GEN_257
                                              ? _slots_21_io_uop_is_amo
                                              : _GEN_248
                                                  ? _slots_20_io_uop_is_amo
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_is_amo
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_is_amo
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_is_amo
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_is_amo
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_is_amo
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_is_amo
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_is_amo
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_is_amo
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_is_amo
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_is_amo
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_is_amo
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_is_amo
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_is_amo
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_is_amo
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_is_amo
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_is_amo
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_is_amo
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_is_amo
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_is_amo
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_is_amo;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_uses_stq =
    _GEN_344
      ? _slots_31_io_uop_uses_stq
      : _GEN_338
          ? _slots_30_io_uop_uses_stq
          : _GEN_329
              ? _slots_29_io_uop_uses_stq
              : _GEN_320
                  ? _slots_28_io_uop_uses_stq
                  : _GEN_311
                      ? _slots_27_io_uop_uses_stq
                      : _GEN_302
                          ? _slots_26_io_uop_uses_stq
                          : _GEN_293
                              ? _slots_25_io_uop_uses_stq
                              : _GEN_284
                                  ? _slots_24_io_uop_uses_stq
                                  : _GEN_275
                                      ? _slots_23_io_uop_uses_stq
                                      : _GEN_266
                                          ? _slots_22_io_uop_uses_stq
                                          : _GEN_257
                                              ? _slots_21_io_uop_uses_stq
                                              : _GEN_248
                                                  ? _slots_20_io_uop_uses_stq
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_uses_stq
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_uses_stq
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_uses_stq
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_uses_stq
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_uses_stq
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_uses_stq
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_uses_stq
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_uses_stq
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_uses_stq
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_uses_stq
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_uses_stq
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_uses_stq
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_uses_stq
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_uses_stq
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_uses_stq
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_uses_stq
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_uses_stq
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_uses_stq
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_uses_stq
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_uses_stq;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_ldst_val =
    _GEN_344
      ? _slots_31_io_uop_ldst_val
      : _GEN_338
          ? _slots_30_io_uop_ldst_val
          : _GEN_329
              ? _slots_29_io_uop_ldst_val
              : _GEN_320
                  ? _slots_28_io_uop_ldst_val
                  : _GEN_311
                      ? _slots_27_io_uop_ldst_val
                      : _GEN_302
                          ? _slots_26_io_uop_ldst_val
                          : _GEN_293
                              ? _slots_25_io_uop_ldst_val
                              : _GEN_284
                                  ? _slots_24_io_uop_ldst_val
                                  : _GEN_275
                                      ? _slots_23_io_uop_ldst_val
                                      : _GEN_266
                                          ? _slots_22_io_uop_ldst_val
                                          : _GEN_257
                                              ? _slots_21_io_uop_ldst_val
                                              : _GEN_248
                                                  ? _slots_20_io_uop_ldst_val
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_ldst_val
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_ldst_val
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_ldst_val
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_ldst_val
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_ldst_val
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_ldst_val
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_ldst_val
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_ldst_val
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_ldst_val
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_ldst_val
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_ldst_val
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_ldst_val
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_ldst_val
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_ldst_val
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_ldst_val
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_ldst_val
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_ldst_val
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_ldst_val
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_ldst_val
                                                                                                                              : _GEN_73
                                                                                                                                & _slots_0_io_uop_ldst_val;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_0_dst_rtype =
    _GEN_344
      ? _slots_31_io_uop_dst_rtype
      : _GEN_338
          ? _slots_30_io_uop_dst_rtype
          : _GEN_329
              ? _slots_29_io_uop_dst_rtype
              : _GEN_320
                  ? _slots_28_io_uop_dst_rtype
                  : _GEN_311
                      ? _slots_27_io_uop_dst_rtype
                      : _GEN_302
                          ? _slots_26_io_uop_dst_rtype
                          : _GEN_293
                              ? _slots_25_io_uop_dst_rtype
                              : _GEN_284
                                  ? _slots_24_io_uop_dst_rtype
                                  : _GEN_275
                                      ? _slots_23_io_uop_dst_rtype
                                      : _GEN_266
                                          ? _slots_22_io_uop_dst_rtype
                                          : _GEN_257
                                              ? _slots_21_io_uop_dst_rtype
                                              : _GEN_248
                                                  ? _slots_20_io_uop_dst_rtype
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_dst_rtype
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_dst_rtype
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_dst_rtype
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_dst_rtype
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_dst_rtype
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_dst_rtype
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_dst_rtype
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_dst_rtype
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_dst_rtype
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_dst_rtype
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_dst_rtype
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_dst_rtype
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_dst_rtype
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_dst_rtype
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_dst_rtype
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_dst_rtype
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_dst_rtype
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_dst_rtype
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_dst_rtype
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_dst_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_0_lrs1_rtype =
    _GEN_344
      ? _slots_31_io_uop_lrs1_rtype
      : _GEN_338
          ? _slots_30_io_uop_lrs1_rtype
          : _GEN_329
              ? _slots_29_io_uop_lrs1_rtype
              : _GEN_320
                  ? _slots_28_io_uop_lrs1_rtype
                  : _GEN_311
                      ? _slots_27_io_uop_lrs1_rtype
                      : _GEN_302
                          ? _slots_26_io_uop_lrs1_rtype
                          : _GEN_293
                              ? _slots_25_io_uop_lrs1_rtype
                              : _GEN_284
                                  ? _slots_24_io_uop_lrs1_rtype
                                  : _GEN_275
                                      ? _slots_23_io_uop_lrs1_rtype
                                      : _GEN_266
                                          ? _slots_22_io_uop_lrs1_rtype
                                          : _GEN_257
                                              ? _slots_21_io_uop_lrs1_rtype
                                              : _GEN_248
                                                  ? _slots_20_io_uop_lrs1_rtype
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_lrs1_rtype
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_lrs1_rtype
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_lrs1_rtype
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_lrs1_rtype
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_lrs1_rtype
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_lrs1_rtype
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_lrs1_rtype
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_lrs1_rtype
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_lrs1_rtype
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_lrs1_rtype
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_lrs1_rtype
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_lrs1_rtype
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_lrs1_rtype
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_lrs1_rtype
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_lrs1_rtype
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_lrs1_rtype
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_lrs1_rtype
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_lrs1_rtype
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_lrs1_rtype
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_lrs1_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:101:31, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_0_lrs2_rtype =
    _GEN_344
      ? _slots_31_io_uop_lrs2_rtype
      : _GEN_338
          ? _slots_30_io_uop_lrs2_rtype
          : _GEN_329
              ? _slots_29_io_uop_lrs2_rtype
              : _GEN_320
                  ? _slots_28_io_uop_lrs2_rtype
                  : _GEN_311
                      ? _slots_27_io_uop_lrs2_rtype
                      : _GEN_302
                          ? _slots_26_io_uop_lrs2_rtype
                          : _GEN_293
                              ? _slots_25_io_uop_lrs2_rtype
                              : _GEN_284
                                  ? _slots_24_io_uop_lrs2_rtype
                                  : _GEN_275
                                      ? _slots_23_io_uop_lrs2_rtype
                                      : _GEN_266
                                          ? _slots_22_io_uop_lrs2_rtype
                                          : _GEN_257
                                              ? _slots_21_io_uop_lrs2_rtype
                                              : _GEN_248
                                                  ? _slots_20_io_uop_lrs2_rtype
                                                  : _GEN_239
                                                      ? _slots_19_io_uop_lrs2_rtype
                                                      : _GEN_230
                                                          ? _slots_18_io_uop_lrs2_rtype
                                                          : _GEN_221
                                                              ? _slots_17_io_uop_lrs2_rtype
                                                              : _GEN_212
                                                                  ? _slots_16_io_uop_lrs2_rtype
                                                                  : _GEN_203
                                                                      ? _slots_15_io_uop_lrs2_rtype
                                                                      : _GEN_194
                                                                          ? _slots_14_io_uop_lrs2_rtype
                                                                          : _GEN_185
                                                                              ? _slots_13_io_uop_lrs2_rtype
                                                                              : _GEN_176
                                                                                  ? _slots_12_io_uop_lrs2_rtype
                                                                                  : _GEN_167
                                                                                      ? _slots_11_io_uop_lrs2_rtype
                                                                                      : _GEN_158
                                                                                          ? _slots_10_io_uop_lrs2_rtype
                                                                                          : _GEN_149
                                                                                              ? _slots_9_io_uop_lrs2_rtype
                                                                                              : _GEN_140
                                                                                                  ? _slots_8_io_uop_lrs2_rtype
                                                                                                  : _GEN_131
                                                                                                      ? _slots_7_io_uop_lrs2_rtype
                                                                                                      : _GEN_122
                                                                                                          ? _slots_6_io_uop_lrs2_rtype
                                                                                                          : _GEN_113
                                                                                                              ? _slots_5_io_uop_lrs2_rtype
                                                                                                              : _GEN_104
                                                                                                                  ? _slots_4_io_uop_lrs2_rtype
                                                                                                                  : _GEN_95
                                                                                                                      ? _slots_3_io_uop_lrs2_rtype
                                                                                                                      : _GEN_86
                                                                                                                          ? _slots_2_io_uop_lrs2_rtype
                                                                                                                          : _GEN_77
                                                                                                                              ? _slots_1_io_uop_lrs2_rtype
                                                                                                                              : _GEN_73
                                                                                                                                  ? _slots_0_io_uop_lrs2_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:102:31, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_1_uopc =
    _GEN_345
      ? _slots_31_io_uop_uopc
      : _GEN_340
          ? _slots_30_io_uop_uopc
          : _GEN_332
              ? _slots_29_io_uop_uopc
              : _GEN_323
                  ? _slots_28_io_uop_uopc
                  : _GEN_314
                      ? _slots_27_io_uop_uopc
                      : _GEN_305
                          ? _slots_26_io_uop_uopc
                          : _GEN_296
                              ? _slots_25_io_uop_uopc
                              : _GEN_287
                                  ? _slots_24_io_uop_uopc
                                  : _GEN_278
                                      ? _slots_23_io_uop_uopc
                                      : _GEN_269
                                          ? _slots_22_io_uop_uopc
                                          : _GEN_260
                                              ? _slots_21_io_uop_uopc
                                              : _GEN_251
                                                  ? _slots_20_io_uop_uopc
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_uopc
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_uopc
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_uopc
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_uopc
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_uopc
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_uopc
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_uopc
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_uopc
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_uopc
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_uopc
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_uopc
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_uopc
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_uopc
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_uopc
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_uopc
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_uopc
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_uopc
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_uopc
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_uopc
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_uopc
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_inst =
    _GEN_345
      ? _slots_31_io_uop_inst
      : _GEN_340
          ? _slots_30_io_uop_inst
          : _GEN_332
              ? _slots_29_io_uop_inst
              : _GEN_323
                  ? _slots_28_io_uop_inst
                  : _GEN_314
                      ? _slots_27_io_uop_inst
                      : _GEN_305
                          ? _slots_26_io_uop_inst
                          : _GEN_296
                              ? _slots_25_io_uop_inst
                              : _GEN_287
                                  ? _slots_24_io_uop_inst
                                  : _GEN_278
                                      ? _slots_23_io_uop_inst
                                      : _GEN_269
                                          ? _slots_22_io_uop_inst
                                          : _GEN_260
                                              ? _slots_21_io_uop_inst
                                              : _GEN_251
                                                  ? _slots_20_io_uop_inst
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_inst
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_inst
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_inst
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_inst
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_inst
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_inst
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_inst
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_inst
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_inst
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_inst
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_inst
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_inst
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_inst
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_inst
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_inst
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_inst
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_inst
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_inst
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_inst
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_inst
                                                                                                                                  : 32'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_debug_inst =
    _GEN_345
      ? _slots_31_io_uop_debug_inst
      : _GEN_340
          ? _slots_30_io_uop_debug_inst
          : _GEN_332
              ? _slots_29_io_uop_debug_inst
              : _GEN_323
                  ? _slots_28_io_uop_debug_inst
                  : _GEN_314
                      ? _slots_27_io_uop_debug_inst
                      : _GEN_305
                          ? _slots_26_io_uop_debug_inst
                          : _GEN_296
                              ? _slots_25_io_uop_debug_inst
                              : _GEN_287
                                  ? _slots_24_io_uop_debug_inst
                                  : _GEN_278
                                      ? _slots_23_io_uop_debug_inst
                                      : _GEN_269
                                          ? _slots_22_io_uop_debug_inst
                                          : _GEN_260
                                              ? _slots_21_io_uop_debug_inst
                                              : _GEN_251
                                                  ? _slots_20_io_uop_debug_inst
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_debug_inst
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_debug_inst
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_debug_inst
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_debug_inst
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_debug_inst
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_debug_inst
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_debug_inst
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_debug_inst
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_debug_inst
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_debug_inst
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_debug_inst
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_debug_inst
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_debug_inst
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_debug_inst
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_debug_inst
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_debug_inst
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_debug_inst
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_debug_inst
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_debug_inst
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_debug_inst
                                                                                                                                  : 32'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_rvc =
    _GEN_345
      ? _slots_31_io_uop_is_rvc
      : _GEN_340
          ? _slots_30_io_uop_is_rvc
          : _GEN_332
              ? _slots_29_io_uop_is_rvc
              : _GEN_323
                  ? _slots_28_io_uop_is_rvc
                  : _GEN_314
                      ? _slots_27_io_uop_is_rvc
                      : _GEN_305
                          ? _slots_26_io_uop_is_rvc
                          : _GEN_296
                              ? _slots_25_io_uop_is_rvc
                              : _GEN_287
                                  ? _slots_24_io_uop_is_rvc
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_rvc
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_rvc
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_rvc
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_rvc
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_rvc
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_rvc
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_rvc
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_rvc
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_rvc
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_rvc
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_rvc
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_rvc
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_rvc
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_rvc
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_rvc
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_rvc
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_rvc
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_rvc
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_rvc
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_rvc
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_rvc
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_rvc
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_rvc
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_rvc;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_debug_pc =
    _GEN_345
      ? _slots_31_io_uop_debug_pc
      : _GEN_340
          ? _slots_30_io_uop_debug_pc
          : _GEN_332
              ? _slots_29_io_uop_debug_pc
              : _GEN_323
                  ? _slots_28_io_uop_debug_pc
                  : _GEN_314
                      ? _slots_27_io_uop_debug_pc
                      : _GEN_305
                          ? _slots_26_io_uop_debug_pc
                          : _GEN_296
                              ? _slots_25_io_uop_debug_pc
                              : _GEN_287
                                  ? _slots_24_io_uop_debug_pc
                                  : _GEN_278
                                      ? _slots_23_io_uop_debug_pc
                                      : _GEN_269
                                          ? _slots_22_io_uop_debug_pc
                                          : _GEN_260
                                              ? _slots_21_io_uop_debug_pc
                                              : _GEN_251
                                                  ? _slots_20_io_uop_debug_pc
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_debug_pc
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_debug_pc
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_debug_pc
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_debug_pc
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_debug_pc
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_debug_pc
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_debug_pc
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_debug_pc
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_debug_pc
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_debug_pc
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_debug_pc
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_debug_pc
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_debug_pc
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_debug_pc
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_debug_pc
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_debug_pc
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_debug_pc
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_debug_pc
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_debug_pc
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_debug_pc
                                                                                                                                  : 40'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_iq_type =
    _GEN_345
      ? _slots_31_io_uop_iq_type
      : _GEN_340
          ? _slots_30_io_uop_iq_type
          : _GEN_332
              ? _slots_29_io_uop_iq_type
              : _GEN_323
                  ? _slots_28_io_uop_iq_type
                  : _GEN_314
                      ? _slots_27_io_uop_iq_type
                      : _GEN_305
                          ? _slots_26_io_uop_iq_type
                          : _GEN_296
                              ? _slots_25_io_uop_iq_type
                              : _GEN_287
                                  ? _slots_24_io_uop_iq_type
                                  : _GEN_278
                                      ? _slots_23_io_uop_iq_type
                                      : _GEN_269
                                          ? _slots_22_io_uop_iq_type
                                          : _GEN_260
                                              ? _slots_21_io_uop_iq_type
                                              : _GEN_251
                                                  ? _slots_20_io_uop_iq_type
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_iq_type
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_iq_type
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_iq_type
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_iq_type
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_iq_type
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_iq_type
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_iq_type
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_iq_type
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_iq_type
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_iq_type
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_iq_type
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_iq_type
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_iq_type
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_iq_type
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_iq_type
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_iq_type
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_iq_type
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_iq_type
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_iq_type
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_iq_type
                                                                                                                                  : 3'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_fu_code =
    _GEN_345
      ? _slots_31_io_uop_fu_code
      : _GEN_340
          ? _slots_30_io_uop_fu_code
          : _GEN_332
              ? _slots_29_io_uop_fu_code
              : _GEN_323
                  ? _slots_28_io_uop_fu_code
                  : _GEN_314
                      ? _slots_27_io_uop_fu_code
                      : _GEN_305
                          ? _slots_26_io_uop_fu_code
                          : _GEN_296
                              ? _slots_25_io_uop_fu_code
                              : _GEN_287
                                  ? _slots_24_io_uop_fu_code
                                  : _GEN_278
                                      ? _slots_23_io_uop_fu_code
                                      : _GEN_269
                                          ? _slots_22_io_uop_fu_code
                                          : _GEN_260
                                              ? _slots_21_io_uop_fu_code
                                              : _GEN_251
                                                  ? _slots_20_io_uop_fu_code
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_fu_code
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_fu_code
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_fu_code
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_fu_code
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_fu_code
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_fu_code
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_fu_code
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_fu_code
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_fu_code
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_fu_code
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_fu_code
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_fu_code
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_fu_code
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_fu_code
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_fu_code
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_fu_code
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_fu_code
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_fu_code
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_fu_code
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_fu_code
                                                                                                                                  : 10'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_iw_state =
    _GEN_345
      ? _slots_31_io_uop_iw_state
      : _GEN_340
          ? _slots_30_io_uop_iw_state
          : _GEN_332
              ? _slots_29_io_uop_iw_state
              : _GEN_323
                  ? _slots_28_io_uop_iw_state
                  : _GEN_314
                      ? _slots_27_io_uop_iw_state
                      : _GEN_305
                          ? _slots_26_io_uop_iw_state
                          : _GEN_296
                              ? _slots_25_io_uop_iw_state
                              : _GEN_287
                                  ? _slots_24_io_uop_iw_state
                                  : _GEN_278
                                      ? _slots_23_io_uop_iw_state
                                      : _GEN_269
                                          ? _slots_22_io_uop_iw_state
                                          : _GEN_260
                                              ? _slots_21_io_uop_iw_state
                                              : _GEN_251
                                                  ? _slots_20_io_uop_iw_state
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_iw_state
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_iw_state
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_iw_state
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_iw_state
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_iw_state
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_iw_state
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_iw_state
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_iw_state
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_iw_state
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_iw_state
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_iw_state
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_iw_state
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_iw_state
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_iw_state
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_iw_state
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_iw_state
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_iw_state
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_iw_state
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_iw_state
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_iw_state
                                                                                                                                  : 2'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:127:84, :153:73
  assign io_iss_uops_1_iw_p1_poisoned =
    _GEN_345
      ? _slots_31_io_uop_iw_p1_poisoned
      : _GEN_340
          ? _slots_30_io_uop_iw_p1_poisoned
          : _GEN_332
              ? _slots_29_io_uop_iw_p1_poisoned
              : _GEN_323
                  ? _slots_28_io_uop_iw_p1_poisoned
                  : _GEN_314
                      ? _slots_27_io_uop_iw_p1_poisoned
                      : _GEN_305
                          ? _slots_26_io_uop_iw_p1_poisoned
                          : _GEN_296
                              ? _slots_25_io_uop_iw_p1_poisoned
                              : _GEN_287
                                  ? _slots_24_io_uop_iw_p1_poisoned
                                  : _GEN_278
                                      ? _slots_23_io_uop_iw_p1_poisoned
                                      : _GEN_269
                                          ? _slots_22_io_uop_iw_p1_poisoned
                                          : _GEN_260
                                              ? _slots_21_io_uop_iw_p1_poisoned
                                              : _GEN_251
                                                  ? _slots_20_io_uop_iw_p1_poisoned
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_iw_p1_poisoned
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_iw_p1_poisoned
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_iw_p1_poisoned
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_iw_p1_poisoned
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_iw_p1_poisoned
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_iw_p1_poisoned
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_iw_p1_poisoned
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_iw_p1_poisoned
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_iw_p1_poisoned
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_iw_p1_poisoned
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_iw_p1_poisoned
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_iw_p1_poisoned
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_iw_p1_poisoned
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_iw_p1_poisoned
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_iw_p1_poisoned
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_iw_p1_poisoned
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_iw_p1_poisoned
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_iw_p1_poisoned
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_iw_p1_poisoned
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_iw_p1_poisoned;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_iw_p2_poisoned =
    _GEN_345
      ? _slots_31_io_uop_iw_p2_poisoned
      : _GEN_340
          ? _slots_30_io_uop_iw_p2_poisoned
          : _GEN_332
              ? _slots_29_io_uop_iw_p2_poisoned
              : _GEN_323
                  ? _slots_28_io_uop_iw_p2_poisoned
                  : _GEN_314
                      ? _slots_27_io_uop_iw_p2_poisoned
                      : _GEN_305
                          ? _slots_26_io_uop_iw_p2_poisoned
                          : _GEN_296
                              ? _slots_25_io_uop_iw_p2_poisoned
                              : _GEN_287
                                  ? _slots_24_io_uop_iw_p2_poisoned
                                  : _GEN_278
                                      ? _slots_23_io_uop_iw_p2_poisoned
                                      : _GEN_269
                                          ? _slots_22_io_uop_iw_p2_poisoned
                                          : _GEN_260
                                              ? _slots_21_io_uop_iw_p2_poisoned
                                              : _GEN_251
                                                  ? _slots_20_io_uop_iw_p2_poisoned
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_iw_p2_poisoned
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_iw_p2_poisoned
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_iw_p2_poisoned
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_iw_p2_poisoned
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_iw_p2_poisoned
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_iw_p2_poisoned
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_iw_p2_poisoned
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_iw_p2_poisoned
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_iw_p2_poisoned
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_iw_p2_poisoned
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_iw_p2_poisoned
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_iw_p2_poisoned
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_iw_p2_poisoned
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_iw_p2_poisoned
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_iw_p2_poisoned
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_iw_p2_poisoned
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_iw_p2_poisoned
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_iw_p2_poisoned
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_iw_p2_poisoned
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_iw_p2_poisoned;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_br =
    _GEN_345
      ? _slots_31_io_uop_is_br
      : _GEN_340
          ? _slots_30_io_uop_is_br
          : _GEN_332
              ? _slots_29_io_uop_is_br
              : _GEN_323
                  ? _slots_28_io_uop_is_br
                  : _GEN_314
                      ? _slots_27_io_uop_is_br
                      : _GEN_305
                          ? _slots_26_io_uop_is_br
                          : _GEN_296
                              ? _slots_25_io_uop_is_br
                              : _GEN_287
                                  ? _slots_24_io_uop_is_br
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_br
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_br
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_br
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_br
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_br
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_br
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_br
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_br
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_br
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_br
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_br
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_br
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_br
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_br
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_br
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_br
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_br
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_br
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_br
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_br
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_br
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_br
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_br
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_br;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_jalr =
    _GEN_345
      ? _slots_31_io_uop_is_jalr
      : _GEN_340
          ? _slots_30_io_uop_is_jalr
          : _GEN_332
              ? _slots_29_io_uop_is_jalr
              : _GEN_323
                  ? _slots_28_io_uop_is_jalr
                  : _GEN_314
                      ? _slots_27_io_uop_is_jalr
                      : _GEN_305
                          ? _slots_26_io_uop_is_jalr
                          : _GEN_296
                              ? _slots_25_io_uop_is_jalr
                              : _GEN_287
                                  ? _slots_24_io_uop_is_jalr
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_jalr
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_jalr
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_jalr
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_jalr
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_jalr
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_jalr
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_jalr
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_jalr
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_jalr
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_jalr
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_jalr
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_jalr
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_jalr
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_jalr
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_jalr
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_jalr
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_jalr
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_jalr
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_jalr
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_jalr
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_jalr
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_jalr
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_jalr
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_jalr;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_jal =
    _GEN_345
      ? _slots_31_io_uop_is_jal
      : _GEN_340
          ? _slots_30_io_uop_is_jal
          : _GEN_332
              ? _slots_29_io_uop_is_jal
              : _GEN_323
                  ? _slots_28_io_uop_is_jal
                  : _GEN_314
                      ? _slots_27_io_uop_is_jal
                      : _GEN_305
                          ? _slots_26_io_uop_is_jal
                          : _GEN_296
                              ? _slots_25_io_uop_is_jal
                              : _GEN_287
                                  ? _slots_24_io_uop_is_jal
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_jal
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_jal
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_jal
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_jal
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_jal
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_jal
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_jal
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_jal
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_jal
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_jal
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_jal
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_jal
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_jal
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_jal
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_jal
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_jal
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_jal
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_jal
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_jal
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_jal
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_jal
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_jal
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_jal
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_jal;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_sfb =
    _GEN_345
      ? _slots_31_io_uop_is_sfb
      : _GEN_340
          ? _slots_30_io_uop_is_sfb
          : _GEN_332
              ? _slots_29_io_uop_is_sfb
              : _GEN_323
                  ? _slots_28_io_uop_is_sfb
                  : _GEN_314
                      ? _slots_27_io_uop_is_sfb
                      : _GEN_305
                          ? _slots_26_io_uop_is_sfb
                          : _GEN_296
                              ? _slots_25_io_uop_is_sfb
                              : _GEN_287
                                  ? _slots_24_io_uop_is_sfb
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_sfb
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_sfb
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_sfb
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_sfb
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_sfb
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_sfb
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_sfb
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_sfb
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_sfb
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_sfb
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_sfb
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_sfb
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_sfb
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_sfb
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_sfb
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_sfb
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_sfb
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_sfb
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_sfb
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_sfb
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_sfb
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_sfb
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_sfb
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_sfb;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_br_mask =
    _GEN_345
      ? _slots_31_io_uop_br_mask
      : _GEN_340
          ? _slots_30_io_uop_br_mask
          : _GEN_332
              ? _slots_29_io_uop_br_mask
              : _GEN_323
                  ? _slots_28_io_uop_br_mask
                  : _GEN_314
                      ? _slots_27_io_uop_br_mask
                      : _GEN_305
                          ? _slots_26_io_uop_br_mask
                          : _GEN_296
                              ? _slots_25_io_uop_br_mask
                              : _GEN_287
                                  ? _slots_24_io_uop_br_mask
                                  : _GEN_278
                                      ? _slots_23_io_uop_br_mask
                                      : _GEN_269
                                          ? _slots_22_io_uop_br_mask
                                          : _GEN_260
                                              ? _slots_21_io_uop_br_mask
                                              : _GEN_251
                                                  ? _slots_20_io_uop_br_mask
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_br_mask
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_br_mask
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_br_mask
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_br_mask
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_br_mask
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_br_mask
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_br_mask
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_br_mask
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_br_mask
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_br_mask
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_br_mask
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_br_mask
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_br_mask
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_br_mask
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_br_mask
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_br_mask
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_br_mask
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_br_mask
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_br_mask
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_br_mask
                                                                                                                                  : 16'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_br_tag =
    _GEN_345
      ? _slots_31_io_uop_br_tag
      : _GEN_340
          ? _slots_30_io_uop_br_tag
          : _GEN_332
              ? _slots_29_io_uop_br_tag
              : _GEN_323
                  ? _slots_28_io_uop_br_tag
                  : _GEN_314
                      ? _slots_27_io_uop_br_tag
                      : _GEN_305
                          ? _slots_26_io_uop_br_tag
                          : _GEN_296
                              ? _slots_25_io_uop_br_tag
                              : _GEN_287
                                  ? _slots_24_io_uop_br_tag
                                  : _GEN_278
                                      ? _slots_23_io_uop_br_tag
                                      : _GEN_269
                                          ? _slots_22_io_uop_br_tag
                                          : _GEN_260
                                              ? _slots_21_io_uop_br_tag
                                              : _GEN_251
                                                  ? _slots_20_io_uop_br_tag
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_br_tag
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_br_tag
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_br_tag
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_br_tag
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_br_tag
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_br_tag
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_br_tag
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_br_tag
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_br_tag
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_br_tag
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_br_tag
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_br_tag
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_br_tag
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_br_tag
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_br_tag
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_br_tag
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_br_tag
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_br_tag
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_br_tag
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_br_tag
                                                                                                                                  : 4'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_ftq_idx =
    _GEN_345
      ? _slots_31_io_uop_ftq_idx
      : _GEN_340
          ? _slots_30_io_uop_ftq_idx
          : _GEN_332
              ? _slots_29_io_uop_ftq_idx
              : _GEN_323
                  ? _slots_28_io_uop_ftq_idx
                  : _GEN_314
                      ? _slots_27_io_uop_ftq_idx
                      : _GEN_305
                          ? _slots_26_io_uop_ftq_idx
                          : _GEN_296
                              ? _slots_25_io_uop_ftq_idx
                              : _GEN_287
                                  ? _slots_24_io_uop_ftq_idx
                                  : _GEN_278
                                      ? _slots_23_io_uop_ftq_idx
                                      : _GEN_269
                                          ? _slots_22_io_uop_ftq_idx
                                          : _GEN_260
                                              ? _slots_21_io_uop_ftq_idx
                                              : _GEN_251
                                                  ? _slots_20_io_uop_ftq_idx
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_ftq_idx
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_ftq_idx
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_ftq_idx
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_ftq_idx
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_ftq_idx
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_ftq_idx
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_ftq_idx
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_ftq_idx
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_ftq_idx
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_ftq_idx
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_ftq_idx
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_ftq_idx
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_ftq_idx
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_ftq_idx
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_ftq_idx
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_ftq_idx
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_ftq_idx
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_ftq_idx
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_ftq_idx
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_ftq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_1_edge_inst =
    _GEN_345
      ? _slots_31_io_uop_edge_inst
      : _GEN_340
          ? _slots_30_io_uop_edge_inst
          : _GEN_332
              ? _slots_29_io_uop_edge_inst
              : _GEN_323
                  ? _slots_28_io_uop_edge_inst
                  : _GEN_314
                      ? _slots_27_io_uop_edge_inst
                      : _GEN_305
                          ? _slots_26_io_uop_edge_inst
                          : _GEN_296
                              ? _slots_25_io_uop_edge_inst
                              : _GEN_287
                                  ? _slots_24_io_uop_edge_inst
                                  : _GEN_278
                                      ? _slots_23_io_uop_edge_inst
                                      : _GEN_269
                                          ? _slots_22_io_uop_edge_inst
                                          : _GEN_260
                                              ? _slots_21_io_uop_edge_inst
                                              : _GEN_251
                                                  ? _slots_20_io_uop_edge_inst
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_edge_inst
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_edge_inst
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_edge_inst
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_edge_inst
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_edge_inst
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_edge_inst
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_edge_inst
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_edge_inst
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_edge_inst
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_edge_inst
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_edge_inst
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_edge_inst
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_edge_inst
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_edge_inst
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_edge_inst
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_edge_inst
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_edge_inst
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_edge_inst
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_edge_inst
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_edge_inst;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_pc_lob =
    _GEN_345
      ? _slots_31_io_uop_pc_lob
      : _GEN_340
          ? _slots_30_io_uop_pc_lob
          : _GEN_332
              ? _slots_29_io_uop_pc_lob
              : _GEN_323
                  ? _slots_28_io_uop_pc_lob
                  : _GEN_314
                      ? _slots_27_io_uop_pc_lob
                      : _GEN_305
                          ? _slots_26_io_uop_pc_lob
                          : _GEN_296
                              ? _slots_25_io_uop_pc_lob
                              : _GEN_287
                                  ? _slots_24_io_uop_pc_lob
                                  : _GEN_278
                                      ? _slots_23_io_uop_pc_lob
                                      : _GEN_269
                                          ? _slots_22_io_uop_pc_lob
                                          : _GEN_260
                                              ? _slots_21_io_uop_pc_lob
                                              : _GEN_251
                                                  ? _slots_20_io_uop_pc_lob
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_pc_lob
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_pc_lob
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_pc_lob
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_pc_lob
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_pc_lob
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_pc_lob
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_pc_lob
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_pc_lob
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_pc_lob
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_pc_lob
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_pc_lob
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_pc_lob
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_pc_lob
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_pc_lob
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_pc_lob
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_pc_lob
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_pc_lob
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_pc_lob
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_pc_lob
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_pc_lob
                                                                                                                                  : 6'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_taken =
    _GEN_345
      ? _slots_31_io_uop_taken
      : _GEN_340
          ? _slots_30_io_uop_taken
          : _GEN_332
              ? _slots_29_io_uop_taken
              : _GEN_323
                  ? _slots_28_io_uop_taken
                  : _GEN_314
                      ? _slots_27_io_uop_taken
                      : _GEN_305
                          ? _slots_26_io_uop_taken
                          : _GEN_296
                              ? _slots_25_io_uop_taken
                              : _GEN_287
                                  ? _slots_24_io_uop_taken
                                  : _GEN_278
                                      ? _slots_23_io_uop_taken
                                      : _GEN_269
                                          ? _slots_22_io_uop_taken
                                          : _GEN_260
                                              ? _slots_21_io_uop_taken
                                              : _GEN_251
                                                  ? _slots_20_io_uop_taken
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_taken
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_taken
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_taken
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_taken
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_taken
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_taken
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_taken
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_taken
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_taken
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_taken
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_taken
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_taken
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_taken
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_taken
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_taken
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_taken
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_taken
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_taken
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_taken
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_taken;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_imm_packed =
    _GEN_345
      ? _slots_31_io_uop_imm_packed
      : _GEN_340
          ? _slots_30_io_uop_imm_packed
          : _GEN_332
              ? _slots_29_io_uop_imm_packed
              : _GEN_323
                  ? _slots_28_io_uop_imm_packed
                  : _GEN_314
                      ? _slots_27_io_uop_imm_packed
                      : _GEN_305
                          ? _slots_26_io_uop_imm_packed
                          : _GEN_296
                              ? _slots_25_io_uop_imm_packed
                              : _GEN_287
                                  ? _slots_24_io_uop_imm_packed
                                  : _GEN_278
                                      ? _slots_23_io_uop_imm_packed
                                      : _GEN_269
                                          ? _slots_22_io_uop_imm_packed
                                          : _GEN_260
                                              ? _slots_21_io_uop_imm_packed
                                              : _GEN_251
                                                  ? _slots_20_io_uop_imm_packed
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_imm_packed
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_imm_packed
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_imm_packed
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_imm_packed
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_imm_packed
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_imm_packed
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_imm_packed
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_imm_packed
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_imm_packed
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_imm_packed
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_imm_packed
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_imm_packed
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_imm_packed
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_imm_packed
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_imm_packed
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_imm_packed
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_imm_packed
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_imm_packed
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_imm_packed
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_imm_packed
                                                                                                                                  : 20'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_csr_addr =
    _GEN_345
      ? _slots_31_io_uop_csr_addr
      : _GEN_340
          ? _slots_30_io_uop_csr_addr
          : _GEN_332
              ? _slots_29_io_uop_csr_addr
              : _GEN_323
                  ? _slots_28_io_uop_csr_addr
                  : _GEN_314
                      ? _slots_27_io_uop_csr_addr
                      : _GEN_305
                          ? _slots_26_io_uop_csr_addr
                          : _GEN_296
                              ? _slots_25_io_uop_csr_addr
                              : _GEN_287
                                  ? _slots_24_io_uop_csr_addr
                                  : _GEN_278
                                      ? _slots_23_io_uop_csr_addr
                                      : _GEN_269
                                          ? _slots_22_io_uop_csr_addr
                                          : _GEN_260
                                              ? _slots_21_io_uop_csr_addr
                                              : _GEN_251
                                                  ? _slots_20_io_uop_csr_addr
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_csr_addr
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_csr_addr
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_csr_addr
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_csr_addr
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_csr_addr
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_csr_addr
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_csr_addr
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_csr_addr
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_csr_addr
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_csr_addr
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_csr_addr
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_csr_addr
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_csr_addr
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_csr_addr
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_csr_addr
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_csr_addr
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_csr_addr
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_csr_addr
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_csr_addr
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_csr_addr
                                                                                                                                  : 12'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_rob_idx =
    _GEN_345
      ? _slots_31_io_uop_rob_idx
      : _GEN_340
          ? _slots_30_io_uop_rob_idx
          : _GEN_332
              ? _slots_29_io_uop_rob_idx
              : _GEN_323
                  ? _slots_28_io_uop_rob_idx
                  : _GEN_314
                      ? _slots_27_io_uop_rob_idx
                      : _GEN_305
                          ? _slots_26_io_uop_rob_idx
                          : _GEN_296
                              ? _slots_25_io_uop_rob_idx
                              : _GEN_287
                                  ? _slots_24_io_uop_rob_idx
                                  : _GEN_278
                                      ? _slots_23_io_uop_rob_idx
                                      : _GEN_269
                                          ? _slots_22_io_uop_rob_idx
                                          : _GEN_260
                                              ? _slots_21_io_uop_rob_idx
                                              : _GEN_251
                                                  ? _slots_20_io_uop_rob_idx
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_rob_idx
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_rob_idx
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_rob_idx
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_rob_idx
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_rob_idx
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_rob_idx
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_rob_idx
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_rob_idx
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_rob_idx
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_rob_idx
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_rob_idx
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_rob_idx
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_rob_idx
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_rob_idx
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_rob_idx
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_rob_idx
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_rob_idx
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_rob_idx
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_rob_idx
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_rob_idx
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_ldq_idx =
    _GEN_345
      ? _slots_31_io_uop_ldq_idx
      : _GEN_340
          ? _slots_30_io_uop_ldq_idx
          : _GEN_332
              ? _slots_29_io_uop_ldq_idx
              : _GEN_323
                  ? _slots_28_io_uop_ldq_idx
                  : _GEN_314
                      ? _slots_27_io_uop_ldq_idx
                      : _GEN_305
                          ? _slots_26_io_uop_ldq_idx
                          : _GEN_296
                              ? _slots_25_io_uop_ldq_idx
                              : _GEN_287
                                  ? _slots_24_io_uop_ldq_idx
                                  : _GEN_278
                                      ? _slots_23_io_uop_ldq_idx
                                      : _GEN_269
                                          ? _slots_22_io_uop_ldq_idx
                                          : _GEN_260
                                              ? _slots_21_io_uop_ldq_idx
                                              : _GEN_251
                                                  ? _slots_20_io_uop_ldq_idx
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_ldq_idx
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_ldq_idx
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_ldq_idx
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_ldq_idx
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_ldq_idx
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_ldq_idx
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_ldq_idx
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_ldq_idx
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_ldq_idx
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_ldq_idx
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_ldq_idx
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_ldq_idx
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_ldq_idx
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_ldq_idx
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_ldq_idx
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_ldq_idx
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_ldq_idx
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_ldq_idx
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_ldq_idx
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_ldq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_1_stq_idx =
    _GEN_345
      ? _slots_31_io_uop_stq_idx
      : _GEN_340
          ? _slots_30_io_uop_stq_idx
          : _GEN_332
              ? _slots_29_io_uop_stq_idx
              : _GEN_323
                  ? _slots_28_io_uop_stq_idx
                  : _GEN_314
                      ? _slots_27_io_uop_stq_idx
                      : _GEN_305
                          ? _slots_26_io_uop_stq_idx
                          : _GEN_296
                              ? _slots_25_io_uop_stq_idx
                              : _GEN_287
                                  ? _slots_24_io_uop_stq_idx
                                  : _GEN_278
                                      ? _slots_23_io_uop_stq_idx
                                      : _GEN_269
                                          ? _slots_22_io_uop_stq_idx
                                          : _GEN_260
                                              ? _slots_21_io_uop_stq_idx
                                              : _GEN_251
                                                  ? _slots_20_io_uop_stq_idx
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_stq_idx
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_stq_idx
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_stq_idx
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_stq_idx
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_stq_idx
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_stq_idx
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_stq_idx
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_stq_idx
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_stq_idx
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_stq_idx
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_stq_idx
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_stq_idx
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_stq_idx
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_stq_idx
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_stq_idx
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_stq_idx
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_stq_idx
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_stq_idx
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_stq_idx
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_stq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_1_rxq_idx =
    _GEN_345
      ? _slots_31_io_uop_rxq_idx
      : _GEN_340
          ? _slots_30_io_uop_rxq_idx
          : _GEN_332
              ? _slots_29_io_uop_rxq_idx
              : _GEN_323
                  ? _slots_28_io_uop_rxq_idx
                  : _GEN_314
                      ? _slots_27_io_uop_rxq_idx
                      : _GEN_305
                          ? _slots_26_io_uop_rxq_idx
                          : _GEN_296
                              ? _slots_25_io_uop_rxq_idx
                              : _GEN_287
                                  ? _slots_24_io_uop_rxq_idx
                                  : _GEN_278
                                      ? _slots_23_io_uop_rxq_idx
                                      : _GEN_269
                                          ? _slots_22_io_uop_rxq_idx
                                          : _GEN_260
                                              ? _slots_21_io_uop_rxq_idx
                                              : _GEN_251
                                                  ? _slots_20_io_uop_rxq_idx
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_rxq_idx
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_rxq_idx
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_rxq_idx
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_rxq_idx
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_rxq_idx
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_rxq_idx
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_rxq_idx
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_rxq_idx
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_rxq_idx
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_rxq_idx
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_rxq_idx
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_rxq_idx
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_rxq_idx
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_rxq_idx
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_rxq_idx
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_rxq_idx
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_rxq_idx
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_rxq_idx
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_rxq_idx
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_rxq_idx
                                                                                                                                  : 2'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:127:84, :153:73
  assign io_iss_uops_1_pdst =
    _GEN_345
      ? _slots_31_io_uop_pdst
      : _GEN_340
          ? _slots_30_io_uop_pdst
          : _GEN_332
              ? _slots_29_io_uop_pdst
              : _GEN_323
                  ? _slots_28_io_uop_pdst
                  : _GEN_314
                      ? _slots_27_io_uop_pdst
                      : _GEN_305
                          ? _slots_26_io_uop_pdst
                          : _GEN_296
                              ? _slots_25_io_uop_pdst
                              : _GEN_287
                                  ? _slots_24_io_uop_pdst
                                  : _GEN_278
                                      ? _slots_23_io_uop_pdst
                                      : _GEN_269
                                          ? _slots_22_io_uop_pdst
                                          : _GEN_260
                                              ? _slots_21_io_uop_pdst
                                              : _GEN_251
                                                  ? _slots_20_io_uop_pdst
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_pdst
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_pdst
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_pdst
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_pdst
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_pdst
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_pdst
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_pdst
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_pdst
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_pdst
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_pdst
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_pdst
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_pdst
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_pdst
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_pdst
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_pdst
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_pdst
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_pdst
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_pdst
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_pdst
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_pdst
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_prs1 =
    _GEN_345
      ? _slots_31_io_uop_prs1
      : _GEN_340
          ? _slots_30_io_uop_prs1
          : _GEN_332
              ? _slots_29_io_uop_prs1
              : _GEN_323
                  ? _slots_28_io_uop_prs1
                  : _GEN_314
                      ? _slots_27_io_uop_prs1
                      : _GEN_305
                          ? _slots_26_io_uop_prs1
                          : _GEN_296
                              ? _slots_25_io_uop_prs1
                              : _GEN_287
                                  ? _slots_24_io_uop_prs1
                                  : _GEN_278
                                      ? _slots_23_io_uop_prs1
                                      : _GEN_269
                                          ? _slots_22_io_uop_prs1
                                          : _GEN_260
                                              ? _slots_21_io_uop_prs1
                                              : _GEN_251
                                                  ? _slots_20_io_uop_prs1
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_prs1
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_prs1
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_prs1
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_prs1
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_prs1
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_prs1
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_prs1
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_prs1
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_prs1
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_prs1
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_prs1
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_prs1
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_prs1
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_prs1
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_prs1
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_prs1
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_prs1
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_prs1
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_prs1
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_prs1
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:98:25, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_prs2 =
    _GEN_345
      ? _slots_31_io_uop_prs2
      : _GEN_340
          ? _slots_30_io_uop_prs2
          : _GEN_332
              ? _slots_29_io_uop_prs2
              : _GEN_323
                  ? _slots_28_io_uop_prs2
                  : _GEN_314
                      ? _slots_27_io_uop_prs2
                      : _GEN_305
                          ? _slots_26_io_uop_prs2
                          : _GEN_296
                              ? _slots_25_io_uop_prs2
                              : _GEN_287
                                  ? _slots_24_io_uop_prs2
                                  : _GEN_278
                                      ? _slots_23_io_uop_prs2
                                      : _GEN_269
                                          ? _slots_22_io_uop_prs2
                                          : _GEN_260
                                              ? _slots_21_io_uop_prs2
                                              : _GEN_251
                                                  ? _slots_20_io_uop_prs2
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_prs2
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_prs2
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_prs2
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_prs2
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_prs2
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_prs2
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_prs2
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_prs2
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_prs2
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_prs2
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_prs2
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_prs2
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_prs2
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_prs2
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_prs2
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_prs2
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_prs2
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_prs2
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_prs2
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_prs2
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:99:25, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_prs3 =
    _GEN_345
      ? _slots_31_io_uop_prs3
      : _GEN_340
          ? _slots_30_io_uop_prs3
          : _GEN_332
              ? _slots_29_io_uop_prs3
              : _GEN_323
                  ? _slots_28_io_uop_prs3
                  : _GEN_314
                      ? _slots_27_io_uop_prs3
                      : _GEN_305
                          ? _slots_26_io_uop_prs3
                          : _GEN_296
                              ? _slots_25_io_uop_prs3
                              : _GEN_287
                                  ? _slots_24_io_uop_prs3
                                  : _GEN_278
                                      ? _slots_23_io_uop_prs3
                                      : _GEN_269
                                          ? _slots_22_io_uop_prs3
                                          : _GEN_260
                                              ? _slots_21_io_uop_prs3
                                              : _GEN_251
                                                  ? _slots_20_io_uop_prs3
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_prs3
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_prs3
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_prs3
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_prs3
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_prs3
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_prs3
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_prs3
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_prs3
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_prs3
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_prs3
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_prs3
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_prs3
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_prs3
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_prs3
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_prs3
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_prs3
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_prs3
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_prs3
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_prs3
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_prs3
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:100:25, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_ppred =
    _GEN_345
      ? _slots_31_io_uop_ppred
      : _GEN_340
          ? _slots_30_io_uop_ppred
          : _GEN_332
              ? _slots_29_io_uop_ppred
              : _GEN_323
                  ? _slots_28_io_uop_ppred
                  : _GEN_314
                      ? _slots_27_io_uop_ppred
                      : _GEN_305
                          ? _slots_26_io_uop_ppred
                          : _GEN_296
                              ? _slots_25_io_uop_ppred
                              : _GEN_287
                                  ? _slots_24_io_uop_ppred
                                  : _GEN_278
                                      ? _slots_23_io_uop_ppred
                                      : _GEN_269
                                          ? _slots_22_io_uop_ppred
                                          : _GEN_260
                                              ? _slots_21_io_uop_ppred
                                              : _GEN_251
                                                  ? _slots_20_io_uop_ppred
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_ppred
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_ppred
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_ppred
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_ppred
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_ppred
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_ppred
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_ppred
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_ppred
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_ppred
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_ppred
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_ppred
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_ppred
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_ppred
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_ppred
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_ppred
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_ppred
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_ppred
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_ppred
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_ppred
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_ppred
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_1_prs1_busy =
    _GEN_345
      ? _slots_31_io_uop_prs1_busy
      : _GEN_340
          ? _slots_30_io_uop_prs1_busy
          : _GEN_332
              ? _slots_29_io_uop_prs1_busy
              : _GEN_323
                  ? _slots_28_io_uop_prs1_busy
                  : _GEN_314
                      ? _slots_27_io_uop_prs1_busy
                      : _GEN_305
                          ? _slots_26_io_uop_prs1_busy
                          : _GEN_296
                              ? _slots_25_io_uop_prs1_busy
                              : _GEN_287
                                  ? _slots_24_io_uop_prs1_busy
                                  : _GEN_278
                                      ? _slots_23_io_uop_prs1_busy
                                      : _GEN_269
                                          ? _slots_22_io_uop_prs1_busy
                                          : _GEN_260
                                              ? _slots_21_io_uop_prs1_busy
                                              : _GEN_251
                                                  ? _slots_20_io_uop_prs1_busy
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_prs1_busy
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_prs1_busy
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_prs1_busy
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_prs1_busy
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_prs1_busy
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_prs1_busy
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_prs1_busy
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_prs1_busy
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_prs1_busy
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_prs1_busy
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_prs1_busy
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_prs1_busy
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_prs1_busy
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_prs1_busy
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_prs1_busy
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_prs1_busy
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_prs1_busy
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_prs1_busy
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_prs1_busy
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_prs1_busy;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_prs2_busy =
    _GEN_345
      ? _slots_31_io_uop_prs2_busy
      : _GEN_340
          ? _slots_30_io_uop_prs2_busy
          : _GEN_332
              ? _slots_29_io_uop_prs2_busy
              : _GEN_323
                  ? _slots_28_io_uop_prs2_busy
                  : _GEN_314
                      ? _slots_27_io_uop_prs2_busy
                      : _GEN_305
                          ? _slots_26_io_uop_prs2_busy
                          : _GEN_296
                              ? _slots_25_io_uop_prs2_busy
                              : _GEN_287
                                  ? _slots_24_io_uop_prs2_busy
                                  : _GEN_278
                                      ? _slots_23_io_uop_prs2_busy
                                      : _GEN_269
                                          ? _slots_22_io_uop_prs2_busy
                                          : _GEN_260
                                              ? _slots_21_io_uop_prs2_busy
                                              : _GEN_251
                                                  ? _slots_20_io_uop_prs2_busy
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_prs2_busy
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_prs2_busy
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_prs2_busy
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_prs2_busy
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_prs2_busy
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_prs2_busy
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_prs2_busy
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_prs2_busy
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_prs2_busy
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_prs2_busy
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_prs2_busy
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_prs2_busy
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_prs2_busy
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_prs2_busy
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_prs2_busy
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_prs2_busy
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_prs2_busy
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_prs2_busy
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_prs2_busy
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_prs2_busy;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_prs3_busy =
    _GEN_345
      ? _slots_31_io_uop_prs3_busy
      : _GEN_340
          ? _slots_30_io_uop_prs3_busy
          : _GEN_332
              ? _slots_29_io_uop_prs3_busy
              : _GEN_323
                  ? _slots_28_io_uop_prs3_busy
                  : _GEN_314
                      ? _slots_27_io_uop_prs3_busy
                      : _GEN_305
                          ? _slots_26_io_uop_prs3_busy
                          : _GEN_296
                              ? _slots_25_io_uop_prs3_busy
                              : _GEN_287
                                  ? _slots_24_io_uop_prs3_busy
                                  : _GEN_278
                                      ? _slots_23_io_uop_prs3_busy
                                      : _GEN_269
                                          ? _slots_22_io_uop_prs3_busy
                                          : _GEN_260
                                              ? _slots_21_io_uop_prs3_busy
                                              : _GEN_251
                                                  ? _slots_20_io_uop_prs3_busy
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_prs3_busy
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_prs3_busy
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_prs3_busy
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_prs3_busy
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_prs3_busy
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_prs3_busy
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_prs3_busy
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_prs3_busy
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_prs3_busy
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_prs3_busy
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_prs3_busy
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_prs3_busy
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_prs3_busy
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_prs3_busy
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_prs3_busy
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_prs3_busy
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_prs3_busy
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_prs3_busy
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_prs3_busy
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_prs3_busy;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_ppred_busy =
    _GEN_345
      ? _slots_31_io_uop_ppred_busy
      : _GEN_340
          ? _slots_30_io_uop_ppred_busy
          : _GEN_332
              ? _slots_29_io_uop_ppred_busy
              : _GEN_323
                  ? _slots_28_io_uop_ppred_busy
                  : _GEN_314
                      ? _slots_27_io_uop_ppred_busy
                      : _GEN_305
                          ? _slots_26_io_uop_ppred_busy
                          : _GEN_296
                              ? _slots_25_io_uop_ppred_busy
                              : _GEN_287
                                  ? _slots_24_io_uop_ppred_busy
                                  : _GEN_278
                                      ? _slots_23_io_uop_ppred_busy
                                      : _GEN_269
                                          ? _slots_22_io_uop_ppred_busy
                                          : _GEN_260
                                              ? _slots_21_io_uop_ppred_busy
                                              : _GEN_251
                                                  ? _slots_20_io_uop_ppred_busy
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_ppred_busy
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_ppred_busy
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_ppred_busy
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_ppred_busy
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_ppred_busy
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_ppred_busy
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_ppred_busy
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_ppred_busy
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_ppred_busy
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_ppred_busy
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_ppred_busy
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_ppred_busy
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_ppred_busy
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_ppred_busy
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_ppred_busy
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_ppred_busy
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_ppred_busy
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_ppred_busy
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_ppred_busy
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_ppred_busy;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_stale_pdst =
    _GEN_345
      ? _slots_31_io_uop_stale_pdst
      : _GEN_340
          ? _slots_30_io_uop_stale_pdst
          : _GEN_332
              ? _slots_29_io_uop_stale_pdst
              : _GEN_323
                  ? _slots_28_io_uop_stale_pdst
                  : _GEN_314
                      ? _slots_27_io_uop_stale_pdst
                      : _GEN_305
                          ? _slots_26_io_uop_stale_pdst
                          : _GEN_296
                              ? _slots_25_io_uop_stale_pdst
                              : _GEN_287
                                  ? _slots_24_io_uop_stale_pdst
                                  : _GEN_278
                                      ? _slots_23_io_uop_stale_pdst
                                      : _GEN_269
                                          ? _slots_22_io_uop_stale_pdst
                                          : _GEN_260
                                              ? _slots_21_io_uop_stale_pdst
                                              : _GEN_251
                                                  ? _slots_20_io_uop_stale_pdst
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_stale_pdst
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_stale_pdst
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_stale_pdst
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_stale_pdst
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_stale_pdst
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_stale_pdst
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_stale_pdst
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_stale_pdst
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_stale_pdst
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_stale_pdst
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_stale_pdst
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_stale_pdst
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_stale_pdst
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_stale_pdst
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_stale_pdst
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_stale_pdst
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_stale_pdst
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_stale_pdst
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_stale_pdst
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_stale_pdst
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_exception =
    _GEN_345
      ? _slots_31_io_uop_exception
      : _GEN_340
          ? _slots_30_io_uop_exception
          : _GEN_332
              ? _slots_29_io_uop_exception
              : _GEN_323
                  ? _slots_28_io_uop_exception
                  : _GEN_314
                      ? _slots_27_io_uop_exception
                      : _GEN_305
                          ? _slots_26_io_uop_exception
                          : _GEN_296
                              ? _slots_25_io_uop_exception
                              : _GEN_287
                                  ? _slots_24_io_uop_exception
                                  : _GEN_278
                                      ? _slots_23_io_uop_exception
                                      : _GEN_269
                                          ? _slots_22_io_uop_exception
                                          : _GEN_260
                                              ? _slots_21_io_uop_exception
                                              : _GEN_251
                                                  ? _slots_20_io_uop_exception
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_exception
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_exception
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_exception
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_exception
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_exception
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_exception
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_exception
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_exception
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_exception
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_exception
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_exception
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_exception
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_exception
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_exception
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_exception
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_exception
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_exception
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_exception
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_exception
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_exception;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_exc_cause =
    _GEN_345
      ? _slots_31_io_uop_exc_cause
      : _GEN_340
          ? _slots_30_io_uop_exc_cause
          : _GEN_332
              ? _slots_29_io_uop_exc_cause
              : _GEN_323
                  ? _slots_28_io_uop_exc_cause
                  : _GEN_314
                      ? _slots_27_io_uop_exc_cause
                      : _GEN_305
                          ? _slots_26_io_uop_exc_cause
                          : _GEN_296
                              ? _slots_25_io_uop_exc_cause
                              : _GEN_287
                                  ? _slots_24_io_uop_exc_cause
                                  : _GEN_278
                                      ? _slots_23_io_uop_exc_cause
                                      : _GEN_269
                                          ? _slots_22_io_uop_exc_cause
                                          : _GEN_260
                                              ? _slots_21_io_uop_exc_cause
                                              : _GEN_251
                                                  ? _slots_20_io_uop_exc_cause
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_exc_cause
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_exc_cause
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_exc_cause
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_exc_cause
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_exc_cause
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_exc_cause
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_exc_cause
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_exc_cause
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_exc_cause
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_exc_cause
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_exc_cause
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_exc_cause
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_exc_cause
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_exc_cause
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_exc_cause
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_exc_cause
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_exc_cause
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_exc_cause
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_exc_cause
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_exc_cause
                                                                                                                                  : 64'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_bypassable =
    _GEN_345
      ? _slots_31_io_uop_bypassable
      : _GEN_340
          ? _slots_30_io_uop_bypassable
          : _GEN_332
              ? _slots_29_io_uop_bypassable
              : _GEN_323
                  ? _slots_28_io_uop_bypassable
                  : _GEN_314
                      ? _slots_27_io_uop_bypassable
                      : _GEN_305
                          ? _slots_26_io_uop_bypassable
                          : _GEN_296
                              ? _slots_25_io_uop_bypassable
                              : _GEN_287
                                  ? _slots_24_io_uop_bypassable
                                  : _GEN_278
                                      ? _slots_23_io_uop_bypassable
                                      : _GEN_269
                                          ? _slots_22_io_uop_bypassable
                                          : _GEN_260
                                              ? _slots_21_io_uop_bypassable
                                              : _GEN_251
                                                  ? _slots_20_io_uop_bypassable
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_bypassable
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_bypassable
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_bypassable
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_bypassable
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_bypassable
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_bypassable
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_bypassable
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_bypassable
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_bypassable
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_bypassable
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_bypassable
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_bypassable
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_bypassable
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_bypassable
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_bypassable
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_bypassable
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_bypassable
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_bypassable
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_bypassable
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_bypassable;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_mem_cmd =
    _GEN_345
      ? _slots_31_io_uop_mem_cmd
      : _GEN_340
          ? _slots_30_io_uop_mem_cmd
          : _GEN_332
              ? _slots_29_io_uop_mem_cmd
              : _GEN_323
                  ? _slots_28_io_uop_mem_cmd
                  : _GEN_314
                      ? _slots_27_io_uop_mem_cmd
                      : _GEN_305
                          ? _slots_26_io_uop_mem_cmd
                          : _GEN_296
                              ? _slots_25_io_uop_mem_cmd
                              : _GEN_287
                                  ? _slots_24_io_uop_mem_cmd
                                  : _GEN_278
                                      ? _slots_23_io_uop_mem_cmd
                                      : _GEN_269
                                          ? _slots_22_io_uop_mem_cmd
                                          : _GEN_260
                                              ? _slots_21_io_uop_mem_cmd
                                              : _GEN_251
                                                  ? _slots_20_io_uop_mem_cmd
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_mem_cmd
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_mem_cmd
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_mem_cmd
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_mem_cmd
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_mem_cmd
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_mem_cmd
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_mem_cmd
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_mem_cmd
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_mem_cmd
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_mem_cmd
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_mem_cmd
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_mem_cmd
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_mem_cmd
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_mem_cmd
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_mem_cmd
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_mem_cmd
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_mem_cmd
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_mem_cmd
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_mem_cmd
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_mem_cmd
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_1_mem_size =
    _GEN_345
      ? _slots_31_io_uop_mem_size
      : _GEN_340
          ? _slots_30_io_uop_mem_size
          : _GEN_332
              ? _slots_29_io_uop_mem_size
              : _GEN_323
                  ? _slots_28_io_uop_mem_size
                  : _GEN_314
                      ? _slots_27_io_uop_mem_size
                      : _GEN_305
                          ? _slots_26_io_uop_mem_size
                          : _GEN_296
                              ? _slots_25_io_uop_mem_size
                              : _GEN_287
                                  ? _slots_24_io_uop_mem_size
                                  : _GEN_278
                                      ? _slots_23_io_uop_mem_size
                                      : _GEN_269
                                          ? _slots_22_io_uop_mem_size
                                          : _GEN_260
                                              ? _slots_21_io_uop_mem_size
                                              : _GEN_251
                                                  ? _slots_20_io_uop_mem_size
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_mem_size
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_mem_size
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_mem_size
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_mem_size
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_mem_size
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_mem_size
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_mem_size
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_mem_size
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_mem_size
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_mem_size
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_mem_size
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_mem_size
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_mem_size
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_mem_size
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_mem_size
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_mem_size
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_mem_size
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_mem_size
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_mem_size
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_mem_size
                                                                                                                                  : 2'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:127:84, :153:73
  assign io_iss_uops_1_mem_signed =
    _GEN_345
      ? _slots_31_io_uop_mem_signed
      : _GEN_340
          ? _slots_30_io_uop_mem_signed
          : _GEN_332
              ? _slots_29_io_uop_mem_signed
              : _GEN_323
                  ? _slots_28_io_uop_mem_signed
                  : _GEN_314
                      ? _slots_27_io_uop_mem_signed
                      : _GEN_305
                          ? _slots_26_io_uop_mem_signed
                          : _GEN_296
                              ? _slots_25_io_uop_mem_signed
                              : _GEN_287
                                  ? _slots_24_io_uop_mem_signed
                                  : _GEN_278
                                      ? _slots_23_io_uop_mem_signed
                                      : _GEN_269
                                          ? _slots_22_io_uop_mem_signed
                                          : _GEN_260
                                              ? _slots_21_io_uop_mem_signed
                                              : _GEN_251
                                                  ? _slots_20_io_uop_mem_signed
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_mem_signed
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_mem_signed
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_mem_signed
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_mem_signed
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_mem_signed
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_mem_signed
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_mem_signed
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_mem_signed
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_mem_signed
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_mem_signed
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_mem_signed
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_mem_signed
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_mem_signed
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_mem_signed
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_mem_signed
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_mem_signed
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_mem_signed
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_mem_signed
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_mem_signed
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_mem_signed;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_fence =
    _GEN_345
      ? _slots_31_io_uop_is_fence
      : _GEN_340
          ? _slots_30_io_uop_is_fence
          : _GEN_332
              ? _slots_29_io_uop_is_fence
              : _GEN_323
                  ? _slots_28_io_uop_is_fence
                  : _GEN_314
                      ? _slots_27_io_uop_is_fence
                      : _GEN_305
                          ? _slots_26_io_uop_is_fence
                          : _GEN_296
                              ? _slots_25_io_uop_is_fence
                              : _GEN_287
                                  ? _slots_24_io_uop_is_fence
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_fence
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_fence
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_fence
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_fence
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_fence
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_fence
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_fence
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_fence
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_fence
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_fence
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_fence
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_fence
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_fence
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_fence
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_fence
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_fence
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_fence
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_fence
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_fence
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_fence
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_fence
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_fence
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_fence
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_fence;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_fencei =
    _GEN_345
      ? _slots_31_io_uop_is_fencei
      : _GEN_340
          ? _slots_30_io_uop_is_fencei
          : _GEN_332
              ? _slots_29_io_uop_is_fencei
              : _GEN_323
                  ? _slots_28_io_uop_is_fencei
                  : _GEN_314
                      ? _slots_27_io_uop_is_fencei
                      : _GEN_305
                          ? _slots_26_io_uop_is_fencei
                          : _GEN_296
                              ? _slots_25_io_uop_is_fencei
                              : _GEN_287
                                  ? _slots_24_io_uop_is_fencei
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_fencei
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_fencei
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_fencei
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_fencei
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_fencei
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_fencei
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_fencei
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_fencei
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_fencei
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_fencei
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_fencei
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_fencei
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_fencei
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_fencei
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_fencei
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_fencei
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_fencei
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_fencei
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_fencei
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_fencei
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_fencei
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_fencei
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_fencei
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_fencei;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_amo =
    _GEN_345
      ? _slots_31_io_uop_is_amo
      : _GEN_340
          ? _slots_30_io_uop_is_amo
          : _GEN_332
              ? _slots_29_io_uop_is_amo
              : _GEN_323
                  ? _slots_28_io_uop_is_amo
                  : _GEN_314
                      ? _slots_27_io_uop_is_amo
                      : _GEN_305
                          ? _slots_26_io_uop_is_amo
                          : _GEN_296
                              ? _slots_25_io_uop_is_amo
                              : _GEN_287
                                  ? _slots_24_io_uop_is_amo
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_amo
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_amo
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_amo
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_amo
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_amo
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_amo
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_amo
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_amo
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_amo
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_amo
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_amo
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_amo
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_amo
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_amo
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_amo
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_amo
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_amo
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_amo
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_amo
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_amo
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_amo
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_amo
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_amo
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_amo;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_uses_ldq =
    _GEN_345
      ? _slots_31_io_uop_uses_ldq
      : _GEN_340
          ? _slots_30_io_uop_uses_ldq
          : _GEN_332
              ? _slots_29_io_uop_uses_ldq
              : _GEN_323
                  ? _slots_28_io_uop_uses_ldq
                  : _GEN_314
                      ? _slots_27_io_uop_uses_ldq
                      : _GEN_305
                          ? _slots_26_io_uop_uses_ldq
                          : _GEN_296
                              ? _slots_25_io_uop_uses_ldq
                              : _GEN_287
                                  ? _slots_24_io_uop_uses_ldq
                                  : _GEN_278
                                      ? _slots_23_io_uop_uses_ldq
                                      : _GEN_269
                                          ? _slots_22_io_uop_uses_ldq
                                          : _GEN_260
                                              ? _slots_21_io_uop_uses_ldq
                                              : _GEN_251
                                                  ? _slots_20_io_uop_uses_ldq
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_uses_ldq
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_uses_ldq
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_uses_ldq
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_uses_ldq
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_uses_ldq
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_uses_ldq
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_uses_ldq
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_uses_ldq
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_uses_ldq
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_uses_ldq
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_uses_ldq
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_uses_ldq
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_uses_ldq
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_uses_ldq
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_uses_ldq
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_uses_ldq
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_uses_ldq
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_uses_ldq
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_uses_ldq
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_uses_ldq;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_uses_stq =
    _GEN_345
      ? _slots_31_io_uop_uses_stq
      : _GEN_340
          ? _slots_30_io_uop_uses_stq
          : _GEN_332
              ? _slots_29_io_uop_uses_stq
              : _GEN_323
                  ? _slots_28_io_uop_uses_stq
                  : _GEN_314
                      ? _slots_27_io_uop_uses_stq
                      : _GEN_305
                          ? _slots_26_io_uop_uses_stq
                          : _GEN_296
                              ? _slots_25_io_uop_uses_stq
                              : _GEN_287
                                  ? _slots_24_io_uop_uses_stq
                                  : _GEN_278
                                      ? _slots_23_io_uop_uses_stq
                                      : _GEN_269
                                          ? _slots_22_io_uop_uses_stq
                                          : _GEN_260
                                              ? _slots_21_io_uop_uses_stq
                                              : _GEN_251
                                                  ? _slots_20_io_uop_uses_stq
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_uses_stq
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_uses_stq
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_uses_stq
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_uses_stq
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_uses_stq
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_uses_stq
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_uses_stq
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_uses_stq
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_uses_stq
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_uses_stq
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_uses_stq
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_uses_stq
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_uses_stq
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_uses_stq
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_uses_stq
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_uses_stq
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_uses_stq
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_uses_stq
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_uses_stq
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_uses_stq;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_sys_pc2epc =
    _GEN_345
      ? _slots_31_io_uop_is_sys_pc2epc
      : _GEN_340
          ? _slots_30_io_uop_is_sys_pc2epc
          : _GEN_332
              ? _slots_29_io_uop_is_sys_pc2epc
              : _GEN_323
                  ? _slots_28_io_uop_is_sys_pc2epc
                  : _GEN_314
                      ? _slots_27_io_uop_is_sys_pc2epc
                      : _GEN_305
                          ? _slots_26_io_uop_is_sys_pc2epc
                          : _GEN_296
                              ? _slots_25_io_uop_is_sys_pc2epc
                              : _GEN_287
                                  ? _slots_24_io_uop_is_sys_pc2epc
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_sys_pc2epc
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_sys_pc2epc
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_sys_pc2epc
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_sys_pc2epc
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_sys_pc2epc
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_sys_pc2epc
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_sys_pc2epc
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_sys_pc2epc
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_sys_pc2epc
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_sys_pc2epc
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_sys_pc2epc
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_sys_pc2epc
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_sys_pc2epc
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_sys_pc2epc
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_sys_pc2epc
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_sys_pc2epc
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_sys_pc2epc
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_sys_pc2epc
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_sys_pc2epc
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_sys_pc2epc
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_sys_pc2epc
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_sys_pc2epc
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_sys_pc2epc
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_sys_pc2epc;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_is_unique =
    _GEN_345
      ? _slots_31_io_uop_is_unique
      : _GEN_340
          ? _slots_30_io_uop_is_unique
          : _GEN_332
              ? _slots_29_io_uop_is_unique
              : _GEN_323
                  ? _slots_28_io_uop_is_unique
                  : _GEN_314
                      ? _slots_27_io_uop_is_unique
                      : _GEN_305
                          ? _slots_26_io_uop_is_unique
                          : _GEN_296
                              ? _slots_25_io_uop_is_unique
                              : _GEN_287
                                  ? _slots_24_io_uop_is_unique
                                  : _GEN_278
                                      ? _slots_23_io_uop_is_unique
                                      : _GEN_269
                                          ? _slots_22_io_uop_is_unique
                                          : _GEN_260
                                              ? _slots_21_io_uop_is_unique
                                              : _GEN_251
                                                  ? _slots_20_io_uop_is_unique
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_is_unique
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_is_unique
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_is_unique
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_is_unique
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_is_unique
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_is_unique
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_is_unique
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_is_unique
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_is_unique
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_is_unique
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_is_unique
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_is_unique
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_is_unique
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_is_unique
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_is_unique
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_is_unique
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_is_unique
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_is_unique
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_is_unique
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_is_unique;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_flush_on_commit =
    _GEN_345
      ? _slots_31_io_uop_flush_on_commit
      : _GEN_340
          ? _slots_30_io_uop_flush_on_commit
          : _GEN_332
              ? _slots_29_io_uop_flush_on_commit
              : _GEN_323
                  ? _slots_28_io_uop_flush_on_commit
                  : _GEN_314
                      ? _slots_27_io_uop_flush_on_commit
                      : _GEN_305
                          ? _slots_26_io_uop_flush_on_commit
                          : _GEN_296
                              ? _slots_25_io_uop_flush_on_commit
                              : _GEN_287
                                  ? _slots_24_io_uop_flush_on_commit
                                  : _GEN_278
                                      ? _slots_23_io_uop_flush_on_commit
                                      : _GEN_269
                                          ? _slots_22_io_uop_flush_on_commit
                                          : _GEN_260
                                              ? _slots_21_io_uop_flush_on_commit
                                              : _GEN_251
                                                  ? _slots_20_io_uop_flush_on_commit
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_flush_on_commit
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_flush_on_commit
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_flush_on_commit
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_flush_on_commit
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_flush_on_commit
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_flush_on_commit
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_flush_on_commit
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_flush_on_commit
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_flush_on_commit
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_flush_on_commit
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_flush_on_commit
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_flush_on_commit
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_flush_on_commit
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_flush_on_commit
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_flush_on_commit
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_flush_on_commit
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_flush_on_commit
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_flush_on_commit
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_flush_on_commit
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_flush_on_commit;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_ldst_is_rs1 =
    _GEN_345
      ? _slots_31_io_uop_ldst_is_rs1
      : _GEN_340
          ? _slots_30_io_uop_ldst_is_rs1
          : _GEN_332
              ? _slots_29_io_uop_ldst_is_rs1
              : _GEN_323
                  ? _slots_28_io_uop_ldst_is_rs1
                  : _GEN_314
                      ? _slots_27_io_uop_ldst_is_rs1
                      : _GEN_305
                          ? _slots_26_io_uop_ldst_is_rs1
                          : _GEN_296
                              ? _slots_25_io_uop_ldst_is_rs1
                              : _GEN_287
                                  ? _slots_24_io_uop_ldst_is_rs1
                                  : _GEN_278
                                      ? _slots_23_io_uop_ldst_is_rs1
                                      : _GEN_269
                                          ? _slots_22_io_uop_ldst_is_rs1
                                          : _GEN_260
                                              ? _slots_21_io_uop_ldst_is_rs1
                                              : _GEN_251
                                                  ? _slots_20_io_uop_ldst_is_rs1
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_ldst_is_rs1
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_ldst_is_rs1
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_ldst_is_rs1
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_ldst_is_rs1
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_ldst_is_rs1
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_ldst_is_rs1
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_ldst_is_rs1
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_ldst_is_rs1
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_ldst_is_rs1
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_ldst_is_rs1
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_ldst_is_rs1
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_ldst_is_rs1
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_ldst_is_rs1
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_ldst_is_rs1
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_ldst_is_rs1
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_ldst_is_rs1
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_ldst_is_rs1
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_ldst_is_rs1
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_ldst_is_rs1
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_ldst_is_rs1;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_ldst =
    _GEN_345
      ? _slots_31_io_uop_ldst
      : _GEN_340
          ? _slots_30_io_uop_ldst
          : _GEN_332
              ? _slots_29_io_uop_ldst
              : _GEN_323
                  ? _slots_28_io_uop_ldst
                  : _GEN_314
                      ? _slots_27_io_uop_ldst
                      : _GEN_305
                          ? _slots_26_io_uop_ldst
                          : _GEN_296
                              ? _slots_25_io_uop_ldst
                              : _GEN_287
                                  ? _slots_24_io_uop_ldst
                                  : _GEN_278
                                      ? _slots_23_io_uop_ldst
                                      : _GEN_269
                                          ? _slots_22_io_uop_ldst
                                          : _GEN_260
                                              ? _slots_21_io_uop_ldst
                                              : _GEN_251
                                                  ? _slots_20_io_uop_ldst
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_ldst
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_ldst
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_ldst
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_ldst
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_ldst
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_ldst
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_ldst
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_ldst
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_ldst
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_ldst
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_ldst
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_ldst
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_ldst
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_ldst
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_ldst
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_ldst
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_ldst
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_ldst
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_ldst
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_ldst
                                                                                                                                  : 6'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_lrs1 =
    _GEN_345
      ? _slots_31_io_uop_lrs1
      : _GEN_340
          ? _slots_30_io_uop_lrs1
          : _GEN_332
              ? _slots_29_io_uop_lrs1
              : _GEN_323
                  ? _slots_28_io_uop_lrs1
                  : _GEN_314
                      ? _slots_27_io_uop_lrs1
                      : _GEN_305
                          ? _slots_26_io_uop_lrs1
                          : _GEN_296
                              ? _slots_25_io_uop_lrs1
                              : _GEN_287
                                  ? _slots_24_io_uop_lrs1
                                  : _GEN_278
                                      ? _slots_23_io_uop_lrs1
                                      : _GEN_269
                                          ? _slots_22_io_uop_lrs1
                                          : _GEN_260
                                              ? _slots_21_io_uop_lrs1
                                              : _GEN_251
                                                  ? _slots_20_io_uop_lrs1
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_lrs1
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_lrs1
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_lrs1
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_lrs1
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_lrs1
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_lrs1
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_lrs1
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_lrs1
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_lrs1
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_lrs1
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_lrs1
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_lrs1
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_lrs1
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_lrs1
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_lrs1
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_lrs1
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_lrs1
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_lrs1
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_lrs1
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_lrs1
                                                                                                                                  : 6'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_lrs2 =
    _GEN_345
      ? _slots_31_io_uop_lrs2
      : _GEN_340
          ? _slots_30_io_uop_lrs2
          : _GEN_332
              ? _slots_29_io_uop_lrs2
              : _GEN_323
                  ? _slots_28_io_uop_lrs2
                  : _GEN_314
                      ? _slots_27_io_uop_lrs2
                      : _GEN_305
                          ? _slots_26_io_uop_lrs2
                          : _GEN_296
                              ? _slots_25_io_uop_lrs2
                              : _GEN_287
                                  ? _slots_24_io_uop_lrs2
                                  : _GEN_278
                                      ? _slots_23_io_uop_lrs2
                                      : _GEN_269
                                          ? _slots_22_io_uop_lrs2
                                          : _GEN_260
                                              ? _slots_21_io_uop_lrs2
                                              : _GEN_251
                                                  ? _slots_20_io_uop_lrs2
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_lrs2
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_lrs2
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_lrs2
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_lrs2
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_lrs2
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_lrs2
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_lrs2
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_lrs2
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_lrs2
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_lrs2
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_lrs2
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_lrs2
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_lrs2
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_lrs2
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_lrs2
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_lrs2
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_lrs2
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_lrs2
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_lrs2
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_lrs2
                                                                                                                                  : 6'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_lrs3 =
    _GEN_345
      ? _slots_31_io_uop_lrs3
      : _GEN_340
          ? _slots_30_io_uop_lrs3
          : _GEN_332
              ? _slots_29_io_uop_lrs3
              : _GEN_323
                  ? _slots_28_io_uop_lrs3
                  : _GEN_314
                      ? _slots_27_io_uop_lrs3
                      : _GEN_305
                          ? _slots_26_io_uop_lrs3
                          : _GEN_296
                              ? _slots_25_io_uop_lrs3
                              : _GEN_287
                                  ? _slots_24_io_uop_lrs3
                                  : _GEN_278
                                      ? _slots_23_io_uop_lrs3
                                      : _GEN_269
                                          ? _slots_22_io_uop_lrs3
                                          : _GEN_260
                                              ? _slots_21_io_uop_lrs3
                                              : _GEN_251
                                                  ? _slots_20_io_uop_lrs3
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_lrs3
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_lrs3
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_lrs3
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_lrs3
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_lrs3
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_lrs3
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_lrs3
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_lrs3
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_lrs3
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_lrs3
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_lrs3
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_lrs3
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_lrs3
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_lrs3
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_lrs3
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_lrs3
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_lrs3
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_lrs3
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_lrs3
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_lrs3
                                                                                                                                  : 6'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_ldst_val =
    _GEN_345
      ? _slots_31_io_uop_ldst_val
      : _GEN_340
          ? _slots_30_io_uop_ldst_val
          : _GEN_332
              ? _slots_29_io_uop_ldst_val
              : _GEN_323
                  ? _slots_28_io_uop_ldst_val
                  : _GEN_314
                      ? _slots_27_io_uop_ldst_val
                      : _GEN_305
                          ? _slots_26_io_uop_ldst_val
                          : _GEN_296
                              ? _slots_25_io_uop_ldst_val
                              : _GEN_287
                                  ? _slots_24_io_uop_ldst_val
                                  : _GEN_278
                                      ? _slots_23_io_uop_ldst_val
                                      : _GEN_269
                                          ? _slots_22_io_uop_ldst_val
                                          : _GEN_260
                                              ? _slots_21_io_uop_ldst_val
                                              : _GEN_251
                                                  ? _slots_20_io_uop_ldst_val
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_ldst_val
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_ldst_val
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_ldst_val
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_ldst_val
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_ldst_val
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_ldst_val
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_ldst_val
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_ldst_val
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_ldst_val
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_ldst_val
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_ldst_val
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_ldst_val
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_ldst_val
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_ldst_val
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_ldst_val
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_ldst_val
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_ldst_val
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_ldst_val
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_ldst_val
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_ldst_val;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_dst_rtype =
    _GEN_345
      ? _slots_31_io_uop_dst_rtype
      : _GEN_340
          ? _slots_30_io_uop_dst_rtype
          : _GEN_332
              ? _slots_29_io_uop_dst_rtype
              : _GEN_323
                  ? _slots_28_io_uop_dst_rtype
                  : _GEN_314
                      ? _slots_27_io_uop_dst_rtype
                      : _GEN_305
                          ? _slots_26_io_uop_dst_rtype
                          : _GEN_296
                              ? _slots_25_io_uop_dst_rtype
                              : _GEN_287
                                  ? _slots_24_io_uop_dst_rtype
                                  : _GEN_278
                                      ? _slots_23_io_uop_dst_rtype
                                      : _GEN_269
                                          ? _slots_22_io_uop_dst_rtype
                                          : _GEN_260
                                              ? _slots_21_io_uop_dst_rtype
                                              : _GEN_251
                                                  ? _slots_20_io_uop_dst_rtype
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_dst_rtype
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_dst_rtype
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_dst_rtype
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_dst_rtype
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_dst_rtype
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_dst_rtype
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_dst_rtype
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_dst_rtype
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_dst_rtype
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_dst_rtype
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_dst_rtype
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_dst_rtype
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_dst_rtype
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_dst_rtype
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_dst_rtype
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_dst_rtype
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_dst_rtype
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_dst_rtype
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_dst_rtype
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_dst_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_1_lrs1_rtype =
    _GEN_345
      ? _slots_31_io_uop_lrs1_rtype
      : _GEN_340
          ? _slots_30_io_uop_lrs1_rtype
          : _GEN_332
              ? _slots_29_io_uop_lrs1_rtype
              : _GEN_323
                  ? _slots_28_io_uop_lrs1_rtype
                  : _GEN_314
                      ? _slots_27_io_uop_lrs1_rtype
                      : _GEN_305
                          ? _slots_26_io_uop_lrs1_rtype
                          : _GEN_296
                              ? _slots_25_io_uop_lrs1_rtype
                              : _GEN_287
                                  ? _slots_24_io_uop_lrs1_rtype
                                  : _GEN_278
                                      ? _slots_23_io_uop_lrs1_rtype
                                      : _GEN_269
                                          ? _slots_22_io_uop_lrs1_rtype
                                          : _GEN_260
                                              ? _slots_21_io_uop_lrs1_rtype
                                              : _GEN_251
                                                  ? _slots_20_io_uop_lrs1_rtype
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_lrs1_rtype
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_lrs1_rtype
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_lrs1_rtype
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_lrs1_rtype
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_lrs1_rtype
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_lrs1_rtype
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_lrs1_rtype
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_lrs1_rtype
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_lrs1_rtype
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_lrs1_rtype
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_lrs1_rtype
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_lrs1_rtype
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_lrs1_rtype
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_lrs1_rtype
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_lrs1_rtype
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_lrs1_rtype
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_lrs1_rtype
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_lrs1_rtype
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_lrs1_rtype
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_lrs1_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:101:31, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_1_lrs2_rtype =
    _GEN_345
      ? _slots_31_io_uop_lrs2_rtype
      : _GEN_340
          ? _slots_30_io_uop_lrs2_rtype
          : _GEN_332
              ? _slots_29_io_uop_lrs2_rtype
              : _GEN_323
                  ? _slots_28_io_uop_lrs2_rtype
                  : _GEN_314
                      ? _slots_27_io_uop_lrs2_rtype
                      : _GEN_305
                          ? _slots_26_io_uop_lrs2_rtype
                          : _GEN_296
                              ? _slots_25_io_uop_lrs2_rtype
                              : _GEN_287
                                  ? _slots_24_io_uop_lrs2_rtype
                                  : _GEN_278
                                      ? _slots_23_io_uop_lrs2_rtype
                                      : _GEN_269
                                          ? _slots_22_io_uop_lrs2_rtype
                                          : _GEN_260
                                              ? _slots_21_io_uop_lrs2_rtype
                                              : _GEN_251
                                                  ? _slots_20_io_uop_lrs2_rtype
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_lrs2_rtype
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_lrs2_rtype
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_lrs2_rtype
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_lrs2_rtype
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_lrs2_rtype
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_lrs2_rtype
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_lrs2_rtype
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_lrs2_rtype
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_lrs2_rtype
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_lrs2_rtype
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_lrs2_rtype
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_lrs2_rtype
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_lrs2_rtype
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_lrs2_rtype
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_lrs2_rtype
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_lrs2_rtype
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_lrs2_rtype
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_lrs2_rtype
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_lrs2_rtype
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_lrs2_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:102:31, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_1_frs3_en =
    _GEN_345
      ? _slots_31_io_uop_frs3_en
      : _GEN_340
          ? _slots_30_io_uop_frs3_en
          : _GEN_332
              ? _slots_29_io_uop_frs3_en
              : _GEN_323
                  ? _slots_28_io_uop_frs3_en
                  : _GEN_314
                      ? _slots_27_io_uop_frs3_en
                      : _GEN_305
                          ? _slots_26_io_uop_frs3_en
                          : _GEN_296
                              ? _slots_25_io_uop_frs3_en
                              : _GEN_287
                                  ? _slots_24_io_uop_frs3_en
                                  : _GEN_278
                                      ? _slots_23_io_uop_frs3_en
                                      : _GEN_269
                                          ? _slots_22_io_uop_frs3_en
                                          : _GEN_260
                                              ? _slots_21_io_uop_frs3_en
                                              : _GEN_251
                                                  ? _slots_20_io_uop_frs3_en
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_frs3_en
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_frs3_en
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_frs3_en
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_frs3_en
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_frs3_en
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_frs3_en
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_frs3_en
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_frs3_en
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_frs3_en
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_frs3_en
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_frs3_en
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_frs3_en
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_frs3_en
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_frs3_en
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_frs3_en
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_frs3_en
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_frs3_en
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_frs3_en
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_frs3_en
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_frs3_en;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_fp_val =
    _GEN_345
      ? _slots_31_io_uop_fp_val
      : _GEN_340
          ? _slots_30_io_uop_fp_val
          : _GEN_332
              ? _slots_29_io_uop_fp_val
              : _GEN_323
                  ? _slots_28_io_uop_fp_val
                  : _GEN_314
                      ? _slots_27_io_uop_fp_val
                      : _GEN_305
                          ? _slots_26_io_uop_fp_val
                          : _GEN_296
                              ? _slots_25_io_uop_fp_val
                              : _GEN_287
                                  ? _slots_24_io_uop_fp_val
                                  : _GEN_278
                                      ? _slots_23_io_uop_fp_val
                                      : _GEN_269
                                          ? _slots_22_io_uop_fp_val
                                          : _GEN_260
                                              ? _slots_21_io_uop_fp_val
                                              : _GEN_251
                                                  ? _slots_20_io_uop_fp_val
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_fp_val
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_fp_val
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_fp_val
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_fp_val
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_fp_val
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_fp_val
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_fp_val
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_fp_val
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_fp_val
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_fp_val
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_fp_val
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_fp_val
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_fp_val
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_fp_val
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_fp_val
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_fp_val
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_fp_val
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_fp_val
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_fp_val
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_fp_val;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_fp_single =
    _GEN_345
      ? _slots_31_io_uop_fp_single
      : _GEN_340
          ? _slots_30_io_uop_fp_single
          : _GEN_332
              ? _slots_29_io_uop_fp_single
              : _GEN_323
                  ? _slots_28_io_uop_fp_single
                  : _GEN_314
                      ? _slots_27_io_uop_fp_single
                      : _GEN_305
                          ? _slots_26_io_uop_fp_single
                          : _GEN_296
                              ? _slots_25_io_uop_fp_single
                              : _GEN_287
                                  ? _slots_24_io_uop_fp_single
                                  : _GEN_278
                                      ? _slots_23_io_uop_fp_single
                                      : _GEN_269
                                          ? _slots_22_io_uop_fp_single
                                          : _GEN_260
                                              ? _slots_21_io_uop_fp_single
                                              : _GEN_251
                                                  ? _slots_20_io_uop_fp_single
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_fp_single
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_fp_single
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_fp_single
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_fp_single
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_fp_single
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_fp_single
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_fp_single
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_fp_single
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_fp_single
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_fp_single
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_fp_single
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_fp_single
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_fp_single
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_fp_single
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_fp_single
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_fp_single
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_fp_single
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_fp_single
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_fp_single
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_fp_single;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_xcpt_pf_if =
    _GEN_345
      ? _slots_31_io_uop_xcpt_pf_if
      : _GEN_340
          ? _slots_30_io_uop_xcpt_pf_if
          : _GEN_332
              ? _slots_29_io_uop_xcpt_pf_if
              : _GEN_323
                  ? _slots_28_io_uop_xcpt_pf_if
                  : _GEN_314
                      ? _slots_27_io_uop_xcpt_pf_if
                      : _GEN_305
                          ? _slots_26_io_uop_xcpt_pf_if
                          : _GEN_296
                              ? _slots_25_io_uop_xcpt_pf_if
                              : _GEN_287
                                  ? _slots_24_io_uop_xcpt_pf_if
                                  : _GEN_278
                                      ? _slots_23_io_uop_xcpt_pf_if
                                      : _GEN_269
                                          ? _slots_22_io_uop_xcpt_pf_if
                                          : _GEN_260
                                              ? _slots_21_io_uop_xcpt_pf_if
                                              : _GEN_251
                                                  ? _slots_20_io_uop_xcpt_pf_if
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_xcpt_pf_if
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_xcpt_pf_if
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_xcpt_pf_if
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_xcpt_pf_if
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_xcpt_pf_if
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_xcpt_pf_if
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_xcpt_pf_if
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_xcpt_pf_if
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_xcpt_pf_if
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_xcpt_pf_if
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_xcpt_pf_if
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_xcpt_pf_if
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_xcpt_pf_if
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_xcpt_pf_if
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_xcpt_pf_if
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_xcpt_pf_if
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_xcpt_pf_if
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_xcpt_pf_if
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_xcpt_pf_if
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_xcpt_pf_if;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_xcpt_ae_if =
    _GEN_345
      ? _slots_31_io_uop_xcpt_ae_if
      : _GEN_340
          ? _slots_30_io_uop_xcpt_ae_if
          : _GEN_332
              ? _slots_29_io_uop_xcpt_ae_if
              : _GEN_323
                  ? _slots_28_io_uop_xcpt_ae_if
                  : _GEN_314
                      ? _slots_27_io_uop_xcpt_ae_if
                      : _GEN_305
                          ? _slots_26_io_uop_xcpt_ae_if
                          : _GEN_296
                              ? _slots_25_io_uop_xcpt_ae_if
                              : _GEN_287
                                  ? _slots_24_io_uop_xcpt_ae_if
                                  : _GEN_278
                                      ? _slots_23_io_uop_xcpt_ae_if
                                      : _GEN_269
                                          ? _slots_22_io_uop_xcpt_ae_if
                                          : _GEN_260
                                              ? _slots_21_io_uop_xcpt_ae_if
                                              : _GEN_251
                                                  ? _slots_20_io_uop_xcpt_ae_if
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_xcpt_ae_if
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_xcpt_ae_if
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_xcpt_ae_if
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_xcpt_ae_if
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_xcpt_ae_if
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_xcpt_ae_if
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_xcpt_ae_if
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_xcpt_ae_if
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_xcpt_ae_if
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_xcpt_ae_if
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_xcpt_ae_if
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_xcpt_ae_if
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_xcpt_ae_if
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_xcpt_ae_if
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_xcpt_ae_if
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_xcpt_ae_if
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_xcpt_ae_if
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_xcpt_ae_if
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_xcpt_ae_if
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_xcpt_ae_if;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_xcpt_ma_if =
    _GEN_345
      ? _slots_31_io_uop_xcpt_ma_if
      : _GEN_340
          ? _slots_30_io_uop_xcpt_ma_if
          : _GEN_332
              ? _slots_29_io_uop_xcpt_ma_if
              : _GEN_323
                  ? _slots_28_io_uop_xcpt_ma_if
                  : _GEN_314
                      ? _slots_27_io_uop_xcpt_ma_if
                      : _GEN_305
                          ? _slots_26_io_uop_xcpt_ma_if
                          : _GEN_296
                              ? _slots_25_io_uop_xcpt_ma_if
                              : _GEN_287
                                  ? _slots_24_io_uop_xcpt_ma_if
                                  : _GEN_278
                                      ? _slots_23_io_uop_xcpt_ma_if
                                      : _GEN_269
                                          ? _slots_22_io_uop_xcpt_ma_if
                                          : _GEN_260
                                              ? _slots_21_io_uop_xcpt_ma_if
                                              : _GEN_251
                                                  ? _slots_20_io_uop_xcpt_ma_if
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_xcpt_ma_if
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_xcpt_ma_if
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_xcpt_ma_if
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_xcpt_ma_if
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_xcpt_ma_if
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_xcpt_ma_if
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_xcpt_ma_if
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_xcpt_ma_if
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_xcpt_ma_if
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_xcpt_ma_if
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_xcpt_ma_if
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_xcpt_ma_if
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_xcpt_ma_if
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_xcpt_ma_if
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_xcpt_ma_if
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_xcpt_ma_if
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_xcpt_ma_if
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_xcpt_ma_if
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_xcpt_ma_if
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_xcpt_ma_if;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_bp_debug_if =
    _GEN_345
      ? _slots_31_io_uop_bp_debug_if
      : _GEN_340
          ? _slots_30_io_uop_bp_debug_if
          : _GEN_332
              ? _slots_29_io_uop_bp_debug_if
              : _GEN_323
                  ? _slots_28_io_uop_bp_debug_if
                  : _GEN_314
                      ? _slots_27_io_uop_bp_debug_if
                      : _GEN_305
                          ? _slots_26_io_uop_bp_debug_if
                          : _GEN_296
                              ? _slots_25_io_uop_bp_debug_if
                              : _GEN_287
                                  ? _slots_24_io_uop_bp_debug_if
                                  : _GEN_278
                                      ? _slots_23_io_uop_bp_debug_if
                                      : _GEN_269
                                          ? _slots_22_io_uop_bp_debug_if
                                          : _GEN_260
                                              ? _slots_21_io_uop_bp_debug_if
                                              : _GEN_251
                                                  ? _slots_20_io_uop_bp_debug_if
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_bp_debug_if
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_bp_debug_if
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_bp_debug_if
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_bp_debug_if
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_bp_debug_if
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_bp_debug_if
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_bp_debug_if
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_bp_debug_if
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_bp_debug_if
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_bp_debug_if
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_bp_debug_if
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_bp_debug_if
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_bp_debug_if
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_bp_debug_if
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_bp_debug_if
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_bp_debug_if
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_bp_debug_if
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_bp_debug_if
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_bp_debug_if
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_bp_debug_if;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_bp_xcpt_if =
    _GEN_345
      ? _slots_31_io_uop_bp_xcpt_if
      : _GEN_340
          ? _slots_30_io_uop_bp_xcpt_if
          : _GEN_332
              ? _slots_29_io_uop_bp_xcpt_if
              : _GEN_323
                  ? _slots_28_io_uop_bp_xcpt_if
                  : _GEN_314
                      ? _slots_27_io_uop_bp_xcpt_if
                      : _GEN_305
                          ? _slots_26_io_uop_bp_xcpt_if
                          : _GEN_296
                              ? _slots_25_io_uop_bp_xcpt_if
                              : _GEN_287
                                  ? _slots_24_io_uop_bp_xcpt_if
                                  : _GEN_278
                                      ? _slots_23_io_uop_bp_xcpt_if
                                      : _GEN_269
                                          ? _slots_22_io_uop_bp_xcpt_if
                                          : _GEN_260
                                              ? _slots_21_io_uop_bp_xcpt_if
                                              : _GEN_251
                                                  ? _slots_20_io_uop_bp_xcpt_if
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_bp_xcpt_if
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_bp_xcpt_if
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_bp_xcpt_if
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_bp_xcpt_if
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_bp_xcpt_if
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_bp_xcpt_if
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_bp_xcpt_if
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_bp_xcpt_if
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_bp_xcpt_if
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_bp_xcpt_if
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_bp_xcpt_if
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_bp_xcpt_if
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_bp_xcpt_if
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_bp_xcpt_if
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_bp_xcpt_if
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_bp_xcpt_if
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_bp_xcpt_if
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_bp_xcpt_if
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_bp_xcpt_if
                                                                                                                              : _GEN_74
                                                                                                                                & _slots_0_io_uop_bp_xcpt_if;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_1_debug_fsrc =
    _GEN_345
      ? _slots_31_io_uop_debug_fsrc
      : _GEN_340
          ? _slots_30_io_uop_debug_fsrc
          : _GEN_332
              ? _slots_29_io_uop_debug_fsrc
              : _GEN_323
                  ? _slots_28_io_uop_debug_fsrc
                  : _GEN_314
                      ? _slots_27_io_uop_debug_fsrc
                      : _GEN_305
                          ? _slots_26_io_uop_debug_fsrc
                          : _GEN_296
                              ? _slots_25_io_uop_debug_fsrc
                              : _GEN_287
                                  ? _slots_24_io_uop_debug_fsrc
                                  : _GEN_278
                                      ? _slots_23_io_uop_debug_fsrc
                                      : _GEN_269
                                          ? _slots_22_io_uop_debug_fsrc
                                          : _GEN_260
                                              ? _slots_21_io_uop_debug_fsrc
                                              : _GEN_251
                                                  ? _slots_20_io_uop_debug_fsrc
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_debug_fsrc
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_debug_fsrc
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_debug_fsrc
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_debug_fsrc
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_debug_fsrc
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_debug_fsrc
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_debug_fsrc
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_debug_fsrc
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_debug_fsrc
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_debug_fsrc
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_debug_fsrc
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_debug_fsrc
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_debug_fsrc
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_debug_fsrc
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_debug_fsrc
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_debug_fsrc
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_debug_fsrc
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_debug_fsrc
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_debug_fsrc
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_debug_fsrc
                                                                                                                                  : 2'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:127:84, :153:73
  assign io_iss_uops_1_debug_tsrc =
    _GEN_345
      ? _slots_31_io_uop_debug_tsrc
      : _GEN_340
          ? _slots_30_io_uop_debug_tsrc
          : _GEN_332
              ? _slots_29_io_uop_debug_tsrc
              : _GEN_323
                  ? _slots_28_io_uop_debug_tsrc
                  : _GEN_314
                      ? _slots_27_io_uop_debug_tsrc
                      : _GEN_305
                          ? _slots_26_io_uop_debug_tsrc
                          : _GEN_296
                              ? _slots_25_io_uop_debug_tsrc
                              : _GEN_287
                                  ? _slots_24_io_uop_debug_tsrc
                                  : _GEN_278
                                      ? _slots_23_io_uop_debug_tsrc
                                      : _GEN_269
                                          ? _slots_22_io_uop_debug_tsrc
                                          : _GEN_260
                                              ? _slots_21_io_uop_debug_tsrc
                                              : _GEN_251
                                                  ? _slots_20_io_uop_debug_tsrc
                                                  : _GEN_242
                                                      ? _slots_19_io_uop_debug_tsrc
                                                      : _GEN_233
                                                          ? _slots_18_io_uop_debug_tsrc
                                                          : _GEN_224
                                                              ? _slots_17_io_uop_debug_tsrc
                                                              : _GEN_215
                                                                  ? _slots_16_io_uop_debug_tsrc
                                                                  : _GEN_206
                                                                      ? _slots_15_io_uop_debug_tsrc
                                                                      : _GEN_197
                                                                          ? _slots_14_io_uop_debug_tsrc
                                                                          : _GEN_188
                                                                              ? _slots_13_io_uop_debug_tsrc
                                                                              : _GEN_179
                                                                                  ? _slots_12_io_uop_debug_tsrc
                                                                                  : _GEN_170
                                                                                      ? _slots_11_io_uop_debug_tsrc
                                                                                      : _GEN_161
                                                                                          ? _slots_10_io_uop_debug_tsrc
                                                                                          : _GEN_152
                                                                                              ? _slots_9_io_uop_debug_tsrc
                                                                                              : _GEN_143
                                                                                                  ? _slots_8_io_uop_debug_tsrc
                                                                                                  : _GEN_134
                                                                                                      ? _slots_7_io_uop_debug_tsrc
                                                                                                      : _GEN_125
                                                                                                          ? _slots_6_io_uop_debug_tsrc
                                                                                                          : _GEN_116
                                                                                                              ? _slots_5_io_uop_debug_tsrc
                                                                                                              : _GEN_107
                                                                                                                  ? _slots_4_io_uop_debug_tsrc
                                                                                                                  : _GEN_98
                                                                                                                      ? _slots_3_io_uop_debug_tsrc
                                                                                                                      : _GEN_89
                                                                                                                          ? _slots_2_io_uop_debug_tsrc
                                                                                                                          : _GEN_80
                                                                                                                              ? _slots_1_io_uop_debug_tsrc
                                                                                                                              : _GEN_74
                                                                                                                                  ? _slots_0_io_uop_debug_tsrc
                                                                                                                                  : 2'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:127:84, :153:73
  assign io_iss_uops_2_uopc =
    _GEN_346
      ? _slots_31_io_uop_uopc
      : _GEN_343
          ? _slots_30_io_uop_uopc
          : _GEN_335
              ? _slots_29_io_uop_uopc
              : _GEN_326
                  ? _slots_28_io_uop_uopc
                  : _GEN_317
                      ? _slots_27_io_uop_uopc
                      : _GEN_308
                          ? _slots_26_io_uop_uopc
                          : _GEN_299
                              ? _slots_25_io_uop_uopc
                              : _GEN_290
                                  ? _slots_24_io_uop_uopc
                                  : _GEN_281
                                      ? _slots_23_io_uop_uopc
                                      : _GEN_272
                                          ? _slots_22_io_uop_uopc
                                          : _GEN_263
                                              ? _slots_21_io_uop_uopc
                                              : _GEN_254
                                                  ? _slots_20_io_uop_uopc
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_uopc
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_uopc
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_uopc
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_uopc
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_uopc
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_uopc
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_uopc
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_uopc
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_uopc
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_uopc
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_uopc
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_uopc
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_uopc
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_uopc
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_uopc
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_uopc
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_uopc
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_uopc
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_uopc
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_uopc
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_is_rvc =
    _GEN_346
      ? _slots_31_io_uop_is_rvc
      : _GEN_343
          ? _slots_30_io_uop_is_rvc
          : _GEN_335
              ? _slots_29_io_uop_is_rvc
              : _GEN_326
                  ? _slots_28_io_uop_is_rvc
                  : _GEN_317
                      ? _slots_27_io_uop_is_rvc
                      : _GEN_308
                          ? _slots_26_io_uop_is_rvc
                          : _GEN_299
                              ? _slots_25_io_uop_is_rvc
                              : _GEN_290
                                  ? _slots_24_io_uop_is_rvc
                                  : _GEN_281
                                      ? _slots_23_io_uop_is_rvc
                                      : _GEN_272
                                          ? _slots_22_io_uop_is_rvc
                                          : _GEN_263
                                              ? _slots_21_io_uop_is_rvc
                                              : _GEN_254
                                                  ? _slots_20_io_uop_is_rvc
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_is_rvc
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_is_rvc
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_is_rvc
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_is_rvc
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_is_rvc
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_is_rvc
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_is_rvc
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_is_rvc
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_is_rvc
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_is_rvc
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_is_rvc
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_is_rvc
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_is_rvc
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_is_rvc
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_is_rvc
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_is_rvc
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_is_rvc
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_is_rvc
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_is_rvc
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_is_rvc;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_fu_code =
    _GEN_346
      ? _slots_31_io_uop_fu_code
      : _GEN_343
          ? _slots_30_io_uop_fu_code
          : _GEN_335
              ? _slots_29_io_uop_fu_code
              : _GEN_326
                  ? _slots_28_io_uop_fu_code
                  : _GEN_317
                      ? _slots_27_io_uop_fu_code
                      : _GEN_308
                          ? _slots_26_io_uop_fu_code
                          : _GEN_299
                              ? _slots_25_io_uop_fu_code
                              : _GEN_290
                                  ? _slots_24_io_uop_fu_code
                                  : _GEN_281
                                      ? _slots_23_io_uop_fu_code
                                      : _GEN_272
                                          ? _slots_22_io_uop_fu_code
                                          : _GEN_263
                                              ? _slots_21_io_uop_fu_code
                                              : _GEN_254
                                                  ? _slots_20_io_uop_fu_code
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_fu_code
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_fu_code
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_fu_code
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_fu_code
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_fu_code
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_fu_code
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_fu_code
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_fu_code
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_fu_code
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_fu_code
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_fu_code
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_fu_code
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_fu_code
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_fu_code
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_fu_code
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_fu_code
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_fu_code
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_fu_code
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_fu_code
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_fu_code
                                                                                                                                  : 10'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_iw_p1_poisoned =
    _GEN_346
      ? _slots_31_io_uop_iw_p1_poisoned
      : _GEN_343
          ? _slots_30_io_uop_iw_p1_poisoned
          : _GEN_335
              ? _slots_29_io_uop_iw_p1_poisoned
              : _GEN_326
                  ? _slots_28_io_uop_iw_p1_poisoned
                  : _GEN_317
                      ? _slots_27_io_uop_iw_p1_poisoned
                      : _GEN_308
                          ? _slots_26_io_uop_iw_p1_poisoned
                          : _GEN_299
                              ? _slots_25_io_uop_iw_p1_poisoned
                              : _GEN_290
                                  ? _slots_24_io_uop_iw_p1_poisoned
                                  : _GEN_281
                                      ? _slots_23_io_uop_iw_p1_poisoned
                                      : _GEN_272
                                          ? _slots_22_io_uop_iw_p1_poisoned
                                          : _GEN_263
                                              ? _slots_21_io_uop_iw_p1_poisoned
                                              : _GEN_254
                                                  ? _slots_20_io_uop_iw_p1_poisoned
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_iw_p1_poisoned
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_iw_p1_poisoned
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_iw_p1_poisoned
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_iw_p1_poisoned
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_iw_p1_poisoned
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_iw_p1_poisoned
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_iw_p1_poisoned
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_iw_p1_poisoned
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_iw_p1_poisoned
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_iw_p1_poisoned
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_iw_p1_poisoned
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_iw_p1_poisoned
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_iw_p1_poisoned
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_iw_p1_poisoned
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_iw_p1_poisoned
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_iw_p1_poisoned
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_iw_p1_poisoned
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_iw_p1_poisoned
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_iw_p1_poisoned
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_iw_p1_poisoned;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_iw_p2_poisoned =
    _GEN_346
      ? _slots_31_io_uop_iw_p2_poisoned
      : _GEN_343
          ? _slots_30_io_uop_iw_p2_poisoned
          : _GEN_335
              ? _slots_29_io_uop_iw_p2_poisoned
              : _GEN_326
                  ? _slots_28_io_uop_iw_p2_poisoned
                  : _GEN_317
                      ? _slots_27_io_uop_iw_p2_poisoned
                      : _GEN_308
                          ? _slots_26_io_uop_iw_p2_poisoned
                          : _GEN_299
                              ? _slots_25_io_uop_iw_p2_poisoned
                              : _GEN_290
                                  ? _slots_24_io_uop_iw_p2_poisoned
                                  : _GEN_281
                                      ? _slots_23_io_uop_iw_p2_poisoned
                                      : _GEN_272
                                          ? _slots_22_io_uop_iw_p2_poisoned
                                          : _GEN_263
                                              ? _slots_21_io_uop_iw_p2_poisoned
                                              : _GEN_254
                                                  ? _slots_20_io_uop_iw_p2_poisoned
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_iw_p2_poisoned
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_iw_p2_poisoned
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_iw_p2_poisoned
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_iw_p2_poisoned
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_iw_p2_poisoned
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_iw_p2_poisoned
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_iw_p2_poisoned
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_iw_p2_poisoned
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_iw_p2_poisoned
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_iw_p2_poisoned
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_iw_p2_poisoned
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_iw_p2_poisoned
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_iw_p2_poisoned
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_iw_p2_poisoned
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_iw_p2_poisoned
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_iw_p2_poisoned
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_iw_p2_poisoned
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_iw_p2_poisoned
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_iw_p2_poisoned
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_iw_p2_poisoned;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_is_br =
    _GEN_346
      ? _slots_31_io_uop_is_br
      : _GEN_343
          ? _slots_30_io_uop_is_br
          : _GEN_335
              ? _slots_29_io_uop_is_br
              : _GEN_326
                  ? _slots_28_io_uop_is_br
                  : _GEN_317
                      ? _slots_27_io_uop_is_br
                      : _GEN_308
                          ? _slots_26_io_uop_is_br
                          : _GEN_299
                              ? _slots_25_io_uop_is_br
                              : _GEN_290
                                  ? _slots_24_io_uop_is_br
                                  : _GEN_281
                                      ? _slots_23_io_uop_is_br
                                      : _GEN_272
                                          ? _slots_22_io_uop_is_br
                                          : _GEN_263
                                              ? _slots_21_io_uop_is_br
                                              : _GEN_254
                                                  ? _slots_20_io_uop_is_br
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_is_br
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_is_br
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_is_br
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_is_br
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_is_br
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_is_br
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_is_br
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_is_br
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_is_br
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_is_br
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_is_br
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_is_br
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_is_br
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_is_br
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_is_br
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_is_br
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_is_br
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_is_br
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_is_br
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_is_br;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_is_jalr =
    _GEN_346
      ? _slots_31_io_uop_is_jalr
      : _GEN_343
          ? _slots_30_io_uop_is_jalr
          : _GEN_335
              ? _slots_29_io_uop_is_jalr
              : _GEN_326
                  ? _slots_28_io_uop_is_jalr
                  : _GEN_317
                      ? _slots_27_io_uop_is_jalr
                      : _GEN_308
                          ? _slots_26_io_uop_is_jalr
                          : _GEN_299
                              ? _slots_25_io_uop_is_jalr
                              : _GEN_290
                                  ? _slots_24_io_uop_is_jalr
                                  : _GEN_281
                                      ? _slots_23_io_uop_is_jalr
                                      : _GEN_272
                                          ? _slots_22_io_uop_is_jalr
                                          : _GEN_263
                                              ? _slots_21_io_uop_is_jalr
                                              : _GEN_254
                                                  ? _slots_20_io_uop_is_jalr
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_is_jalr
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_is_jalr
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_is_jalr
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_is_jalr
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_is_jalr
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_is_jalr
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_is_jalr
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_is_jalr
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_is_jalr
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_is_jalr
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_is_jalr
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_is_jalr
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_is_jalr
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_is_jalr
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_is_jalr
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_is_jalr
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_is_jalr
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_is_jalr
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_is_jalr
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_is_jalr;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_is_jal =
    _GEN_346
      ? _slots_31_io_uop_is_jal
      : _GEN_343
          ? _slots_30_io_uop_is_jal
          : _GEN_335
              ? _slots_29_io_uop_is_jal
              : _GEN_326
                  ? _slots_28_io_uop_is_jal
                  : _GEN_317
                      ? _slots_27_io_uop_is_jal
                      : _GEN_308
                          ? _slots_26_io_uop_is_jal
                          : _GEN_299
                              ? _slots_25_io_uop_is_jal
                              : _GEN_290
                                  ? _slots_24_io_uop_is_jal
                                  : _GEN_281
                                      ? _slots_23_io_uop_is_jal
                                      : _GEN_272
                                          ? _slots_22_io_uop_is_jal
                                          : _GEN_263
                                              ? _slots_21_io_uop_is_jal
                                              : _GEN_254
                                                  ? _slots_20_io_uop_is_jal
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_is_jal
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_is_jal
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_is_jal
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_is_jal
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_is_jal
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_is_jal
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_is_jal
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_is_jal
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_is_jal
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_is_jal
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_is_jal
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_is_jal
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_is_jal
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_is_jal
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_is_jal
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_is_jal
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_is_jal
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_is_jal
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_is_jal
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_is_jal;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_is_sfb =
    _GEN_346
      ? _slots_31_io_uop_is_sfb
      : _GEN_343
          ? _slots_30_io_uop_is_sfb
          : _GEN_335
              ? _slots_29_io_uop_is_sfb
              : _GEN_326
                  ? _slots_28_io_uop_is_sfb
                  : _GEN_317
                      ? _slots_27_io_uop_is_sfb
                      : _GEN_308
                          ? _slots_26_io_uop_is_sfb
                          : _GEN_299
                              ? _slots_25_io_uop_is_sfb
                              : _GEN_290
                                  ? _slots_24_io_uop_is_sfb
                                  : _GEN_281
                                      ? _slots_23_io_uop_is_sfb
                                      : _GEN_272
                                          ? _slots_22_io_uop_is_sfb
                                          : _GEN_263
                                              ? _slots_21_io_uop_is_sfb
                                              : _GEN_254
                                                  ? _slots_20_io_uop_is_sfb
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_is_sfb
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_is_sfb
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_is_sfb
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_is_sfb
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_is_sfb
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_is_sfb
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_is_sfb
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_is_sfb
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_is_sfb
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_is_sfb
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_is_sfb
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_is_sfb
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_is_sfb
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_is_sfb
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_is_sfb
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_is_sfb
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_is_sfb
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_is_sfb
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_is_sfb
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_is_sfb;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_br_mask =
    _GEN_346
      ? _slots_31_io_uop_br_mask
      : _GEN_343
          ? _slots_30_io_uop_br_mask
          : _GEN_335
              ? _slots_29_io_uop_br_mask
              : _GEN_326
                  ? _slots_28_io_uop_br_mask
                  : _GEN_317
                      ? _slots_27_io_uop_br_mask
                      : _GEN_308
                          ? _slots_26_io_uop_br_mask
                          : _GEN_299
                              ? _slots_25_io_uop_br_mask
                              : _GEN_290
                                  ? _slots_24_io_uop_br_mask
                                  : _GEN_281
                                      ? _slots_23_io_uop_br_mask
                                      : _GEN_272
                                          ? _slots_22_io_uop_br_mask
                                          : _GEN_263
                                              ? _slots_21_io_uop_br_mask
                                              : _GEN_254
                                                  ? _slots_20_io_uop_br_mask
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_br_mask
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_br_mask
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_br_mask
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_br_mask
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_br_mask
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_br_mask
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_br_mask
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_br_mask
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_br_mask
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_br_mask
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_br_mask
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_br_mask
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_br_mask
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_br_mask
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_br_mask
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_br_mask
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_br_mask
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_br_mask
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_br_mask
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_br_mask
                                                                                                                                  : 16'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_br_tag =
    _GEN_346
      ? _slots_31_io_uop_br_tag
      : _GEN_343
          ? _slots_30_io_uop_br_tag
          : _GEN_335
              ? _slots_29_io_uop_br_tag
              : _GEN_326
                  ? _slots_28_io_uop_br_tag
                  : _GEN_317
                      ? _slots_27_io_uop_br_tag
                      : _GEN_308
                          ? _slots_26_io_uop_br_tag
                          : _GEN_299
                              ? _slots_25_io_uop_br_tag
                              : _GEN_290
                                  ? _slots_24_io_uop_br_tag
                                  : _GEN_281
                                      ? _slots_23_io_uop_br_tag
                                      : _GEN_272
                                          ? _slots_22_io_uop_br_tag
                                          : _GEN_263
                                              ? _slots_21_io_uop_br_tag
                                              : _GEN_254
                                                  ? _slots_20_io_uop_br_tag
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_br_tag
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_br_tag
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_br_tag
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_br_tag
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_br_tag
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_br_tag
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_br_tag
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_br_tag
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_br_tag
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_br_tag
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_br_tag
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_br_tag
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_br_tag
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_br_tag
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_br_tag
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_br_tag
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_br_tag
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_br_tag
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_br_tag
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_br_tag
                                                                                                                                  : 4'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_ftq_idx =
    _GEN_346
      ? _slots_31_io_uop_ftq_idx
      : _GEN_343
          ? _slots_30_io_uop_ftq_idx
          : _GEN_335
              ? _slots_29_io_uop_ftq_idx
              : _GEN_326
                  ? _slots_28_io_uop_ftq_idx
                  : _GEN_317
                      ? _slots_27_io_uop_ftq_idx
                      : _GEN_308
                          ? _slots_26_io_uop_ftq_idx
                          : _GEN_299
                              ? _slots_25_io_uop_ftq_idx
                              : _GEN_290
                                  ? _slots_24_io_uop_ftq_idx
                                  : _GEN_281
                                      ? _slots_23_io_uop_ftq_idx
                                      : _GEN_272
                                          ? _slots_22_io_uop_ftq_idx
                                          : _GEN_263
                                              ? _slots_21_io_uop_ftq_idx
                                              : _GEN_254
                                                  ? _slots_20_io_uop_ftq_idx
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_ftq_idx
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_ftq_idx
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_ftq_idx
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_ftq_idx
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_ftq_idx
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_ftq_idx
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_ftq_idx
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_ftq_idx
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_ftq_idx
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_ftq_idx
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_ftq_idx
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_ftq_idx
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_ftq_idx
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_ftq_idx
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_ftq_idx
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_ftq_idx
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_ftq_idx
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_ftq_idx
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_ftq_idx
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_ftq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_2_edge_inst =
    _GEN_346
      ? _slots_31_io_uop_edge_inst
      : _GEN_343
          ? _slots_30_io_uop_edge_inst
          : _GEN_335
              ? _slots_29_io_uop_edge_inst
              : _GEN_326
                  ? _slots_28_io_uop_edge_inst
                  : _GEN_317
                      ? _slots_27_io_uop_edge_inst
                      : _GEN_308
                          ? _slots_26_io_uop_edge_inst
                          : _GEN_299
                              ? _slots_25_io_uop_edge_inst
                              : _GEN_290
                                  ? _slots_24_io_uop_edge_inst
                                  : _GEN_281
                                      ? _slots_23_io_uop_edge_inst
                                      : _GEN_272
                                          ? _slots_22_io_uop_edge_inst
                                          : _GEN_263
                                              ? _slots_21_io_uop_edge_inst
                                              : _GEN_254
                                                  ? _slots_20_io_uop_edge_inst
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_edge_inst
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_edge_inst
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_edge_inst
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_edge_inst
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_edge_inst
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_edge_inst
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_edge_inst
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_edge_inst
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_edge_inst
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_edge_inst
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_edge_inst
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_edge_inst
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_edge_inst
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_edge_inst
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_edge_inst
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_edge_inst
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_edge_inst
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_edge_inst
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_edge_inst
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_edge_inst;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_pc_lob =
    _GEN_346
      ? _slots_31_io_uop_pc_lob
      : _GEN_343
          ? _slots_30_io_uop_pc_lob
          : _GEN_335
              ? _slots_29_io_uop_pc_lob
              : _GEN_326
                  ? _slots_28_io_uop_pc_lob
                  : _GEN_317
                      ? _slots_27_io_uop_pc_lob
                      : _GEN_308
                          ? _slots_26_io_uop_pc_lob
                          : _GEN_299
                              ? _slots_25_io_uop_pc_lob
                              : _GEN_290
                                  ? _slots_24_io_uop_pc_lob
                                  : _GEN_281
                                      ? _slots_23_io_uop_pc_lob
                                      : _GEN_272
                                          ? _slots_22_io_uop_pc_lob
                                          : _GEN_263
                                              ? _slots_21_io_uop_pc_lob
                                              : _GEN_254
                                                  ? _slots_20_io_uop_pc_lob
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_pc_lob
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_pc_lob
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_pc_lob
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_pc_lob
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_pc_lob
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_pc_lob
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_pc_lob
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_pc_lob
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_pc_lob
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_pc_lob
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_pc_lob
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_pc_lob
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_pc_lob
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_pc_lob
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_pc_lob
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_pc_lob
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_pc_lob
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_pc_lob
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_pc_lob
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_pc_lob
                                                                                                                                  : 6'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_taken =
    _GEN_346
      ? _slots_31_io_uop_taken
      : _GEN_343
          ? _slots_30_io_uop_taken
          : _GEN_335
              ? _slots_29_io_uop_taken
              : _GEN_326
                  ? _slots_28_io_uop_taken
                  : _GEN_317
                      ? _slots_27_io_uop_taken
                      : _GEN_308
                          ? _slots_26_io_uop_taken
                          : _GEN_299
                              ? _slots_25_io_uop_taken
                              : _GEN_290
                                  ? _slots_24_io_uop_taken
                                  : _GEN_281
                                      ? _slots_23_io_uop_taken
                                      : _GEN_272
                                          ? _slots_22_io_uop_taken
                                          : _GEN_263
                                              ? _slots_21_io_uop_taken
                                              : _GEN_254
                                                  ? _slots_20_io_uop_taken
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_taken
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_taken
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_taken
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_taken
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_taken
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_taken
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_taken
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_taken
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_taken
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_taken
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_taken
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_taken
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_taken
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_taken
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_taken
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_taken
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_taken
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_taken
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_taken
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_taken;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_imm_packed =
    _GEN_346
      ? _slots_31_io_uop_imm_packed
      : _GEN_343
          ? _slots_30_io_uop_imm_packed
          : _GEN_335
              ? _slots_29_io_uop_imm_packed
              : _GEN_326
                  ? _slots_28_io_uop_imm_packed
                  : _GEN_317
                      ? _slots_27_io_uop_imm_packed
                      : _GEN_308
                          ? _slots_26_io_uop_imm_packed
                          : _GEN_299
                              ? _slots_25_io_uop_imm_packed
                              : _GEN_290
                                  ? _slots_24_io_uop_imm_packed
                                  : _GEN_281
                                      ? _slots_23_io_uop_imm_packed
                                      : _GEN_272
                                          ? _slots_22_io_uop_imm_packed
                                          : _GEN_263
                                              ? _slots_21_io_uop_imm_packed
                                              : _GEN_254
                                                  ? _slots_20_io_uop_imm_packed
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_imm_packed
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_imm_packed
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_imm_packed
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_imm_packed
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_imm_packed
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_imm_packed
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_imm_packed
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_imm_packed
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_imm_packed
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_imm_packed
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_imm_packed
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_imm_packed
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_imm_packed
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_imm_packed
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_imm_packed
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_imm_packed
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_imm_packed
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_imm_packed
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_imm_packed
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_imm_packed
                                                                                                                                  : 20'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_rob_idx =
    _GEN_346
      ? _slots_31_io_uop_rob_idx
      : _GEN_343
          ? _slots_30_io_uop_rob_idx
          : _GEN_335
              ? _slots_29_io_uop_rob_idx
              : _GEN_326
                  ? _slots_28_io_uop_rob_idx
                  : _GEN_317
                      ? _slots_27_io_uop_rob_idx
                      : _GEN_308
                          ? _slots_26_io_uop_rob_idx
                          : _GEN_299
                              ? _slots_25_io_uop_rob_idx
                              : _GEN_290
                                  ? _slots_24_io_uop_rob_idx
                                  : _GEN_281
                                      ? _slots_23_io_uop_rob_idx
                                      : _GEN_272
                                          ? _slots_22_io_uop_rob_idx
                                          : _GEN_263
                                              ? _slots_21_io_uop_rob_idx
                                              : _GEN_254
                                                  ? _slots_20_io_uop_rob_idx
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_rob_idx
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_rob_idx
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_rob_idx
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_rob_idx
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_rob_idx
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_rob_idx
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_rob_idx
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_rob_idx
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_rob_idx
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_rob_idx
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_rob_idx
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_rob_idx
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_rob_idx
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_rob_idx
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_rob_idx
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_rob_idx
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_rob_idx
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_rob_idx
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_rob_idx
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_rob_idx
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_ldq_idx =
    _GEN_346
      ? _slots_31_io_uop_ldq_idx
      : _GEN_343
          ? _slots_30_io_uop_ldq_idx
          : _GEN_335
              ? _slots_29_io_uop_ldq_idx
              : _GEN_326
                  ? _slots_28_io_uop_ldq_idx
                  : _GEN_317
                      ? _slots_27_io_uop_ldq_idx
                      : _GEN_308
                          ? _slots_26_io_uop_ldq_idx
                          : _GEN_299
                              ? _slots_25_io_uop_ldq_idx
                              : _GEN_290
                                  ? _slots_24_io_uop_ldq_idx
                                  : _GEN_281
                                      ? _slots_23_io_uop_ldq_idx
                                      : _GEN_272
                                          ? _slots_22_io_uop_ldq_idx
                                          : _GEN_263
                                              ? _slots_21_io_uop_ldq_idx
                                              : _GEN_254
                                                  ? _slots_20_io_uop_ldq_idx
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_ldq_idx
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_ldq_idx
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_ldq_idx
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_ldq_idx
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_ldq_idx
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_ldq_idx
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_ldq_idx
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_ldq_idx
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_ldq_idx
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_ldq_idx
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_ldq_idx
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_ldq_idx
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_ldq_idx
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_ldq_idx
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_ldq_idx
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_ldq_idx
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_ldq_idx
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_ldq_idx
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_ldq_idx
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_ldq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_2_stq_idx =
    _GEN_346
      ? _slots_31_io_uop_stq_idx
      : _GEN_343
          ? _slots_30_io_uop_stq_idx
          : _GEN_335
              ? _slots_29_io_uop_stq_idx
              : _GEN_326
                  ? _slots_28_io_uop_stq_idx
                  : _GEN_317
                      ? _slots_27_io_uop_stq_idx
                      : _GEN_308
                          ? _slots_26_io_uop_stq_idx
                          : _GEN_299
                              ? _slots_25_io_uop_stq_idx
                              : _GEN_290
                                  ? _slots_24_io_uop_stq_idx
                                  : _GEN_281
                                      ? _slots_23_io_uop_stq_idx
                                      : _GEN_272
                                          ? _slots_22_io_uop_stq_idx
                                          : _GEN_263
                                              ? _slots_21_io_uop_stq_idx
                                              : _GEN_254
                                                  ? _slots_20_io_uop_stq_idx
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_stq_idx
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_stq_idx
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_stq_idx
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_stq_idx
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_stq_idx
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_stq_idx
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_stq_idx
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_stq_idx
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_stq_idx
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_stq_idx
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_stq_idx
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_stq_idx
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_stq_idx
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_stq_idx
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_stq_idx
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_stq_idx
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_stq_idx
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_stq_idx
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_stq_idx
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_stq_idx
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_2_pdst =
    _GEN_346
      ? _slots_31_io_uop_pdst
      : _GEN_343
          ? _slots_30_io_uop_pdst
          : _GEN_335
              ? _slots_29_io_uop_pdst
              : _GEN_326
                  ? _slots_28_io_uop_pdst
                  : _GEN_317
                      ? _slots_27_io_uop_pdst
                      : _GEN_308
                          ? _slots_26_io_uop_pdst
                          : _GEN_299
                              ? _slots_25_io_uop_pdst
                              : _GEN_290
                                  ? _slots_24_io_uop_pdst
                                  : _GEN_281
                                      ? _slots_23_io_uop_pdst
                                      : _GEN_272
                                          ? _slots_22_io_uop_pdst
                                          : _GEN_263
                                              ? _slots_21_io_uop_pdst
                                              : _GEN_254
                                                  ? _slots_20_io_uop_pdst
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_pdst
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_pdst
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_pdst
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_pdst
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_pdst
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_pdst
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_pdst
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_pdst
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_pdst
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_pdst
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_pdst
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_pdst
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_pdst
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_pdst
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_pdst
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_pdst
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_pdst
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_pdst
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_pdst
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_pdst
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_prs1 =
    _GEN_346
      ? _slots_31_io_uop_prs1
      : _GEN_343
          ? _slots_30_io_uop_prs1
          : _GEN_335
              ? _slots_29_io_uop_prs1
              : _GEN_326
                  ? _slots_28_io_uop_prs1
                  : _GEN_317
                      ? _slots_27_io_uop_prs1
                      : _GEN_308
                          ? _slots_26_io_uop_prs1
                          : _GEN_299
                              ? _slots_25_io_uop_prs1
                              : _GEN_290
                                  ? _slots_24_io_uop_prs1
                                  : _GEN_281
                                      ? _slots_23_io_uop_prs1
                                      : _GEN_272
                                          ? _slots_22_io_uop_prs1
                                          : _GEN_263
                                              ? _slots_21_io_uop_prs1
                                              : _GEN_254
                                                  ? _slots_20_io_uop_prs1
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_prs1
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_prs1
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_prs1
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_prs1
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_prs1
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_prs1
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_prs1
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_prs1
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_prs1
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_prs1
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_prs1
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_prs1
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_prs1
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_prs1
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_prs1
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_prs1
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_prs1
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_prs1
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_prs1
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_prs1
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:98:25, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_prs2 =
    _GEN_346
      ? _slots_31_io_uop_prs2
      : _GEN_343
          ? _slots_30_io_uop_prs2
          : _GEN_335
              ? _slots_29_io_uop_prs2
              : _GEN_326
                  ? _slots_28_io_uop_prs2
                  : _GEN_317
                      ? _slots_27_io_uop_prs2
                      : _GEN_308
                          ? _slots_26_io_uop_prs2
                          : _GEN_299
                              ? _slots_25_io_uop_prs2
                              : _GEN_290
                                  ? _slots_24_io_uop_prs2
                                  : _GEN_281
                                      ? _slots_23_io_uop_prs2
                                      : _GEN_272
                                          ? _slots_22_io_uop_prs2
                                          : _GEN_263
                                              ? _slots_21_io_uop_prs2
                                              : _GEN_254
                                                  ? _slots_20_io_uop_prs2
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_prs2
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_prs2
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_prs2
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_prs2
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_prs2
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_prs2
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_prs2
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_prs2
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_prs2
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_prs2
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_prs2
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_prs2
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_prs2
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_prs2
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_prs2
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_prs2
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_prs2
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_prs2
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_prs2
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_prs2
                                                                                                                                  : 7'h0;	// consts.scala:270:20, issue-unit-age-ordered.scala:99:25, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_bypassable =
    _GEN_346
      ? _slots_31_io_uop_bypassable
      : _GEN_343
          ? _slots_30_io_uop_bypassable
          : _GEN_335
              ? _slots_29_io_uop_bypassable
              : _GEN_326
                  ? _slots_28_io_uop_bypassable
                  : _GEN_317
                      ? _slots_27_io_uop_bypassable
                      : _GEN_308
                          ? _slots_26_io_uop_bypassable
                          : _GEN_299
                              ? _slots_25_io_uop_bypassable
                              : _GEN_290
                                  ? _slots_24_io_uop_bypassable
                                  : _GEN_281
                                      ? _slots_23_io_uop_bypassable
                                      : _GEN_272
                                          ? _slots_22_io_uop_bypassable
                                          : _GEN_263
                                              ? _slots_21_io_uop_bypassable
                                              : _GEN_254
                                                  ? _slots_20_io_uop_bypassable
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_bypassable
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_bypassable
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_bypassable
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_bypassable
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_bypassable
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_bypassable
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_bypassable
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_bypassable
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_bypassable
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_bypassable
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_bypassable
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_bypassable
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_bypassable
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_bypassable
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_bypassable
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_bypassable
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_bypassable
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_bypassable
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_bypassable
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_bypassable;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_mem_cmd =
    _GEN_346
      ? _slots_31_io_uop_mem_cmd
      : _GEN_343
          ? _slots_30_io_uop_mem_cmd
          : _GEN_335
              ? _slots_29_io_uop_mem_cmd
              : _GEN_326
                  ? _slots_28_io_uop_mem_cmd
                  : _GEN_317
                      ? _slots_27_io_uop_mem_cmd
                      : _GEN_308
                          ? _slots_26_io_uop_mem_cmd
                          : _GEN_299
                              ? _slots_25_io_uop_mem_cmd
                              : _GEN_290
                                  ? _slots_24_io_uop_mem_cmd
                                  : _GEN_281
                                      ? _slots_23_io_uop_mem_cmd
                                      : _GEN_272
                                          ? _slots_22_io_uop_mem_cmd
                                          : _GEN_263
                                              ? _slots_21_io_uop_mem_cmd
                                              : _GEN_254
                                                  ? _slots_20_io_uop_mem_cmd
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_mem_cmd
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_mem_cmd
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_mem_cmd
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_mem_cmd
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_mem_cmd
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_mem_cmd
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_mem_cmd
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_mem_cmd
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_mem_cmd
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_mem_cmd
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_mem_cmd
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_mem_cmd
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_mem_cmd
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_mem_cmd
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_mem_cmd
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_mem_cmd
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_mem_cmd
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_mem_cmd
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_mem_cmd
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_mem_cmd
                                                                                                                                  : 5'h0;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73, :154:28
  assign io_iss_uops_2_is_amo =
    _GEN_346
      ? _slots_31_io_uop_is_amo
      : _GEN_343
          ? _slots_30_io_uop_is_amo
          : _GEN_335
              ? _slots_29_io_uop_is_amo
              : _GEN_326
                  ? _slots_28_io_uop_is_amo
                  : _GEN_317
                      ? _slots_27_io_uop_is_amo
                      : _GEN_308
                          ? _slots_26_io_uop_is_amo
                          : _GEN_299
                              ? _slots_25_io_uop_is_amo
                              : _GEN_290
                                  ? _slots_24_io_uop_is_amo
                                  : _GEN_281
                                      ? _slots_23_io_uop_is_amo
                                      : _GEN_272
                                          ? _slots_22_io_uop_is_amo
                                          : _GEN_263
                                              ? _slots_21_io_uop_is_amo
                                              : _GEN_254
                                                  ? _slots_20_io_uop_is_amo
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_is_amo
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_is_amo
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_is_amo
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_is_amo
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_is_amo
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_is_amo
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_is_amo
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_is_amo
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_is_amo
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_is_amo
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_is_amo
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_is_amo
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_is_amo
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_is_amo
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_is_amo
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_is_amo
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_is_amo
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_is_amo
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_is_amo
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_is_amo;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_uses_stq =
    _GEN_346
      ? _slots_31_io_uop_uses_stq
      : _GEN_343
          ? _slots_30_io_uop_uses_stq
          : _GEN_335
              ? _slots_29_io_uop_uses_stq
              : _GEN_326
                  ? _slots_28_io_uop_uses_stq
                  : _GEN_317
                      ? _slots_27_io_uop_uses_stq
                      : _GEN_308
                          ? _slots_26_io_uop_uses_stq
                          : _GEN_299
                              ? _slots_25_io_uop_uses_stq
                              : _GEN_290
                                  ? _slots_24_io_uop_uses_stq
                                  : _GEN_281
                                      ? _slots_23_io_uop_uses_stq
                                      : _GEN_272
                                          ? _slots_22_io_uop_uses_stq
                                          : _GEN_263
                                              ? _slots_21_io_uop_uses_stq
                                              : _GEN_254
                                                  ? _slots_20_io_uop_uses_stq
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_uses_stq
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_uses_stq
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_uses_stq
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_uses_stq
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_uses_stq
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_uses_stq
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_uses_stq
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_uses_stq
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_uses_stq
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_uses_stq
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_uses_stq
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_uses_stq
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_uses_stq
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_uses_stq
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_uses_stq
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_uses_stq
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_uses_stq
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_uses_stq
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_uses_stq
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_uses_stq;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_ldst_val =
    _GEN_346
      ? _slots_31_io_uop_ldst_val
      : _GEN_343
          ? _slots_30_io_uop_ldst_val
          : _GEN_335
              ? _slots_29_io_uop_ldst_val
              : _GEN_326
                  ? _slots_28_io_uop_ldst_val
                  : _GEN_317
                      ? _slots_27_io_uop_ldst_val
                      : _GEN_308
                          ? _slots_26_io_uop_ldst_val
                          : _GEN_299
                              ? _slots_25_io_uop_ldst_val
                              : _GEN_290
                                  ? _slots_24_io_uop_ldst_val
                                  : _GEN_281
                                      ? _slots_23_io_uop_ldst_val
                                      : _GEN_272
                                          ? _slots_22_io_uop_ldst_val
                                          : _GEN_263
                                              ? _slots_21_io_uop_ldst_val
                                              : _GEN_254
                                                  ? _slots_20_io_uop_ldst_val
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_ldst_val
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_ldst_val
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_ldst_val
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_ldst_val
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_ldst_val
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_ldst_val
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_ldst_val
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_ldst_val
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_ldst_val
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_ldst_val
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_ldst_val
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_ldst_val
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_ldst_val
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_ldst_val
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_ldst_val
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_ldst_val
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_ldst_val
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_ldst_val
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_ldst_val
                                                                                                                              : _GEN_75
                                                                                                                                & _slots_0_io_uop_ldst_val;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:153:73
  assign io_iss_uops_2_dst_rtype =
    _GEN_346
      ? _slots_31_io_uop_dst_rtype
      : _GEN_343
          ? _slots_30_io_uop_dst_rtype
          : _GEN_335
              ? _slots_29_io_uop_dst_rtype
              : _GEN_326
                  ? _slots_28_io_uop_dst_rtype
                  : _GEN_317
                      ? _slots_27_io_uop_dst_rtype
                      : _GEN_308
                          ? _slots_26_io_uop_dst_rtype
                          : _GEN_299
                              ? _slots_25_io_uop_dst_rtype
                              : _GEN_290
                                  ? _slots_24_io_uop_dst_rtype
                                  : _GEN_281
                                      ? _slots_23_io_uop_dst_rtype
                                      : _GEN_272
                                          ? _slots_22_io_uop_dst_rtype
                                          : _GEN_263
                                              ? _slots_21_io_uop_dst_rtype
                                              : _GEN_254
                                                  ? _slots_20_io_uop_dst_rtype
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_dst_rtype
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_dst_rtype
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_dst_rtype
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_dst_rtype
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_dst_rtype
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_dst_rtype
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_dst_rtype
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_dst_rtype
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_dst_rtype
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_dst_rtype
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_dst_rtype
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_dst_rtype
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_dst_rtype
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_dst_rtype
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_dst_rtype
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_dst_rtype
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_dst_rtype
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_dst_rtype
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_dst_rtype
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_dst_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:96:22, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_2_lrs1_rtype =
    _GEN_346
      ? _slots_31_io_uop_lrs1_rtype
      : _GEN_343
          ? _slots_30_io_uop_lrs1_rtype
          : _GEN_335
              ? _slots_29_io_uop_lrs1_rtype
              : _GEN_326
                  ? _slots_28_io_uop_lrs1_rtype
                  : _GEN_317
                      ? _slots_27_io_uop_lrs1_rtype
                      : _GEN_308
                          ? _slots_26_io_uop_lrs1_rtype
                          : _GEN_299
                              ? _slots_25_io_uop_lrs1_rtype
                              : _GEN_290
                                  ? _slots_24_io_uop_lrs1_rtype
                                  : _GEN_281
                                      ? _slots_23_io_uop_lrs1_rtype
                                      : _GEN_272
                                          ? _slots_22_io_uop_lrs1_rtype
                                          : _GEN_263
                                              ? _slots_21_io_uop_lrs1_rtype
                                              : _GEN_254
                                                  ? _slots_20_io_uop_lrs1_rtype
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_lrs1_rtype
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_lrs1_rtype
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_lrs1_rtype
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_lrs1_rtype
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_lrs1_rtype
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_lrs1_rtype
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_lrs1_rtype
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_lrs1_rtype
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_lrs1_rtype
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_lrs1_rtype
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_lrs1_rtype
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_lrs1_rtype
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_lrs1_rtype
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_lrs1_rtype
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_lrs1_rtype
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_lrs1_rtype
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_lrs1_rtype
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_lrs1_rtype
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_lrs1_rtype
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_lrs1_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:101:31, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
  assign io_iss_uops_2_lrs2_rtype =
    _GEN_346
      ? _slots_31_io_uop_lrs2_rtype
      : _GEN_343
          ? _slots_30_io_uop_lrs2_rtype
          : _GEN_335
              ? _slots_29_io_uop_lrs2_rtype
              : _GEN_326
                  ? _slots_28_io_uop_lrs2_rtype
                  : _GEN_317
                      ? _slots_27_io_uop_lrs2_rtype
                      : _GEN_308
                          ? _slots_26_io_uop_lrs2_rtype
                          : _GEN_299
                              ? _slots_25_io_uop_lrs2_rtype
                              : _GEN_290
                                  ? _slots_24_io_uop_lrs2_rtype
                                  : _GEN_281
                                      ? _slots_23_io_uop_lrs2_rtype
                                      : _GEN_272
                                          ? _slots_22_io_uop_lrs2_rtype
                                          : _GEN_263
                                              ? _slots_21_io_uop_lrs2_rtype
                                              : _GEN_254
                                                  ? _slots_20_io_uop_lrs2_rtype
                                                  : _GEN_245
                                                      ? _slots_19_io_uop_lrs2_rtype
                                                      : _GEN_236
                                                          ? _slots_18_io_uop_lrs2_rtype
                                                          : _GEN_227
                                                              ? _slots_17_io_uop_lrs2_rtype
                                                              : _GEN_218
                                                                  ? _slots_16_io_uop_lrs2_rtype
                                                                  : _GEN_209
                                                                      ? _slots_15_io_uop_lrs2_rtype
                                                                      : _GEN_200
                                                                          ? _slots_14_io_uop_lrs2_rtype
                                                                          : _GEN_191
                                                                              ? _slots_13_io_uop_lrs2_rtype
                                                                              : _GEN_182
                                                                                  ? _slots_12_io_uop_lrs2_rtype
                                                                                  : _GEN_173
                                                                                      ? _slots_11_io_uop_lrs2_rtype
                                                                                      : _GEN_164
                                                                                          ? _slots_10_io_uop_lrs2_rtype
                                                                                          : _GEN_155
                                                                                              ? _slots_9_io_uop_lrs2_rtype
                                                                                              : _GEN_146
                                                                                                  ? _slots_8_io_uop_lrs2_rtype
                                                                                                  : _GEN_137
                                                                                                      ? _slots_7_io_uop_lrs2_rtype
                                                                                                      : _GEN_128
                                                                                                          ? _slots_6_io_uop_lrs2_rtype
                                                                                                          : _GEN_119
                                                                                                              ? _slots_5_io_uop_lrs2_rtype
                                                                                                              : _GEN_110
                                                                                                                  ? _slots_4_io_uop_lrs2_rtype
                                                                                                                  : _GEN_101
                                                                                                                      ? _slots_3_io_uop_lrs2_rtype
                                                                                                                      : _GEN_92
                                                                                                                          ? _slots_2_io_uop_lrs2_rtype
                                                                                                                          : _GEN_83
                                                                                                                              ? _slots_1_io_uop_lrs2_rtype
                                                                                                                              : _GEN_75
                                                                                                                                  ? _slots_0_io_uop_lrs2_rtype
                                                                                                                                  : 2'h2;	// issue-unit-age-ordered.scala:102:31, :118:{40,56,76}, :121:24, issue-unit.scala:129:30, :153:73
endmodule

